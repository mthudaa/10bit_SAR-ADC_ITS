magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect 238 1527 268 1561
rect 302 1527 340 1561
rect 374 1527 412 1561
rect 446 1527 484 1561
rect 518 1527 556 1561
rect 590 1527 628 1561
rect 662 1527 700 1561
rect 734 1527 772 1561
rect 806 1527 844 1561
rect 878 1527 916 1561
rect 950 1527 988 1561
rect 1022 1527 1060 1561
rect 1094 1527 1132 1561
rect 1166 1527 1204 1561
rect 1238 1527 1276 1561
rect 1310 1527 1348 1561
rect 1382 1527 1420 1561
rect 1454 1527 1492 1561
rect 1526 1527 1564 1561
rect 1598 1527 1636 1561
rect 1670 1527 1708 1561
rect 1742 1527 1780 1561
rect 1814 1527 1852 1561
rect 1886 1527 1924 1561
rect 1958 1527 1996 1561
rect 2030 1527 2068 1561
rect 2102 1527 2140 1561
rect 2174 1527 2212 1561
rect 2246 1527 2284 1561
rect 2318 1527 2356 1561
rect 2390 1527 2428 1561
rect 2462 1527 2500 1561
rect 2534 1527 2572 1561
rect 2606 1527 2644 1561
rect 2678 1527 2716 1561
rect 2750 1527 2788 1561
rect 2822 1527 2852 1561
rect 238 -123 262 -89
rect 296 -123 334 -89
rect 368 -123 406 -89
rect 440 -123 478 -89
rect 512 -123 550 -89
rect 584 -123 622 -89
rect 656 -123 694 -89
rect 728 -123 766 -89
rect 800 -123 838 -89
rect 872 -123 910 -89
rect 944 -123 982 -89
rect 1016 -123 1054 -89
rect 1088 -123 1126 -89
rect 1160 -123 1198 -89
rect 1232 -123 1270 -89
rect 1304 -123 1342 -89
rect 1376 -123 1414 -89
rect 1448 -123 1486 -89
rect 1520 -123 1544 -89
<< viali >>
rect 268 1527 302 1561
rect 340 1527 374 1561
rect 412 1527 446 1561
rect 484 1527 518 1561
rect 556 1527 590 1561
rect 628 1527 662 1561
rect 700 1527 734 1561
rect 772 1527 806 1561
rect 844 1527 878 1561
rect 916 1527 950 1561
rect 988 1527 1022 1561
rect 1060 1527 1094 1561
rect 1132 1527 1166 1561
rect 1204 1527 1238 1561
rect 1276 1527 1310 1561
rect 1348 1527 1382 1561
rect 1420 1527 1454 1561
rect 1492 1527 1526 1561
rect 1564 1527 1598 1561
rect 1636 1527 1670 1561
rect 1708 1527 1742 1561
rect 1780 1527 1814 1561
rect 1852 1527 1886 1561
rect 1924 1527 1958 1561
rect 1996 1527 2030 1561
rect 2068 1527 2102 1561
rect 2140 1527 2174 1561
rect 2212 1527 2246 1561
rect 2284 1527 2318 1561
rect 2356 1527 2390 1561
rect 2428 1527 2462 1561
rect 2500 1527 2534 1561
rect 2572 1527 2606 1561
rect 2644 1527 2678 1561
rect 2716 1527 2750 1561
rect 2788 1527 2822 1561
rect 262 -123 296 -89
rect 334 -123 368 -89
rect 406 -123 440 -89
rect 478 -123 512 -89
rect 550 -123 584 -89
rect 622 -123 656 -89
rect 694 -123 728 -89
rect 766 -123 800 -89
rect 838 -123 872 -89
rect 910 -123 944 -89
rect 982 -123 1016 -89
rect 1054 -123 1088 -89
rect 1126 -123 1160 -89
rect 1198 -123 1232 -89
rect 1270 -123 1304 -89
rect 1342 -123 1376 -89
rect 1414 -123 1448 -89
rect 1486 -123 1520 -89
<< metal1 >>
rect 106 1561 2984 1597
rect 106 1527 268 1561
rect 302 1527 340 1561
rect 374 1527 412 1561
rect 446 1527 484 1561
rect 518 1527 556 1561
rect 590 1527 628 1561
rect 662 1527 700 1561
rect 734 1527 772 1561
rect 806 1527 844 1561
rect 878 1527 916 1561
rect 950 1527 988 1561
rect 1022 1527 1060 1561
rect 1094 1527 1132 1561
rect 1166 1527 1204 1561
rect 1238 1527 1276 1561
rect 1310 1527 1348 1561
rect 1382 1527 1420 1561
rect 1454 1527 1492 1561
rect 1526 1527 1564 1561
rect 1598 1527 1636 1561
rect 1670 1527 1708 1561
rect 1742 1527 1780 1561
rect 1814 1527 1852 1561
rect 1886 1527 1924 1561
rect 1958 1527 1996 1561
rect 2030 1527 2068 1561
rect 2102 1527 2140 1561
rect 2174 1527 2212 1561
rect 2246 1527 2284 1561
rect 2318 1527 2356 1561
rect 2390 1527 2428 1561
rect 2462 1527 2500 1561
rect 2534 1527 2572 1561
rect 2606 1527 2644 1561
rect 2678 1527 2716 1561
rect 2750 1527 2788 1561
rect 2822 1527 2984 1561
rect 106 1521 2984 1527
rect 325 1447 2765 1521
rect 106 1377 284 1401
rect 106 1325 176 1377
rect 228 1325 284 1377
rect 106 1301 284 1325
rect 325 1061 2765 1255
rect 106 915 284 1015
rect 106 569 2984 869
rect 106 423 284 523
rect 316 183 1466 376
rect 166 113 284 137
rect 166 61 176 113
rect 228 61 284 113
rect 166 37 284 61
rect 316 -83 1466 -9
rect 106 -89 2984 -83
rect 106 -123 262 -89
rect 296 -123 334 -89
rect 368 -123 406 -89
rect 440 -123 478 -89
rect 512 -123 550 -89
rect 584 -123 622 -89
rect 656 -123 694 -89
rect 728 -123 766 -89
rect 800 -123 838 -89
rect 872 -123 910 -89
rect 944 -123 982 -89
rect 1016 -123 1054 -89
rect 1088 -123 1126 -89
rect 1160 -123 1198 -89
rect 1232 -123 1270 -89
rect 1304 -123 1342 -89
rect 1376 -123 1414 -89
rect 1448 -123 1486 -89
rect 1520 -123 2984 -89
rect 106 -159 2984 -123
<< via1 >>
rect 176 1325 228 1377
rect 176 61 228 113
<< metal2 >>
rect 176 1377 228 1411
rect 176 113 228 1325
rect 176 27 228 61
use sky130_fd_pr__nfet_01v8_54GLWN  sky130_fd_pr__nfet_01v8_54GLWN_0
timestamp 1750100919
transform 0 1 891 -1 0 87
box -236 -775 236 775
use sky130_fd_pr__pfet_01v8_NMY8JJ  sky130_fd_pr__pfet_01v8_NMY8JJ_0
timestamp 1750100919
transform 0 1 1545 -1 0 965
box -246 -1439 246 1439
use sky130_fd_pr__pfet_01v8_NMY8JJ  XM1
timestamp 1750100919
transform 0 1 1545 -1 0 1351
box -246 -1439 246 1439
use sky130_fd_pr__nfet_01v8_54GLWN  XM3
timestamp 1750100919
transform 0 1 891 -1 0 473
box -236 -775 236 775
<< labels >>
flabel metal1 s 106 1521 238 1597 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 106 1301 176 1401 0 FreeSans 500 0 0 0 IN
port 2 nsew
flabel metal1 s 106 915 284 1015 0 FreeSans 500 0 0 0 CKB
port 3 nsew
flabel metal1 s 106 423 284 523 0 FreeSans 500 0 0 0 CK
port 4 nsew
flabel metal1 s 106 -159 238 -83 0 FreeSans 500 0 0 0 VSS
port 5 nsew
flabel metal1 s 2802 673 2934 749 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
