* NGSPICE file created from sar10b.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hs__fill_8 abstract view
.subckt sky130_fd_sc_hs__fill_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__dfrtp_1 abstract view
.subckt sky130_fd_sc_hs__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__fill_2 abstract view
.subckt sky130_fd_sc_hs__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__dfrtp_2 abstract view
.subckt sky130_fd_sc_hs__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__decap_4 abstract view
.subckt sky130_fd_sc_hs__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__fill_1 abstract view
.subckt sky130_fd_sc_hs__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__clkbuf_1 abstract view
.subckt sky130_fd_sc_hs__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hs__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__and2_1 abstract view
.subckt sky130_fd_sc_hs__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__xor2_1 abstract view
.subckt sky130_fd_sc_hs__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__clkbuf_16 abstract view
.subckt sky130_fd_sc_hs__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nor2_1 abstract view
.subckt sky130_fd_sc_hs__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__a21bo_1 abstract view
.subckt sky130_fd_sc_hs__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__o21a_1 abstract view
.subckt sky130_fd_sc_hs__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__or3b_1 abstract view
.subckt sky130_fd_sc_hs__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nand2_1 abstract view
.subckt sky130_fd_sc_hs__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__or4bb_1 abstract view
.subckt sky130_fd_sc_hs__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__clkbuf_2 abstract view
.subckt sky130_fd_sc_hs__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__buf_8 abstract view
.subckt sky130_fd_sc_hs__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__clkbuf_4 abstract view
.subckt sky130_fd_sc_hs__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__dfxtp_4 abstract view
.subckt sky130_fd_sc_hs__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__dfxtp_1 abstract view
.subckt sky130_fd_sc_hs__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nor3_1 abstract view
.subckt sky130_fd_sc_hs__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__a21oi_1 abstract view
.subckt sky130_fd_sc_hs__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__and3_1 abstract view
.subckt sky130_fd_sc_hs__and3_1 A B C VGND VNB VPB VPWR X
.ends

.subckt sar10b CF[0] CF[1] CF[2] CF[3] CF[4] CF[5] CF[6] CF[7] CF[8] CF[9] CKO CKS
+ CKSB CLK CMP_N CMP_P DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7]
+ DATA[8] DATA[9] EN RDY SWN[0] SWN[1] SWN[2] SWN[3] SWN[4] SWN[5] SWN[6] SWN[7] SWN[8]
+ SWN[9] SWP[0] SWP[1] SWP[2] SWP[3] SWP[4] SWP[5] SWP[6] SWP[7] SWP[8] SWP[9] VGND
+ VPWR
XFILLER_0_3_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_83_ cyclic_flag_0.FINAL net38 net3 VGND VGND VPWR VPWR net18 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_34_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_0_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_66_ net12 net1 net16 VGND VGND VPWR VPWR net35 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_9_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_49_ net4 net14 net16 VGND VGND VPWR VPWR cyclic_flag_0.FINAL sky130_fd_sc_hs__dfrtp_2
XPHY_EDGE_ROW_28_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_12_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_6_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
Xoutput42 net42 VGND VGND VPWR VPWR SWP[4] sky130_fd_sc_hs__clkbuf_1
Xoutput31 net31 VGND VGND VPWR VPWR SWN[3] sky130_fd_sc_hs__clkbuf_1
Xoutput20 net20 VGND VGND VPWR VPWR DATA[2] sky130_fd_sc_hs__clkbuf_1
Xoutput7 net7 VGND VGND VPWR VPWR CF[2] sky130_fd_sc_hs__clkbuf_1
XTAP_TAPCELL_ROW_24_107 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_15_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_82_ cyclic_flag_0.FINAL net39 net3 VGND VGND VPWR VPWR net19 sky130_fd_sc_hs__dfrtp_1
XPHY_EDGE_ROW_0_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_65_ net13 net1 net16 VGND VGND VPWR VPWR net36 sky130_fd_sc_hs__dfrtp_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_48_ net4 net13 net16 VGND VGND VPWR VPWR net14 sky130_fd_sc_hs__dfrtp_1
XTAP_TAPCELL_ROW_18_98 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_79 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_21_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_34_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_1_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
Xoutput43 net43 VGND VGND VPWR VPWR SWP[5] sky130_fd_sc_hs__clkbuf_1
Xoutput32 net32 VGND VGND VPWR VPWR SWN[4] sky130_fd_sc_hs__clkbuf_1
Xoutput21 net21 VGND VGND VPWR VPWR DATA[3] sky130_fd_sc_hs__clkbuf_1
Xoutput8 net8 VGND VGND VPWR VPWR CF[3] sky130_fd_sc_hs__clkbuf_1
Xoutput10 net10 VGND VGND VPWR VPWR CF[5] sky130_fd_sc_hs__clkbuf_1
XTAP_TAPCELL_ROW_24_108 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_7_83 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_81_ cyclic_flag_0.FINAL net40 net3 VGND VGND VPWR VPWR net20 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XTAP_TAPCELL_ROW_12_89 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_64_ net14 net1 net16 VGND VGND VPWR VPWR net37 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_24_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_47_ net4 net12 net16 VGND VGND VPWR VPWR net13 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_18_99 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_19_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_27_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_32_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_16_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
Xoutput44 net44 VGND VGND VPWR VPWR SWP[6] sky130_fd_sc_hs__clkbuf_1
Xoutput33 net33 VGND VGND VPWR VPWR SWN[5] sky130_fd_sc_hs__clkbuf_1
Xoutput22 net22 VGND VGND VPWR VPWR DATA[4] sky130_fd_sc_hs__clkbuf_1
Xoutput9 net9 VGND VGND VPWR VPWR CF[4] sky130_fd_sc_hs__clkbuf_1
Xoutput11 net11 VGND VGND VPWR VPWR CF[6] sky130_fd_sc_hs__clkbuf_1
XTAP_TAPCELL_ROW_32_120 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_27_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_27_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_80_ cyclic_flag_0.FINAL net41 net3 VGND VGND VPWR VPWR net21 sky130_fd_sc_hs__dfrtp_1
XTAP_TAPCELL_ROW_20_101 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_63_ net5 net2 net16 VGND VGND VPWR VPWR net38 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_29_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_0_70 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_46_ net4 net11 net16 VGND VGND VPWR VPWR net12 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_34_6 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_29_ net3 _12_ VGND VGND VPWR VPWR _13_ sky130_fd_sc_hs__and2_1
XFILLER_0_32_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_6_80 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
Xoutput45 net45 VGND VGND VPWR VPWR SWP[7] sky130_fd_sc_hs__clkbuf_1
Xoutput12 net12 VGND VGND VPWR VPWR CF[7] sky130_fd_sc_hs__clkbuf_1
Xoutput34 net34 VGND VGND VPWR VPWR SWN[6] sky130_fd_sc_hs__clkbuf_1
Xoutput23 net23 VGND VGND VPWR VPWR DATA[5] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_27_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_11_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_7_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_13_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_19_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_20_102 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_62_ net6 net2 net16 VGND VGND VPWR VPWR net39 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_4_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_0_71 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_10_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_45_ net4 net10 net16 VGND VGND VPWR VPWR net11 sky130_fd_sc_hs__dfrtp_1
X_28_ clk_div_0.COUNT\[1\] clk_div_0.COUNT\[0\] VGND VGND VPWR VPWR _12_ sky130_fd_sc_hs__xor2_1
XFILLER_0_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_7_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_32_76 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_6_81 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
Xoutput46 net46 VGND VGND VPWR VPWR SWP[8] sky130_fd_sc_hs__clkbuf_1
XPHY_EDGE_ROW_33_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_32_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
Xoutput13 net13 VGND VGND VPWR VPWR CF[8] sky130_fd_sc_hs__clkbuf_1
Xoutput35 net35 VGND VGND VPWR VPWR SWN[7] sky130_fd_sc_hs__clkbuf_1
Xoutput24 net24 VGND VGND VPWR VPWR DATA[6] sky130_fd_sc_hs__clkbuf_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_61_ net7 net2 net16 VGND VGND VPWR VPWR net40 sky130_fd_sc_hs__dfrtp_1
XPHY_EDGE_ROW_20_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
Xclkbuf_1_1__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_1_1__leaf_CLK sky130_fd_sc_hs__clkbuf_16
XFILLER_0_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_13_91 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_72 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_44_ net4 net9 net16 VGND VGND VPWR VPWR net10 sky130_fd_sc_hs__dfrtp_1
X_27_ clk_div_0.COUNT\[0\] _08_ VGND VGND VPWR VPWR _02_ sky130_fd_sc_hs__nor2_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_21_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_1_77 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_16_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
Xoutput47 net47 VGND VGND VPWR VPWR SWP[9] sky130_fd_sc_hs__clkbuf_1
Xoutput14 net14 VGND VGND VPWR VPWR CF[9] sky130_fd_sc_hs__clkbuf_1
Xoutput36 net36 VGND VGND VPWR VPWR SWN[8] sky130_fd_sc_hs__clkbuf_1
Xoutput25 net25 VGND VGND VPWR VPWR DATA[7] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_60_ net8 net2 net16 VGND VGND VPWR VPWR net41 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_10_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_43_ net4 net8 net16 VGND VGND VPWR VPWR net9 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_26_ _11_ VGND VGND VPWR VPWR _01_ sky130_fd_sc_hs__clkbuf_1
XFILLER_0_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_32_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
Xoutput15 net15 VGND VGND VPWR VPWR CKO sky130_fd_sc_hs__clkbuf_1
Xoutput26 net26 VGND VGND VPWR VPWR DATA[8] sky130_fd_sc_hs__clkbuf_1
XTAP_TAPCELL_ROW_26_110 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
Xoutput37 net37 VGND VGND VPWR VPWR SWN[9] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_27_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_27_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_7_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_13_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_42_ net4 net7 net16 VGND VGND VPWR VPWR net8 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_25_ net16 _10_ _09_ VGND VGND VPWR VPWR _11_ sky130_fd_sc_hs__a21bo_1
XFILLER_0_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
Xoutput16 net16 VGND VGND VPWR VPWR CKS sky130_fd_sc_hs__clkbuf_1
Xoutput38 net38 VGND VGND VPWR VPWR SWP[0] sky130_fd_sc_hs__clkbuf_1
Xoutput27 net27 VGND VGND VPWR VPWR DATA[9] sky130_fd_sc_hs__clkbuf_1
XTAP_TAPCELL_ROW_26_111 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_9_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_30_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_7_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_24_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_41_ net4 net6 net16 VGND VGND VPWR VPWR net7 sky130_fd_sc_hs__dfrtp_1
XPHY_EDGE_ROW_24_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_24_ net3 _07_ VGND VGND VPWR VPWR _10_ sky130_fd_sc_hs__and2_1
XFILLER_0_32_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_27_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
Xoutput39 net39 VGND VGND VPWR VPWR SWP[1] sky130_fd_sc_hs__clkbuf_1
Xoutput28 net28 VGND VGND VPWR VPWR SWN[0] sky130_fd_sc_hs__clkbuf_1
Xoutput17 net17 VGND VGND VPWR VPWR CKSB sky130_fd_sc_hs__clkbuf_1
XPHY_EDGE_ROW_11_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_27_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_2_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_28_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_40_ net4 net5 net16 VGND VGND VPWR VPWR net6 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_10_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_9_85 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_23_ net17 _08_ _09_ VGND VGND VPWR VPWR _00_ sky130_fd_sc_hs__o21a_1
XFILLER_0_1_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_21_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_25_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
Xoutput18 net18 VGND VGND VPWR VPWR DATA[0] sky130_fd_sc_hs__clkbuf_1
Xoutput29 net29 VGND VGND VPWR VPWR SWN[1] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_16_95 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_76 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_5_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_19_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_22_ _07_ net16 net3 VGND VGND VPWR VPWR _09_ sky130_fd_sc_hs__or3b_1
XFILLER_0_1_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_10_86 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_16_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
Xoutput19 net19 VGND VGND VPWR VPWR DATA[1] sky130_fd_sc_hs__clkbuf_1
XTAP_TAPCELL_ROW_23_106 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_96 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_24_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_4_49 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_21_ net3 _07_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hs__nand2_1
XTAP_TAPCELL_ROW_10_87 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_32_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_27_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_33_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_28_60 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_4_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_18_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_3_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_20_ clk_div_0.COUNT\[1\] clk_div_0.COUNT\[0\] clk_div_0.COUNT\[2\] clk_div_0.COUNT\[3\]
+ VGND VGND VPWR VPWR _07_ sky130_fd_sc_hs__or4bb_1
XFILLER_0_11_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
Xinput1 CMP_N VGND VGND VPWR VPWR net1 sky130_fd_sc_hs__clkbuf_2
XFILLER_0_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_32_119 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_7_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_23_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_32_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_3_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
Xinput2 CMP_P VGND VGND VPWR VPWR net2 sky130_fd_sc_hs__clkbuf_2
X_79_ cyclic_flag_0.FINAL net42 net3 VGND VGND VPWR VPWR net22 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_17_30 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_17_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_8_72 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_14_75 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_25_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_25_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_5_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_78_ cyclic_flag_0.FINAL net43 net3 VGND VGND VPWR VPWR net23 sky130_fd_sc_hs__dfrtp_1
Xinput3 EN VGND VGND VPWR VPWR net3 sky130_fd_sc_hs__buf_8
XFILLER_0_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_29_115 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_33_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_28_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_30_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
Xinput4 RDY VGND VGND VPWR VPWR net4 sky130_fd_sc_hs__clkbuf_4
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_77_ cyclic_flag_0.FINAL net44 net3 VGND VGND VPWR VPWR net24 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_33_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_21_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_25_32 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_76_ cyclic_flag_0.FINAL net45 net3 VGND VGND VPWR VPWR net25 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_11_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_23_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_59_ net9 net2 net16 VGND VGND VPWR VPWR net42 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_33_87 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_26_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_10_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_28_76 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_75_ cyclic_flag_0.FINAL net46 net3 VGND VGND VPWR VPWR net26 sky130_fd_sc_hs__dfrtp_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_58_ net10 net2 net16 VGND VGND VPWR VPWR net43 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_33_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_7_82 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_8_10 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_30_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_25_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XTAP_TAPCELL_ROW_14_92 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_74_ cyclic_flag_0.FINAL net47 net3 VGND VGND VPWR VPWR net27 sky130_fd_sc_hs__dfrtp_1
XTAP_TAPCELL_ROW_1_73 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_22_57 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_34_122 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_57_ net11 net2 net16 VGND VGND VPWR VPWR net44 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_33_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_33_89 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_30_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_14_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_25_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_10_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_14_93 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_73_ net5 net1 net16 VGND VGND VPWR VPWR net28 sky130_fd_sc_hs__dfrtp_1
XTAP_TAPCELL_ROW_34_123 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_56_ net12 net2 net16 VGND VGND VPWR VPWR net45 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_2_46 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_33_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_39_ net4 net16 net16 VGND VGND VPWR VPWR net5 sky130_fd_sc_hs__dfrtp_1
XTAP_TAPCELL_ROW_22_104 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_14_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_18_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_30_69 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_30_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_17_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_72_ net6 net1 net16 VGND VGND VPWR VPWR net29 sky130_fd_sc_hs__dfrtp_1
XPHY_EDGE_ROW_2_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_34_124 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_55_ net13 net2 net16 VGND VGND VPWR VPWR net46 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_33_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_38_ clknet_1_1__leaf_CLK _01_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hs__dfxtp_4
XTAP_TAPCELL_ROW_22_105 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_31_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_31_91 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_15_92 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_71_ net7 net1 net16 VGND VGND VPWR VPWR net30 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_54_ net14 net2 net16 VGND VGND VPWR VPWR net47 sky130_fd_sc_hs__dfrtp_1
XTAP_TAPCELL_ROW_19_100 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_23_92 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_37_ clknet_1_0__leaf_CLK _00_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hs__dfxtp_1
XFILLER_0_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_8_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_14_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_25_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_70_ net8 net1 net16 VGND VGND VPWR VPWR net31 sky130_fd_sc_hs__dfrtp_1
Xclkbuf_0_CLK CLK VGND VGND VPWR VPWR clknet_0_CLK sky130_fd_sc_hs__clkbuf_16
X_53_ clknet_1_1__leaf_CLK _05_ VGND VGND VPWR VPWR clk_div_0.COUNT\[3\] sky130_fd_sc_hs__dfxtp_1
XFILLER_0_22_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_31_118 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_17_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_36_ _17_ VGND VGND VPWR VPWR _05_ sky130_fd_sc_hs__clkbuf_1
XFILLER_0_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_19_ _06_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hs__clkbuf_1
XFILLER_0_18_60 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_30_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_4_77 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_6_70 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_28_113 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_2_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_52_ clknet_1_1__leaf_CLK _04_ VGND VGND VPWR VPWR clk_div_0.COUNT\[2\] sky130_fd_sc_hs__dfxtp_1
XFILLER_0_12_51 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_33_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_35_ _10_ _16_ VGND VGND VPWR VPWR _17_ sky130_fd_sc_hs__and2_1
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_34_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_18_ net16 cyclic_flag_0.FINAL VGND VGND VPWR VPWR _06_ sky130_fd_sc_hs__and2_1
XTAP_TAPCELL_ROW_17_97 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_78 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_9_92 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_31_83 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_28_114 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_22_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_51_ clknet_1_0__leaf_CLK _03_ VGND VGND VPWR VPWR clk_div_0.COUNT\[1\] sky130_fd_sc_hs__dfxtp_1
XTAP_TAPCELL_ROW_11_88 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_34_ clk_div_0.COUNT\[3\] _14_ VGND VGND VPWR VPWR _16_ sky130_fd_sc_hs__xor2_1
XFILLER_0_23_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_25_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_8_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_31_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_15_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_6_72 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_50_ clknet_1_0__leaf_CLK _02_ VGND VGND VPWR VPWR clk_div_0.COUNT\[0\] sky130_fd_sc_hs__dfxtp_1
X_33_ _08_ _14_ _15_ VGND VGND VPWR VPWR _04_ sky130_fd_sc_hs__nor3_1
XFILLER_0_23_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_23_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_34_51 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_18_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_29_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_15_42 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_12_76 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_32_ clk_div_0.COUNT\[1\] clk_div_0.COUNT\[0\] clk_div_0.COUNT\[2\] VGND VGND VPWR
+ VPWR _15_ sky130_fd_sc_hs__a21oi_1
XFILLER_0_34_30 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_19_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_29_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_9_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XTAP_TAPCELL_ROW_25_109 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_31_ clk_div_0.COUNT\[1\] clk_div_0.COUNT\[0\] clk_div_0.COUNT\[2\] VGND VGND VPWR
+ VPWR _14_ sky130_fd_sc_hs__and3_1
XFILLER_0_23_32 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XTAP_TAPCELL_ROW_12_90 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_31_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_29_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_13_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_16_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_33_121 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_30_ _13_ VGND VGND VPWR VPWR _03_ sky130_fd_sc_hs__clkbuf_1
XFILLER_0_3_87 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_29_32 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_30_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_15_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_23_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_21_103 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_17_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_23_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_8_83 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_29_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_31_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_2_74 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_116 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_34_35 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_18_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_34_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_8_84 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_24_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_29_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_9_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_8_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_34_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_26_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_32_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_15_94 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_75 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_117 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_23_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_69_ net9 net1 net16 VGND VGND VPWR VPWR net32 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_9_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_60 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_15_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_15_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_21_92 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XTAP_TAPCELL_ROW_27_112 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_23_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_34_59 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_68_ net10 net1 net16 VGND VGND VPWR VPWR net33 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_29_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_20_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_31_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
Xoutput40 net40 VGND VGND VPWR VPWR SWP[2] sky130_fd_sc_hs__clkbuf_1
Xoutput5 net5 VGND VGND VPWR VPWR CF[0] sky130_fd_sc_hs__clkbuf_1
XFILLER_0_27_92 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
Xclkbuf_1_0__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_1_0__leaf_CLK sky130_fd_sc_hs__clkbuf_16
XFILLER_0_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_18_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_67_ net11 net1 net16 VGND VGND VPWR VPWR net34 sky130_fd_sc_hs__dfrtp_1
XFILLER_0_29_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_0_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_9_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_15_18 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_26_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_32_60 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
Xoutput41 net41 VGND VGND VPWR VPWR SWP[3] sky130_fd_sc_hs__clkbuf_1
Xoutput30 net30 VGND VGND VPWR VPWR SWN[2] sky130_fd_sc_hs__clkbuf_1
Xoutput6 net6 VGND VGND VPWR VPWR CF[1] sky130_fd_sc_hs__clkbuf_1
.ends

