magic
tech sky130A
magscale 1 2
timestamp 1749307785
<< metal3 >>
rect -2704 4332 -1532 4360
rect -2704 3508 -1616 4332
rect -1552 3508 -1532 4332
rect -2704 3480 -1532 3508
rect -1292 4332 -120 4360
rect -1292 3508 -204 4332
rect -140 3508 -120 4332
rect -1292 3480 -120 3508
rect 120 4332 1292 4360
rect 120 3508 1208 4332
rect 1272 3508 1292 4332
rect 120 3480 1292 3508
rect 1532 4332 2704 4360
rect 1532 3508 2620 4332
rect 2684 3508 2704 4332
rect 1532 3480 2704 3508
rect -2704 3212 -1532 3240
rect -2704 2388 -1616 3212
rect -1552 2388 -1532 3212
rect -2704 2360 -1532 2388
rect -1292 3212 -120 3240
rect -1292 2388 -204 3212
rect -140 2388 -120 3212
rect -1292 2360 -120 2388
rect 120 3212 1292 3240
rect 120 2388 1208 3212
rect 1272 2388 1292 3212
rect 120 2360 1292 2388
rect 1532 3212 2704 3240
rect 1532 2388 2620 3212
rect 2684 2388 2704 3212
rect 1532 2360 2704 2388
rect -2704 2092 -1532 2120
rect -2704 1268 -1616 2092
rect -1552 1268 -1532 2092
rect -2704 1240 -1532 1268
rect -1292 2092 -120 2120
rect -1292 1268 -204 2092
rect -140 1268 -120 2092
rect -1292 1240 -120 1268
rect 120 2092 1292 2120
rect 120 1268 1208 2092
rect 1272 1268 1292 2092
rect 120 1240 1292 1268
rect 1532 2092 2704 2120
rect 1532 1268 2620 2092
rect 2684 1268 2704 2092
rect 1532 1240 2704 1268
rect -2704 972 -1532 1000
rect -2704 148 -1616 972
rect -1552 148 -1532 972
rect -2704 120 -1532 148
rect -1292 972 -120 1000
rect -1292 148 -204 972
rect -140 148 -120 972
rect -1292 120 -120 148
rect 120 972 1292 1000
rect 120 148 1208 972
rect 1272 148 1292 972
rect 120 120 1292 148
rect 1532 972 2704 1000
rect 1532 148 2620 972
rect 2684 148 2704 972
rect 1532 120 2704 148
rect -2704 -148 -1532 -120
rect -2704 -972 -1616 -148
rect -1552 -972 -1532 -148
rect -2704 -1000 -1532 -972
rect -1292 -148 -120 -120
rect -1292 -972 -204 -148
rect -140 -972 -120 -148
rect -1292 -1000 -120 -972
rect 120 -148 1292 -120
rect 120 -972 1208 -148
rect 1272 -972 1292 -148
rect 120 -1000 1292 -972
rect 1532 -148 2704 -120
rect 1532 -972 2620 -148
rect 2684 -972 2704 -148
rect 1532 -1000 2704 -972
rect -2704 -1268 -1532 -1240
rect -2704 -2092 -1616 -1268
rect -1552 -2092 -1532 -1268
rect -2704 -2120 -1532 -2092
rect -1292 -1268 -120 -1240
rect -1292 -2092 -204 -1268
rect -140 -2092 -120 -1268
rect -1292 -2120 -120 -2092
rect 120 -1268 1292 -1240
rect 120 -2092 1208 -1268
rect 1272 -2092 1292 -1268
rect 120 -2120 1292 -2092
rect 1532 -1268 2704 -1240
rect 1532 -2092 2620 -1268
rect 2684 -2092 2704 -1268
rect 1532 -2120 2704 -2092
rect -2704 -2388 -1532 -2360
rect -2704 -3212 -1616 -2388
rect -1552 -3212 -1532 -2388
rect -2704 -3240 -1532 -3212
rect -1292 -2388 -120 -2360
rect -1292 -3212 -204 -2388
rect -140 -3212 -120 -2388
rect -1292 -3240 -120 -3212
rect 120 -2388 1292 -2360
rect 120 -3212 1208 -2388
rect 1272 -3212 1292 -2388
rect 120 -3240 1292 -3212
rect 1532 -2388 2704 -2360
rect 1532 -3212 2620 -2388
rect 2684 -3212 2704 -2388
rect 1532 -3240 2704 -3212
rect -2704 -3508 -1532 -3480
rect -2704 -4332 -1616 -3508
rect -1552 -4332 -1532 -3508
rect -2704 -4360 -1532 -4332
rect -1292 -3508 -120 -3480
rect -1292 -4332 -204 -3508
rect -140 -4332 -120 -3508
rect -1292 -4360 -120 -4332
rect 120 -3508 1292 -3480
rect 120 -4332 1208 -3508
rect 1272 -4332 1292 -3508
rect 120 -4360 1292 -4332
rect 1532 -3508 2704 -3480
rect 1532 -4332 2620 -3508
rect 2684 -4332 2704 -3508
rect 1532 -4360 2704 -4332
<< via3 >>
rect -1616 3508 -1552 4332
rect -204 3508 -140 4332
rect 1208 3508 1272 4332
rect 2620 3508 2684 4332
rect -1616 2388 -1552 3212
rect -204 2388 -140 3212
rect 1208 2388 1272 3212
rect 2620 2388 2684 3212
rect -1616 1268 -1552 2092
rect -204 1268 -140 2092
rect 1208 1268 1272 2092
rect 2620 1268 2684 2092
rect -1616 148 -1552 972
rect -204 148 -140 972
rect 1208 148 1272 972
rect 2620 148 2684 972
rect -1616 -972 -1552 -148
rect -204 -972 -140 -148
rect 1208 -972 1272 -148
rect 2620 -972 2684 -148
rect -1616 -2092 -1552 -1268
rect -204 -2092 -140 -1268
rect 1208 -2092 1272 -1268
rect 2620 -2092 2684 -1268
rect -1616 -3212 -1552 -2388
rect -204 -3212 -140 -2388
rect 1208 -3212 1272 -2388
rect 2620 -3212 2684 -2388
rect -1616 -4332 -1552 -3508
rect -204 -4332 -140 -3508
rect 1208 -4332 1272 -3508
rect 2620 -4332 2684 -3508
<< mimcap >>
rect -2664 4280 -1864 4320
rect -2664 3560 -2624 4280
rect -1904 3560 -1864 4280
rect -2664 3520 -1864 3560
rect -1252 4280 -452 4320
rect -1252 3560 -1212 4280
rect -492 3560 -452 4280
rect -1252 3520 -452 3560
rect 160 4280 960 4320
rect 160 3560 200 4280
rect 920 3560 960 4280
rect 160 3520 960 3560
rect 1572 4280 2372 4320
rect 1572 3560 1612 4280
rect 2332 3560 2372 4280
rect 1572 3520 2372 3560
rect -2664 3160 -1864 3200
rect -2664 2440 -2624 3160
rect -1904 2440 -1864 3160
rect -2664 2400 -1864 2440
rect -1252 3160 -452 3200
rect -1252 2440 -1212 3160
rect -492 2440 -452 3160
rect -1252 2400 -452 2440
rect 160 3160 960 3200
rect 160 2440 200 3160
rect 920 2440 960 3160
rect 160 2400 960 2440
rect 1572 3160 2372 3200
rect 1572 2440 1612 3160
rect 2332 2440 2372 3160
rect 1572 2400 2372 2440
rect -2664 2040 -1864 2080
rect -2664 1320 -2624 2040
rect -1904 1320 -1864 2040
rect -2664 1280 -1864 1320
rect -1252 2040 -452 2080
rect -1252 1320 -1212 2040
rect -492 1320 -452 2040
rect -1252 1280 -452 1320
rect 160 2040 960 2080
rect 160 1320 200 2040
rect 920 1320 960 2040
rect 160 1280 960 1320
rect 1572 2040 2372 2080
rect 1572 1320 1612 2040
rect 2332 1320 2372 2040
rect 1572 1280 2372 1320
rect -2664 920 -1864 960
rect -2664 200 -2624 920
rect -1904 200 -1864 920
rect -2664 160 -1864 200
rect -1252 920 -452 960
rect -1252 200 -1212 920
rect -492 200 -452 920
rect -1252 160 -452 200
rect 160 920 960 960
rect 160 200 200 920
rect 920 200 960 920
rect 160 160 960 200
rect 1572 920 2372 960
rect 1572 200 1612 920
rect 2332 200 2372 920
rect 1572 160 2372 200
rect -2664 -200 -1864 -160
rect -2664 -920 -2624 -200
rect -1904 -920 -1864 -200
rect -2664 -960 -1864 -920
rect -1252 -200 -452 -160
rect -1252 -920 -1212 -200
rect -492 -920 -452 -200
rect -1252 -960 -452 -920
rect 160 -200 960 -160
rect 160 -920 200 -200
rect 920 -920 960 -200
rect 160 -960 960 -920
rect 1572 -200 2372 -160
rect 1572 -920 1612 -200
rect 2332 -920 2372 -200
rect 1572 -960 2372 -920
rect -2664 -1320 -1864 -1280
rect -2664 -2040 -2624 -1320
rect -1904 -2040 -1864 -1320
rect -2664 -2080 -1864 -2040
rect -1252 -1320 -452 -1280
rect -1252 -2040 -1212 -1320
rect -492 -2040 -452 -1320
rect -1252 -2080 -452 -2040
rect 160 -1320 960 -1280
rect 160 -2040 200 -1320
rect 920 -2040 960 -1320
rect 160 -2080 960 -2040
rect 1572 -1320 2372 -1280
rect 1572 -2040 1612 -1320
rect 2332 -2040 2372 -1320
rect 1572 -2080 2372 -2040
rect -2664 -2440 -1864 -2400
rect -2664 -3160 -2624 -2440
rect -1904 -3160 -1864 -2440
rect -2664 -3200 -1864 -3160
rect -1252 -2440 -452 -2400
rect -1252 -3160 -1212 -2440
rect -492 -3160 -452 -2440
rect -1252 -3200 -452 -3160
rect 160 -2440 960 -2400
rect 160 -3160 200 -2440
rect 920 -3160 960 -2440
rect 160 -3200 960 -3160
rect 1572 -2440 2372 -2400
rect 1572 -3160 1612 -2440
rect 2332 -3160 2372 -2440
rect 1572 -3200 2372 -3160
rect -2664 -3560 -1864 -3520
rect -2664 -4280 -2624 -3560
rect -1904 -4280 -1864 -3560
rect -2664 -4320 -1864 -4280
rect -1252 -3560 -452 -3520
rect -1252 -4280 -1212 -3560
rect -492 -4280 -452 -3560
rect -1252 -4320 -452 -4280
rect 160 -3560 960 -3520
rect 160 -4280 200 -3560
rect 920 -4280 960 -3560
rect 160 -4320 960 -4280
rect 1572 -3560 2372 -3520
rect 1572 -4280 1612 -3560
rect 2332 -4280 2372 -3560
rect 1572 -4320 2372 -4280
<< mimcapcontact >>
rect -2624 3560 -1904 4280
rect -1212 3560 -492 4280
rect 200 3560 920 4280
rect 1612 3560 2332 4280
rect -2624 2440 -1904 3160
rect -1212 2440 -492 3160
rect 200 2440 920 3160
rect 1612 2440 2332 3160
rect -2624 1320 -1904 2040
rect -1212 1320 -492 2040
rect 200 1320 920 2040
rect 1612 1320 2332 2040
rect -2624 200 -1904 920
rect -1212 200 -492 920
rect 200 200 920 920
rect 1612 200 2332 920
rect -2624 -920 -1904 -200
rect -1212 -920 -492 -200
rect 200 -920 920 -200
rect 1612 -920 2332 -200
rect -2624 -2040 -1904 -1320
rect -1212 -2040 -492 -1320
rect 200 -2040 920 -1320
rect 1612 -2040 2332 -1320
rect -2624 -3160 -1904 -2440
rect -1212 -3160 -492 -2440
rect 200 -3160 920 -2440
rect 1612 -3160 2332 -2440
rect -2624 -4280 -1904 -3560
rect -1212 -4280 -492 -3560
rect 200 -4280 920 -3560
rect 1612 -4280 2332 -3560
<< metal4 >>
rect -2316 4281 -2212 4480
rect -1636 4332 -1532 4480
rect -2625 4280 -1903 4281
rect -2625 3560 -2624 4280
rect -1904 3560 -1903 4280
rect -2625 3559 -1903 3560
rect -2316 3161 -2212 3559
rect -1636 3508 -1616 4332
rect -1552 3508 -1532 4332
rect -904 4281 -800 4480
rect -224 4332 -120 4480
rect -1213 4280 -491 4281
rect -1213 3560 -1212 4280
rect -492 3560 -491 4280
rect -1213 3559 -491 3560
rect -1636 3212 -1532 3508
rect -2625 3160 -1903 3161
rect -2625 2440 -2624 3160
rect -1904 2440 -1903 3160
rect -2625 2439 -1903 2440
rect -2316 2041 -2212 2439
rect -1636 2388 -1616 3212
rect -1552 2388 -1532 3212
rect -904 3161 -800 3559
rect -224 3508 -204 4332
rect -140 3508 -120 4332
rect 508 4281 612 4480
rect 1188 4332 1292 4480
rect 199 4280 921 4281
rect 199 3560 200 4280
rect 920 3560 921 4280
rect 199 3559 921 3560
rect -224 3212 -120 3508
rect -1213 3160 -491 3161
rect -1213 2440 -1212 3160
rect -492 2440 -491 3160
rect -1213 2439 -491 2440
rect -1636 2092 -1532 2388
rect -2625 2040 -1903 2041
rect -2625 1320 -2624 2040
rect -1904 1320 -1903 2040
rect -2625 1319 -1903 1320
rect -2316 921 -2212 1319
rect -1636 1268 -1616 2092
rect -1552 1268 -1532 2092
rect -904 2041 -800 2439
rect -224 2388 -204 3212
rect -140 2388 -120 3212
rect 508 3161 612 3559
rect 1188 3508 1208 4332
rect 1272 3508 1292 4332
rect 1920 4281 2024 4480
rect 2600 4332 2704 4480
rect 1611 4280 2333 4281
rect 1611 3560 1612 4280
rect 2332 3560 2333 4280
rect 1611 3559 2333 3560
rect 1188 3212 1292 3508
rect 199 3160 921 3161
rect 199 2440 200 3160
rect 920 2440 921 3160
rect 199 2439 921 2440
rect -224 2092 -120 2388
rect -1213 2040 -491 2041
rect -1213 1320 -1212 2040
rect -492 1320 -491 2040
rect -1213 1319 -491 1320
rect -1636 972 -1532 1268
rect -2625 920 -1903 921
rect -2625 200 -2624 920
rect -1904 200 -1903 920
rect -2625 199 -1903 200
rect -2316 -199 -2212 199
rect -1636 148 -1616 972
rect -1552 148 -1532 972
rect -904 921 -800 1319
rect -224 1268 -204 2092
rect -140 1268 -120 2092
rect 508 2041 612 2439
rect 1188 2388 1208 3212
rect 1272 2388 1292 3212
rect 1920 3161 2024 3559
rect 2600 3508 2620 4332
rect 2684 3508 2704 4332
rect 2600 3212 2704 3508
rect 1611 3160 2333 3161
rect 1611 2440 1612 3160
rect 2332 2440 2333 3160
rect 1611 2439 2333 2440
rect 1188 2092 1292 2388
rect 199 2040 921 2041
rect 199 1320 200 2040
rect 920 1320 921 2040
rect 199 1319 921 1320
rect -224 972 -120 1268
rect -1213 920 -491 921
rect -1213 200 -1212 920
rect -492 200 -491 920
rect -1213 199 -491 200
rect -1636 -148 -1532 148
rect -2625 -200 -1903 -199
rect -2625 -920 -2624 -200
rect -1904 -920 -1903 -200
rect -2625 -921 -1903 -920
rect -2316 -1319 -2212 -921
rect -1636 -972 -1616 -148
rect -1552 -972 -1532 -148
rect -904 -199 -800 199
rect -224 148 -204 972
rect -140 148 -120 972
rect 508 921 612 1319
rect 1188 1268 1208 2092
rect 1272 1268 1292 2092
rect 1920 2041 2024 2439
rect 2600 2388 2620 3212
rect 2684 2388 2704 3212
rect 2600 2092 2704 2388
rect 1611 2040 2333 2041
rect 1611 1320 1612 2040
rect 2332 1320 2333 2040
rect 1611 1319 2333 1320
rect 1188 972 1292 1268
rect 199 920 921 921
rect 199 200 200 920
rect 920 200 921 920
rect 199 199 921 200
rect -224 -148 -120 148
rect -1213 -200 -491 -199
rect -1213 -920 -1212 -200
rect -492 -920 -491 -200
rect -1213 -921 -491 -920
rect -1636 -1268 -1532 -972
rect -2625 -1320 -1903 -1319
rect -2625 -2040 -2624 -1320
rect -1904 -2040 -1903 -1320
rect -2625 -2041 -1903 -2040
rect -2316 -2439 -2212 -2041
rect -1636 -2092 -1616 -1268
rect -1552 -2092 -1532 -1268
rect -904 -1319 -800 -921
rect -224 -972 -204 -148
rect -140 -972 -120 -148
rect 508 -199 612 199
rect 1188 148 1208 972
rect 1272 148 1292 972
rect 1920 921 2024 1319
rect 2600 1268 2620 2092
rect 2684 1268 2704 2092
rect 2600 972 2704 1268
rect 1611 920 2333 921
rect 1611 200 1612 920
rect 2332 200 2333 920
rect 1611 199 2333 200
rect 1188 -148 1292 148
rect 199 -200 921 -199
rect 199 -920 200 -200
rect 920 -920 921 -200
rect 199 -921 921 -920
rect -224 -1268 -120 -972
rect -1213 -1320 -491 -1319
rect -1213 -2040 -1212 -1320
rect -492 -2040 -491 -1320
rect -1213 -2041 -491 -2040
rect -1636 -2388 -1532 -2092
rect -2625 -2440 -1903 -2439
rect -2625 -3160 -2624 -2440
rect -1904 -3160 -1903 -2440
rect -2625 -3161 -1903 -3160
rect -2316 -3559 -2212 -3161
rect -1636 -3212 -1616 -2388
rect -1552 -3212 -1532 -2388
rect -904 -2439 -800 -2041
rect -224 -2092 -204 -1268
rect -140 -2092 -120 -1268
rect 508 -1319 612 -921
rect 1188 -972 1208 -148
rect 1272 -972 1292 -148
rect 1920 -199 2024 199
rect 2600 148 2620 972
rect 2684 148 2704 972
rect 2600 -148 2704 148
rect 1611 -200 2333 -199
rect 1611 -920 1612 -200
rect 2332 -920 2333 -200
rect 1611 -921 2333 -920
rect 1188 -1268 1292 -972
rect 199 -1320 921 -1319
rect 199 -2040 200 -1320
rect 920 -2040 921 -1320
rect 199 -2041 921 -2040
rect -224 -2388 -120 -2092
rect -1213 -2440 -491 -2439
rect -1213 -3160 -1212 -2440
rect -492 -3160 -491 -2440
rect -1213 -3161 -491 -3160
rect -1636 -3508 -1532 -3212
rect -2625 -3560 -1903 -3559
rect -2625 -4280 -2624 -3560
rect -1904 -4280 -1903 -3560
rect -2625 -4281 -1903 -4280
rect -2316 -4480 -2212 -4281
rect -1636 -4332 -1616 -3508
rect -1552 -4332 -1532 -3508
rect -904 -3559 -800 -3161
rect -224 -3212 -204 -2388
rect -140 -3212 -120 -2388
rect 508 -2439 612 -2041
rect 1188 -2092 1208 -1268
rect 1272 -2092 1292 -1268
rect 1920 -1319 2024 -921
rect 2600 -972 2620 -148
rect 2684 -972 2704 -148
rect 2600 -1268 2704 -972
rect 1611 -1320 2333 -1319
rect 1611 -2040 1612 -1320
rect 2332 -2040 2333 -1320
rect 1611 -2041 2333 -2040
rect 1188 -2388 1292 -2092
rect 199 -2440 921 -2439
rect 199 -3160 200 -2440
rect 920 -3160 921 -2440
rect 199 -3161 921 -3160
rect -224 -3508 -120 -3212
rect -1213 -3560 -491 -3559
rect -1213 -4280 -1212 -3560
rect -492 -4280 -491 -3560
rect -1213 -4281 -491 -4280
rect -1636 -4480 -1532 -4332
rect -904 -4480 -800 -4281
rect -224 -4332 -204 -3508
rect -140 -4332 -120 -3508
rect 508 -3559 612 -3161
rect 1188 -3212 1208 -2388
rect 1272 -3212 1292 -2388
rect 1920 -2439 2024 -2041
rect 2600 -2092 2620 -1268
rect 2684 -2092 2704 -1268
rect 2600 -2388 2704 -2092
rect 1611 -2440 2333 -2439
rect 1611 -3160 1612 -2440
rect 2332 -3160 2333 -2440
rect 1611 -3161 2333 -3160
rect 1188 -3508 1292 -3212
rect 199 -3560 921 -3559
rect 199 -4280 200 -3560
rect 920 -4280 921 -3560
rect 199 -4281 921 -4280
rect -224 -4480 -120 -4332
rect 508 -4480 612 -4281
rect 1188 -4332 1208 -3508
rect 1272 -4332 1292 -3508
rect 1920 -3559 2024 -3161
rect 2600 -3212 2620 -2388
rect 2684 -3212 2704 -2388
rect 2600 -3508 2704 -3212
rect 1611 -3560 2333 -3559
rect 1611 -4280 1612 -3560
rect 2332 -4280 2333 -3560
rect 1611 -4281 2333 -4280
rect 1188 -4480 1292 -4332
rect 1920 -4480 2024 -4281
rect 2600 -4332 2620 -3508
rect 2684 -4332 2704 -3508
rect 2600 -4480 2704 -4332
<< properties >>
string FIXED_BBOX 1532 3480 2412 4360
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 4.0 l 4.0 val 35.04 carea 2.00 cperi 0.19 nx 4 ny 8 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
