../mag/x10b_adc.pex.spice