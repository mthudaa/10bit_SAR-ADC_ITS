magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect 238 1527 272 1561
rect 306 1527 344 1561
rect 378 1527 416 1561
rect 450 1527 488 1561
rect 522 1527 560 1561
rect 594 1527 632 1561
rect 666 1527 704 1561
rect 738 1527 776 1561
rect 810 1527 848 1561
rect 882 1527 920 1561
rect 954 1527 992 1561
rect 1026 1527 1064 1561
rect 1098 1527 1136 1561
rect 1170 1527 1208 1561
rect 1242 1527 1280 1561
rect 1314 1527 1352 1561
rect 1386 1527 1424 1561
rect 1458 1527 1496 1561
rect 1530 1527 1568 1561
rect 1602 1527 1640 1561
rect 1674 1527 1712 1561
rect 1746 1527 1784 1561
rect 1818 1527 1856 1561
rect 1890 1527 1928 1561
rect 1962 1527 1996 1561
rect 238 -123 268 -89
rect 302 -123 340 -89
rect 374 -123 412 -89
rect 446 -123 484 -89
rect 518 -123 556 -89
rect 590 -123 628 -89
rect 662 -123 700 -89
rect 734 -123 772 -89
rect 806 -123 844 -89
rect 878 -123 916 -89
rect 950 -123 988 -89
rect 1022 -123 1060 -89
rect 1094 -123 1124 -89
<< viali >>
rect 272 1527 306 1561
rect 344 1527 378 1561
rect 416 1527 450 1561
rect 488 1527 522 1561
rect 560 1527 594 1561
rect 632 1527 666 1561
rect 704 1527 738 1561
rect 776 1527 810 1561
rect 848 1527 882 1561
rect 920 1527 954 1561
rect 992 1527 1026 1561
rect 1064 1527 1098 1561
rect 1136 1527 1170 1561
rect 1208 1527 1242 1561
rect 1280 1527 1314 1561
rect 1352 1527 1386 1561
rect 1424 1527 1458 1561
rect 1496 1527 1530 1561
rect 1568 1527 1602 1561
rect 1640 1527 1674 1561
rect 1712 1527 1746 1561
rect 1784 1527 1818 1561
rect 1856 1527 1890 1561
rect 1928 1527 1962 1561
rect 268 -123 302 -89
rect 340 -123 374 -89
rect 412 -123 446 -89
rect 484 -123 518 -89
rect 556 -123 590 -89
rect 628 -123 662 -89
rect 700 -123 734 -89
rect 772 -123 806 -89
rect 844 -123 878 -89
rect 916 -123 950 -89
rect 988 -123 1022 -89
rect 1060 -123 1094 -89
<< metal1 >>
rect 106 1561 2128 1597
rect 106 1527 272 1561
rect 306 1527 344 1561
rect 378 1527 416 1561
rect 450 1527 488 1561
rect 522 1527 560 1561
rect 594 1527 632 1561
rect 666 1527 704 1561
rect 738 1527 776 1561
rect 810 1527 848 1561
rect 882 1527 920 1561
rect 954 1527 992 1561
rect 1026 1527 1064 1561
rect 1098 1527 1136 1561
rect 1170 1527 1208 1561
rect 1242 1527 1280 1561
rect 1314 1527 1352 1561
rect 1386 1527 1424 1561
rect 1458 1527 1496 1561
rect 1530 1527 1568 1561
rect 1602 1527 1640 1561
rect 1674 1527 1712 1561
rect 1746 1527 1784 1561
rect 1818 1527 1856 1561
rect 1890 1527 1928 1561
rect 1962 1527 2128 1561
rect 106 1521 2128 1527
rect 325 1447 1909 1521
rect 106 1377 283 1401
rect 106 1325 176 1377
rect 228 1325 283 1377
rect 106 1301 283 1325
rect 325 1061 1909 1255
rect 106 915 284 1015
rect 106 570 2128 869
rect 106 423 284 523
rect 316 183 1046 377
rect 166 113 284 137
rect 166 61 176 113
rect 228 61 284 113
rect 166 37 284 61
rect 316 -83 1046 -9
rect 106 -89 2128 -83
rect 106 -123 268 -89
rect 302 -123 340 -89
rect 374 -123 412 -89
rect 446 -123 484 -89
rect 518 -123 556 -89
rect 590 -123 628 -89
rect 662 -123 700 -89
rect 734 -123 772 -89
rect 806 -123 844 -89
rect 878 -123 916 -89
rect 950 -123 988 -89
rect 1022 -123 1060 -89
rect 1094 -123 2128 -89
rect 106 -159 2128 -123
<< via1 >>
rect 176 1325 228 1377
rect 176 61 228 113
<< metal2 >>
rect 176 1377 228 1411
rect 176 113 228 1325
rect 176 27 228 61
use sky130_fd_pr__nfet_01v8_KT5VMN  sky130_fd_pr__nfet_01v8_KT5VMN_0
timestamp 1750100919
transform 0 1 681 -1 0 87
box -236 -565 236 565
use sky130_fd_pr__pfet_01v8_NMYCWJ  sky130_fd_pr__pfet_01v8_NMYCWJ_0
timestamp 1750100919
transform 0 1 1117 -1 0 965
box -246 -1011 246 1011
use sky130_fd_pr__pfet_01v8_NMYCWJ  XM1
timestamp 1750100919
transform 0 1 1117 -1 0 1351
box -246 -1011 246 1011
use sky130_fd_pr__nfet_01v8_KT5VMN  XM3
timestamp 1750100919
transform 0 1 681 -1 0 473
box -236 -565 236 565
<< labels >>
flabel metal1 s 106 1521 238 1597 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 106 1301 176 1401 0 FreeSans 500 0 0 0 IN
port 2 nsew
flabel metal1 s 106 915 284 1015 0 FreeSans 500 0 0 0 CKB
port 3 nsew
flabel metal1 s 106 423 284 523 0 FreeSans 500 0 0 0 CK
port 4 nsew
flabel metal1 s 106 -159 238 -83 0 FreeSans 500 0 0 0 VSS
port 5 nsew
flabel metal1 s 1962 666 2074 747 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
