magic
tech sky130A
magscale 1 2
timestamp 1748800002
<< metal1 >>
rect -228 1302 -218 1400
rect -118 1302 61 1400
rect -1628 1168 -1618 1228
rect -1518 1168 42 1228
rect -628 1017 -618 1077
rect -518 1017 42 1077
rect -828 841 -818 901
rect -718 841 51 901
rect -428 636 -418 734
rect -318 636 116 734
rect -1028 293 -1018 353
rect -918 293 45 353
rect -1228 138 -1218 198
rect -1118 138 44 198
rect -228 -106 -218 68
rect -118 -106 91 68
rect -628 -712 -618 -612
rect -518 -712 67 -612
rect 8552 -1058 13463 -758
rect 13563 -1058 13573 -758
rect -828 -1204 -818 -1104
rect -718 -1204 -18 -1104
rect -1828 -1590 -1818 -1490
rect -1718 -1590 49 -1490
rect -428 -1862 -418 -1710
rect -318 -1862 59 -1710
rect 13453 -1902 13463 -1868
rect -27 -2078 -17 -1986
rect 83 -2078 93 -1986
rect 4476 -2162 4510 -1902
rect 13226 -1936 13463 -1902
rect 13453 -1970 13463 -1936
rect 13563 -1970 13573 -1868
rect 13253 -2078 13263 -1986
rect 13363 -2078 13373 -1986
rect -228 -2354 -218 -2202
rect -118 -2354 57 -2202
rect 13453 -2394 13463 -2360
rect 13218 -2428 13463 -2394
rect 13453 -2462 13463 -2428
rect 13563 -2462 13573 -2360
rect -1228 -2570 -1218 -2478
rect -1118 -2570 -17 -2478
rect 83 -2570 93 -2478
rect 13253 -2570 13263 -2478
rect 13363 -2570 13373 -2478
rect -1428 -2688 -1418 -2586
rect -1318 -2620 -1308 -2586
rect -1318 -2654 126 -2620
rect -1318 -2688 -1308 -2654
rect -428 -2846 -418 -2694
rect -318 -2846 51 -2694
rect -27 -3062 -17 -2970
rect 83 -3062 93 -2970
rect -1428 -3180 -1418 -3078
rect -1318 -3112 -1308 -3078
rect -1318 -3146 109 -3112
rect 4476 -3146 4510 -2886
rect 13253 -3062 13263 -2970
rect 13363 -3062 13373 -2970
rect -1318 -3180 -1308 -3146
rect -228 -3262 -218 -3186
rect -118 -3262 84 -3186
<< via1 >>
rect -218 1302 -118 1400
rect -1618 1168 -1518 1228
rect -618 1017 -518 1077
rect -818 841 -718 901
rect -418 636 -318 734
rect -1018 293 -918 353
rect -1218 138 -1118 198
rect -218 -106 -118 68
rect -618 -712 -518 -612
rect 13463 -1058 13563 -758
rect -818 -1204 -718 -1104
rect -1818 -1590 -1718 -1490
rect -418 -1862 -318 -1710
rect -17 -2078 83 -1986
rect 13463 -1970 13563 -1868
rect 13263 -2078 13363 -1986
rect -218 -2354 -118 -2202
rect 13463 -2462 13563 -2360
rect -1218 -2570 -1118 -2478
rect -17 -2570 83 -2478
rect 13263 -2570 13363 -2478
rect -1418 -2688 -1318 -2586
rect -418 -2846 -318 -2694
rect -17 -3062 83 -2970
rect -1418 -3180 -1318 -3078
rect 13263 -3062 13363 -2970
rect -218 -3262 -118 -3186
<< metal2 >>
rect -218 1400 -118 1410
rect -1818 -1490 -1718 1400
rect -1818 -3272 -1718 -1590
rect -1618 1228 -1518 1400
rect -1618 -3272 -1518 1168
rect -1418 -2586 -1318 1400
rect -1418 -3078 -1318 -2688
rect -1418 -3272 -1318 -3180
rect -1218 198 -1118 1400
rect -1218 -2478 -1118 138
rect -1218 -3272 -1118 -2570
rect -1018 353 -918 1400
rect -1018 -1986 -918 293
rect -1018 -3272 -918 -2078
rect -818 901 -718 1400
rect -818 -1104 -718 841
rect -818 -3272 -718 -1204
rect -618 1077 -518 1400
rect -618 -612 -518 1017
rect -618 -3272 -518 -712
rect -418 734 -318 1400
rect -418 -1710 -318 636
rect -418 -2694 -318 -1862
rect -418 -3272 -318 -2846
rect -218 68 -118 1302
rect -218 -2202 -118 -106
rect 13463 -758 13563 -748
rect 13463 -1868 13563 -1058
rect -218 -3186 -118 -2354
rect -17 -1986 83 -1976
rect -17 -2478 83 -2078
rect -17 -2970 83 -2570
rect -17 -3072 83 -3062
rect 13263 -1986 13363 -1976
rect 13263 -2478 13363 -2078
rect 13263 -2970 13363 -2570
rect 13263 -3072 13363 -3062
rect 13463 -2360 13563 -1970
rect 13463 -3262 13563 -2462
rect -218 -3272 -118 -3262
<< via2 >>
rect -1018 -2078 -918 -1986
rect 13263 -2078 13363 -1986
<< metal3 >>
rect -1028 -1986 -908 -1981
rect 13253 -1986 13373 -1981
rect -1028 -2078 -1018 -1986
rect -918 -2078 13263 -1986
rect 13363 -2078 13373 -1986
rect -1028 -2083 -908 -2078
rect 13253 -2083 13373 -2078
use dac_sw_1  dac_sw_1_0
timestamp 1746262095
transform 1 0 -124 0 -1 -189
box 106 -159 8976 1597
use nooverlap_clk  nooverlap_clk_0
timestamp 1748785634
transform -1 0 2909 0 1 4745
box -701 -4775 2927 -3345
use tg_sw_1  tg_sw_1_0
timestamp 1748683470
transform -1 0 13310 0 1 -2225
box -53 -53 13327 439
use tg_sw_1  tg_sw_1_1
timestamp 1748683470
transform 1 0 36 0 -1 -2331
box -53 -53 13327 439
use tg_sw_1  tg_sw_1_2
timestamp 1748683470
transform -1 0 13310 0 1 -3209
box -53 -53 13327 439
<< labels >>
flabel metal1 13244 -973 13344 -839 0 FreeSans 400 0 0 0 DAC_OUT
port 6 nsew
flabel metal2 -182 -393 -142 -353 0 FreeSans 480 0 0 0 VSSA
port 8 nsew
flabel metal2 -393 -382 -353 -342 0 FreeSans 480 0 0 0 VDDA
port 9 nsew
flabel metal2 -1384 -382 -1344 -342 0 FreeSans 480 0 0 0 VCM
port 10 nsew
flabel metal2 -1593 -388 -1553 -348 0 FreeSans 480 0 0 0 CKI
port 11 nsew
flabel metal2 -1786 -378 -1746 -338 0 FreeSans 480 0 0 0 BI
port 13 nsew
<< end >>
