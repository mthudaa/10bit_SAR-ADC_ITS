magic
tech sky130A
magscale 1 2
timestamp 1749411235
<< metal1 >>
rect -224 2900 -214 2996
rect -118 2900 5318 2996
rect 5414 2900 5424 2996
rect -32 2708 -22 2804
rect 74 2708 2306 2804
rect 2404 2708 5126 2804
rect 5222 2708 5232 2804
rect 2195 2516 2306 2612
rect 2404 2516 2414 2612
rect 368 2423 378 2475
rect 430 2466 440 2475
rect 430 2432 609 2466
rect 430 2423 440 2432
rect 2296 2301 2306 2399
rect 2404 2301 2414 2399
rect 2095 1888 2410 1940
rect 160 1379 170 1388
rect -214 1345 170 1379
rect 160 1336 170 1345
rect 222 1379 232 1388
rect 222 1345 613 1379
rect 222 1336 232 1345
rect 264 1305 274 1314
rect -214 1271 274 1305
rect 264 1262 274 1271
rect 326 1305 336 1314
rect 326 1271 636 1305
rect 326 1262 336 1271
rect -224 1132 -214 1228
rect -118 1132 496 1228
rect 2210 1132 2306 1228
rect 4990 1132 5318 1228
rect 5414 1132 5424 1228
rect 368 1089 378 1098
rect -214 1055 378 1089
rect 368 1046 378 1055
rect 430 1089 440 1098
rect 430 1055 671 1089
rect 430 1046 440 1055
rect 160 972 170 1024
rect 222 1015 232 1024
rect 222 981 624 1015
rect 222 972 232 981
rect 4983 888 5414 928
rect 4984 676 5414 716
rect 4990 597 5414 637
rect 2095 406 2519 458
rect 2296 -39 2306 59
rect 2404 -39 2414 59
rect 264 -115 274 -63
rect 326 -72 336 -63
rect 326 -106 637 -72
rect 326 -115 336 -106
rect 2204 -252 2306 -156
rect 2404 -252 2414 -156
rect -32 -444 -22 -348
rect 74 -444 2306 -348
rect 2404 -444 3552 -348
rect 3648 -444 5126 -348
rect 5222 -444 5232 -348
rect -224 -636 -214 -540
rect -118 -636 5318 -540
rect 5414 -636 5424 -540
<< via1 >>
rect -214 2900 -118 2996
rect 5318 2900 5414 2996
rect -22 2708 74 2804
rect 2306 2708 2404 2804
rect 5126 2708 5222 2804
rect 2306 2516 2404 2612
rect 378 2423 430 2475
rect 2306 2301 2404 2399
rect 170 1336 222 1388
rect 274 1262 326 1314
rect -214 1132 -118 1228
rect 5318 1132 5414 1228
rect 378 1046 430 1098
rect 170 972 222 1024
rect 2306 -39 2404 59
rect 274 -115 326 -63
rect 2306 -252 2404 -156
rect -22 -444 74 -348
rect 2306 -444 2404 -348
rect 3552 -444 3648 -348
rect 5126 -444 5222 -348
rect -214 -636 -118 -540
rect 5318 -636 5414 -540
<< metal2 >>
rect -214 2996 -118 3006
rect -214 1228 -118 2900
rect 5318 2996 5414 3006
rect -214 -540 -118 1132
rect -22 2804 74 2814
rect -22 -348 74 2708
rect 2306 2804 2404 2814
rect 2306 2612 2404 2708
rect 378 2475 430 2485
rect 170 1388 222 1398
rect 170 1024 222 1336
rect 170 962 222 972
rect 274 1314 326 1324
rect 274 -63 326 1262
rect 378 1098 430 2423
rect 2306 2399 2404 2516
rect 2306 2291 2404 2301
rect 5126 2804 5222 2814
rect 378 1036 430 1046
rect 274 -125 326 -115
rect 2306 59 2404 69
rect -22 -454 74 -444
rect 2306 -156 2404 -39
rect 2306 -348 2404 -252
rect 2306 -454 2404 -444
rect 3552 -348 3648 210
rect 3552 -454 3648 -444
rect 5126 -348 5222 2708
rect 5126 -454 5222 -444
rect 5318 1228 5414 2900
rect -214 -646 -118 -636
rect 5318 -540 5414 1132
rect 5318 -646 5414 -636
use delay_gate_ori  delay_gate_ori_0
timestamp 1749411235
transform 1 0 1371 0 -1 2130
box -875 -482 853 998
use delay_gate_ori  delay_gate_ori_1
timestamp 1749411235
transform 1 0 1371 0 1 230
box -875 -482 853 998
use phase_detector  phase_detector_0
timestamp 1749411235
transform 1 0 2324 0 1 -47
box -28 -2 2706 2456
<< labels >>
flabel metal1 412 2934 442 2964 0 FreeSans 400 0 0 0 VDD
port 0 nsew
flabel metal1 392 2748 422 2778 0 FreeSans 400 0 0 0 VSS
port 1 nsew
flabel metal1 -93 1271 -59 1305 0 FreeSans 400 0 0 0 VINP
port 3 nsew
flabel metal1 -92 1055 -58 1089 0 FreeSans 400 0 0 0 VINN
port 4 nsew
flabel metal1 5245 888 5285 928 0 FreeSans 400 0 0 0 RDY
port 5 nsew
flabel metal1 5253 676 5293 716 0 FreeSans 400 0 0 0 OUTP
port 6 nsew
flabel metal1 5249 597 5289 637 0 FreeSans 400 0 0 0 OUTN
port 8 nsew
flabel metal1 -103 1345 -69 1379 0 FreeSans 400 0 0 0 CLK
port 10 nsew
<< end >>
