magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect -17 369 9 403
rect 43 369 81 403
rect 115 369 153 403
rect 187 369 225 403
rect 259 369 297 403
rect 331 369 369 403
rect 403 369 441 403
rect 475 369 513 403
rect 547 369 585 403
rect 619 369 657 403
rect 691 369 729 403
rect 763 369 801 403
rect 835 369 873 403
rect 907 369 945 403
rect 979 369 1017 403
rect 1051 369 1089 403
rect 1123 369 1161 403
rect 1195 369 1233 403
rect 1267 369 1305 403
rect 1339 369 1377 403
rect 1411 369 1449 403
rect 1483 369 1521 403
rect 1555 369 1593 403
rect 1627 369 1665 403
rect 1699 369 1737 403
rect 1771 369 1809 403
rect 1843 369 1881 403
rect 1915 369 1953 403
rect 1987 369 2025 403
rect 2059 369 2097 403
rect 2131 369 2169 403
rect 2203 369 2241 403
rect 2275 369 2313 403
rect 2347 369 2385 403
rect 2419 369 2457 403
rect 2491 369 2529 403
rect 2563 369 2601 403
rect 2635 369 2673 403
rect 2707 369 2745 403
rect 2779 369 2817 403
rect 2851 369 2889 403
rect 2923 369 2961 403
rect 2995 369 3033 403
rect 3067 369 3105 403
rect 3139 369 3177 403
rect 3211 369 3249 403
rect 3283 369 3321 403
rect 3355 369 3393 403
rect 3427 369 3465 403
rect 3499 369 3537 403
rect 3571 369 3609 403
rect 3643 369 3681 403
rect 3715 369 3753 403
rect 3787 369 3825 403
rect 3859 369 3897 403
rect 3931 369 3969 403
rect 4003 369 4041 403
rect 4075 369 4113 403
rect 4147 369 4185 403
rect 4219 369 4257 403
rect 4291 369 4329 403
rect 4363 369 4401 403
rect 4435 369 4473 403
rect 4507 369 4545 403
rect 4579 369 4617 403
rect 4651 369 4689 403
rect 4723 369 4761 403
rect 4795 369 4833 403
rect 4867 369 4905 403
rect 4939 369 4977 403
rect 5011 369 5049 403
rect 5083 369 5121 403
rect 5155 369 5193 403
rect 5227 369 5265 403
rect 5299 369 5337 403
rect 5371 369 5409 403
rect 5443 369 5481 403
rect 5515 369 5553 403
rect 5587 369 5625 403
rect 5659 369 5697 403
rect 5731 369 5769 403
rect 5803 369 5841 403
rect 5875 369 5913 403
rect 5947 369 5985 403
rect 6019 369 6057 403
rect 6091 369 6129 403
rect 6163 369 6201 403
rect 6235 369 6273 403
rect 6307 369 6345 403
rect 6379 369 6417 403
rect 6451 369 6489 403
rect 6523 369 6561 403
rect 6595 369 6633 403
rect 6667 369 6705 403
rect 6739 369 6777 403
rect 6811 369 6849 403
rect 6883 369 6921 403
rect 6955 369 6993 403
rect 7027 369 7065 403
rect 7099 369 7137 403
rect 7171 369 7209 403
rect 7243 369 7281 403
rect 7315 369 7353 403
rect 7387 369 7425 403
rect 7459 369 7497 403
rect 7531 369 7569 403
rect 7603 369 7641 403
rect 7675 369 7713 403
rect 7747 369 7785 403
rect 7819 369 7857 403
rect 7891 369 7929 403
rect 7963 369 8001 403
rect 8035 369 8073 403
rect 8107 369 8145 403
rect 8179 369 8217 403
rect 8251 369 8289 403
rect 8323 369 8361 403
rect 8395 369 8433 403
rect 8467 369 8505 403
rect 8539 369 8577 403
rect 8611 369 8649 403
rect 8683 369 8721 403
rect 8755 369 8781 403
rect 8853 -17 8859 17
rect 8893 -17 8931 17
rect 8965 -17 9003 17
rect 9037 -17 9075 17
rect 9109 -17 9147 17
rect 9181 -17 9219 17
rect 9253 -17 9291 17
rect 9325 -17 9363 17
rect 9397 -17 9435 17
rect 9469 -17 9507 17
rect 9541 -17 9579 17
rect 9613 -17 9651 17
rect 9685 -17 9723 17
rect 9757 -17 9795 17
rect 9829 -17 9867 17
rect 9901 -17 9939 17
rect 9973 -17 10011 17
rect 10045 -17 10083 17
rect 10117 -17 10155 17
rect 10189 -17 10227 17
rect 10261 -17 10299 17
rect 10333 -17 10371 17
rect 10405 -17 10443 17
rect 10477 -17 10515 17
rect 10549 -17 10587 17
rect 10621 -17 10659 17
rect 10693 -17 10731 17
rect 10765 -17 10803 17
rect 10837 -17 10875 17
rect 10909 -17 10947 17
rect 10981 -17 11019 17
rect 11053 -17 11091 17
rect 11125 -17 11163 17
rect 11197 -17 11235 17
rect 11269 -17 11307 17
rect 11341 -17 11379 17
rect 11413 -17 11451 17
rect 11485 -17 11523 17
rect 11557 -17 11595 17
rect 11629 -17 11667 17
rect 11701 -17 11739 17
rect 11773 -17 11811 17
rect 11845 -17 11883 17
rect 11917 -17 11955 17
rect 11989 -17 12027 17
rect 12061 -17 12099 17
rect 12133 -17 12171 17
rect 12205 -17 12243 17
rect 12277 -17 12315 17
rect 12349 -17 12387 17
rect 12421 -17 12459 17
rect 12493 -17 12531 17
rect 12565 -17 12603 17
rect 12637 -17 12675 17
rect 12709 -17 12747 17
rect 12781 -17 12819 17
rect 12853 -17 12891 17
rect 12925 -17 12963 17
rect 12997 -17 13035 17
rect 13069 -17 13107 17
rect 13141 -17 13179 17
rect 13213 -17 13251 17
rect 13285 -17 13291 17
<< viali >>
rect 9 369 43 403
rect 81 369 115 403
rect 153 369 187 403
rect 225 369 259 403
rect 297 369 331 403
rect 369 369 403 403
rect 441 369 475 403
rect 513 369 547 403
rect 585 369 619 403
rect 657 369 691 403
rect 729 369 763 403
rect 801 369 835 403
rect 873 369 907 403
rect 945 369 979 403
rect 1017 369 1051 403
rect 1089 369 1123 403
rect 1161 369 1195 403
rect 1233 369 1267 403
rect 1305 369 1339 403
rect 1377 369 1411 403
rect 1449 369 1483 403
rect 1521 369 1555 403
rect 1593 369 1627 403
rect 1665 369 1699 403
rect 1737 369 1771 403
rect 1809 369 1843 403
rect 1881 369 1915 403
rect 1953 369 1987 403
rect 2025 369 2059 403
rect 2097 369 2131 403
rect 2169 369 2203 403
rect 2241 369 2275 403
rect 2313 369 2347 403
rect 2385 369 2419 403
rect 2457 369 2491 403
rect 2529 369 2563 403
rect 2601 369 2635 403
rect 2673 369 2707 403
rect 2745 369 2779 403
rect 2817 369 2851 403
rect 2889 369 2923 403
rect 2961 369 2995 403
rect 3033 369 3067 403
rect 3105 369 3139 403
rect 3177 369 3211 403
rect 3249 369 3283 403
rect 3321 369 3355 403
rect 3393 369 3427 403
rect 3465 369 3499 403
rect 3537 369 3571 403
rect 3609 369 3643 403
rect 3681 369 3715 403
rect 3753 369 3787 403
rect 3825 369 3859 403
rect 3897 369 3931 403
rect 3969 369 4003 403
rect 4041 369 4075 403
rect 4113 369 4147 403
rect 4185 369 4219 403
rect 4257 369 4291 403
rect 4329 369 4363 403
rect 4401 369 4435 403
rect 4473 369 4507 403
rect 4545 369 4579 403
rect 4617 369 4651 403
rect 4689 369 4723 403
rect 4761 369 4795 403
rect 4833 369 4867 403
rect 4905 369 4939 403
rect 4977 369 5011 403
rect 5049 369 5083 403
rect 5121 369 5155 403
rect 5193 369 5227 403
rect 5265 369 5299 403
rect 5337 369 5371 403
rect 5409 369 5443 403
rect 5481 369 5515 403
rect 5553 369 5587 403
rect 5625 369 5659 403
rect 5697 369 5731 403
rect 5769 369 5803 403
rect 5841 369 5875 403
rect 5913 369 5947 403
rect 5985 369 6019 403
rect 6057 369 6091 403
rect 6129 369 6163 403
rect 6201 369 6235 403
rect 6273 369 6307 403
rect 6345 369 6379 403
rect 6417 369 6451 403
rect 6489 369 6523 403
rect 6561 369 6595 403
rect 6633 369 6667 403
rect 6705 369 6739 403
rect 6777 369 6811 403
rect 6849 369 6883 403
rect 6921 369 6955 403
rect 6993 369 7027 403
rect 7065 369 7099 403
rect 7137 369 7171 403
rect 7209 369 7243 403
rect 7281 369 7315 403
rect 7353 369 7387 403
rect 7425 369 7459 403
rect 7497 369 7531 403
rect 7569 369 7603 403
rect 7641 369 7675 403
rect 7713 369 7747 403
rect 7785 369 7819 403
rect 7857 369 7891 403
rect 7929 369 7963 403
rect 8001 369 8035 403
rect 8073 369 8107 403
rect 8145 369 8179 403
rect 8217 369 8251 403
rect 8289 369 8323 403
rect 8361 369 8395 403
rect 8433 369 8467 403
rect 8505 369 8539 403
rect 8577 369 8611 403
rect 8649 369 8683 403
rect 8721 369 8755 403
rect 8859 -17 8893 17
rect 8931 -17 8965 17
rect 9003 -17 9037 17
rect 9075 -17 9109 17
rect 9147 -17 9181 17
rect 9219 -17 9253 17
rect 9291 -17 9325 17
rect 9363 -17 9397 17
rect 9435 -17 9469 17
rect 9507 -17 9541 17
rect 9579 -17 9613 17
rect 9651 -17 9685 17
rect 9723 -17 9757 17
rect 9795 -17 9829 17
rect 9867 -17 9901 17
rect 9939 -17 9973 17
rect 10011 -17 10045 17
rect 10083 -17 10117 17
rect 10155 -17 10189 17
rect 10227 -17 10261 17
rect 10299 -17 10333 17
rect 10371 -17 10405 17
rect 10443 -17 10477 17
rect 10515 -17 10549 17
rect 10587 -17 10621 17
rect 10659 -17 10693 17
rect 10731 -17 10765 17
rect 10803 -17 10837 17
rect 10875 -17 10909 17
rect 10947 -17 10981 17
rect 11019 -17 11053 17
rect 11091 -17 11125 17
rect 11163 -17 11197 17
rect 11235 -17 11269 17
rect 11307 -17 11341 17
rect 11379 -17 11413 17
rect 11451 -17 11485 17
rect 11523 -17 11557 17
rect 11595 -17 11629 17
rect 11667 -17 11701 17
rect 11739 -17 11773 17
rect 11811 -17 11845 17
rect 11883 -17 11917 17
rect 11955 -17 11989 17
rect 12027 -17 12061 17
rect 12099 -17 12133 17
rect 12171 -17 12205 17
rect 12243 -17 12277 17
rect 12315 -17 12349 17
rect 12387 -17 12421 17
rect 12459 -17 12493 17
rect 12531 -17 12565 17
rect 12603 -17 12637 17
rect 12675 -17 12709 17
rect 12747 -17 12781 17
rect 12819 -17 12853 17
rect 12891 -17 12925 17
rect 12963 -17 12997 17
rect 13035 -17 13069 17
rect 13107 -17 13141 17
rect 13179 -17 13213 17
rect 13251 -17 13285 17
<< metal1 >>
rect -53 403 13327 439
rect -53 369 9 403
rect 43 369 81 403
rect 115 369 153 403
rect 187 369 225 403
rect 259 369 297 403
rect 331 369 369 403
rect 403 369 441 403
rect 475 369 513 403
rect 547 369 585 403
rect 619 369 657 403
rect 691 369 729 403
rect 763 369 801 403
rect 835 369 873 403
rect 907 369 945 403
rect 979 369 1017 403
rect 1051 369 1089 403
rect 1123 369 1161 403
rect 1195 369 1233 403
rect 1267 369 1305 403
rect 1339 369 1377 403
rect 1411 369 1449 403
rect 1483 369 1521 403
rect 1555 369 1593 403
rect 1627 369 1665 403
rect 1699 369 1737 403
rect 1771 369 1809 403
rect 1843 369 1881 403
rect 1915 369 1953 403
rect 1987 369 2025 403
rect 2059 369 2097 403
rect 2131 369 2169 403
rect 2203 369 2241 403
rect 2275 369 2313 403
rect 2347 369 2385 403
rect 2419 369 2457 403
rect 2491 369 2529 403
rect 2563 369 2601 403
rect 2635 369 2673 403
rect 2707 369 2745 403
rect 2779 369 2817 403
rect 2851 369 2889 403
rect 2923 369 2961 403
rect 2995 369 3033 403
rect 3067 369 3105 403
rect 3139 369 3177 403
rect 3211 369 3249 403
rect 3283 369 3321 403
rect 3355 369 3393 403
rect 3427 369 3465 403
rect 3499 369 3537 403
rect 3571 369 3609 403
rect 3643 369 3681 403
rect 3715 369 3753 403
rect 3787 369 3825 403
rect 3859 369 3897 403
rect 3931 369 3969 403
rect 4003 369 4041 403
rect 4075 369 4113 403
rect 4147 369 4185 403
rect 4219 369 4257 403
rect 4291 369 4329 403
rect 4363 369 4401 403
rect 4435 369 4473 403
rect 4507 369 4545 403
rect 4579 369 4617 403
rect 4651 369 4689 403
rect 4723 369 4761 403
rect 4795 369 4833 403
rect 4867 369 4905 403
rect 4939 369 4977 403
rect 5011 369 5049 403
rect 5083 369 5121 403
rect 5155 369 5193 403
rect 5227 369 5265 403
rect 5299 369 5337 403
rect 5371 369 5409 403
rect 5443 369 5481 403
rect 5515 369 5553 403
rect 5587 369 5625 403
rect 5659 369 5697 403
rect 5731 369 5769 403
rect 5803 369 5841 403
rect 5875 369 5913 403
rect 5947 369 5985 403
rect 6019 369 6057 403
rect 6091 369 6129 403
rect 6163 369 6201 403
rect 6235 369 6273 403
rect 6307 369 6345 403
rect 6379 369 6417 403
rect 6451 369 6489 403
rect 6523 369 6561 403
rect 6595 369 6633 403
rect 6667 369 6705 403
rect 6739 369 6777 403
rect 6811 369 6849 403
rect 6883 369 6921 403
rect 6955 369 6993 403
rect 7027 369 7065 403
rect 7099 369 7137 403
rect 7171 369 7209 403
rect 7243 369 7281 403
rect 7315 369 7353 403
rect 7387 369 7425 403
rect 7459 369 7497 403
rect 7531 369 7569 403
rect 7603 369 7641 403
rect 7675 369 7713 403
rect 7747 369 7785 403
rect 7819 369 7857 403
rect 7891 369 7929 403
rect 7963 369 8001 403
rect 8035 369 8073 403
rect 8107 369 8145 403
rect 8179 369 8217 403
rect 8251 369 8289 403
rect 8323 369 8361 403
rect 8395 369 8433 403
rect 8467 369 8505 403
rect 8539 369 8577 403
rect 8611 369 8649 403
rect 8683 369 8721 403
rect 8755 369 13327 403
rect -53 363 13327 369
rect -53 289 13117 323
rect -53 147 125 239
rect 13149 147 13327 239
rect 166 63 13327 97
rect -53 17 13327 23
rect -53 -17 8859 17
rect 8893 -17 8931 17
rect 8965 -17 9003 17
rect 9037 -17 9075 17
rect 9109 -17 9147 17
rect 9181 -17 9219 17
rect 9253 -17 9291 17
rect 9325 -17 9363 17
rect 9397 -17 9435 17
rect 9469 -17 9507 17
rect 9541 -17 9579 17
rect 9613 -17 9651 17
rect 9685 -17 9723 17
rect 9757 -17 9795 17
rect 9829 -17 9867 17
rect 9901 -17 9939 17
rect 9973 -17 10011 17
rect 10045 -17 10083 17
rect 10117 -17 10155 17
rect 10189 -17 10227 17
rect 10261 -17 10299 17
rect 10333 -17 10371 17
rect 10405 -17 10443 17
rect 10477 -17 10515 17
rect 10549 -17 10587 17
rect 10621 -17 10659 17
rect 10693 -17 10731 17
rect 10765 -17 10803 17
rect 10837 -17 10875 17
rect 10909 -17 10947 17
rect 10981 -17 11019 17
rect 11053 -17 11091 17
rect 11125 -17 11163 17
rect 11197 -17 11235 17
rect 11269 -17 11307 17
rect 11341 -17 11379 17
rect 11413 -17 11451 17
rect 11485 -17 11523 17
rect 11557 -17 11595 17
rect 11629 -17 11667 17
rect 11701 -17 11739 17
rect 11773 -17 11811 17
rect 11845 -17 11883 17
rect 11917 -17 11955 17
rect 11989 -17 12027 17
rect 12061 -17 12099 17
rect 12133 -17 12171 17
rect 12205 -17 12243 17
rect 12277 -17 12315 17
rect 12349 -17 12387 17
rect 12421 -17 12459 17
rect 12493 -17 12531 17
rect 12565 -17 12603 17
rect 12637 -17 12675 17
rect 12709 -17 12747 17
rect 12781 -17 12819 17
rect 12853 -17 12891 17
rect 12925 -17 12963 17
rect 12997 -17 13035 17
rect 13069 -17 13107 17
rect 13141 -17 13179 17
rect 13213 -17 13251 17
rect 13285 -17 13327 17
rect -53 -53 13327 -17
use sky130_fd_pr__pfet_01v8_C9QZQZ  sky130_fd_pr__pfet_01v8_C9QZQZ_0
timestamp 1750100919
transform 0 1 4382 -1 0 193
box -246 -4435 246 4435
use sky130_fd_pr__nfet_01v8_MKNP2D  XM2
timestamp 1750100919
transform 0 1 11072 -1 0 193
box -236 -2245 236 2245
<< labels >>
flabel metal1 s -36 408 -22 422 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s -32 -37 -18 -23 0 FreeSans 500 0 0 0 VSS
port 2 nsew
flabel metal1 s -42 184 -28 198 0 FreeSans 500 0 0 0 SWP
port 3 nsew
flabel metal1 s -42 299 -28 313 0 FreeSans 500 0 0 0 IN
port 4 nsew
flabel metal1 s 13302 179 13316 193 0 FreeSans 500 0 0 0 SWN
port 5 nsew
flabel metal1 s 13306 74 13320 88 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
