magic
tech sky130A
magscale 1 2
timestamp 1749060920
<< nwell >>
rect -194 -398 194 364
<< pmos >>
rect -100 -336 100 264
<< pdiff >>
rect -158 252 -100 264
rect -158 -324 -146 252
rect -112 -324 -100 252
rect -158 -336 -100 -324
rect 100 252 158 264
rect 100 -324 112 252
rect 146 -324 158 252
rect 100 -336 158 -324
<< pdiffc >>
rect -146 -324 -112 252
rect 112 -324 146 252
<< poly >>
rect -58 345 58 361
rect -58 328 -42 345
rect -100 311 -42 328
rect 42 328 58 345
rect 42 311 100 328
rect -100 264 100 311
rect -100 -362 100 -336
<< polycont >>
rect -42 311 42 345
<< locali >>
rect -58 311 -42 345
rect 42 311 58 345
rect -146 252 -112 268
rect -146 -340 -112 -324
rect 112 252 146 268
rect 112 -340 146 -324
<< viali >>
rect -42 311 42 345
rect -146 -324 -112 252
rect 112 -324 146 252
<< metal1 >>
rect -54 345 54 351
rect -54 311 -42 345
rect 42 311 54 345
rect -54 305 54 311
rect -152 252 -106 264
rect -152 -324 -146 252
rect -112 -324 -106 252
rect -152 -336 -106 -324
rect 106 252 152 264
rect 106 -324 112 252
rect 146 -324 152 252
rect 106 -336 152 -324
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.0 l 1.0 m 1 nf 1 diffcov 100 polycov 50 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
