/home/mthudaa/vlsi/8bit_SAR-ADC_ITS/magic/th_dif_sw.pex.spice