magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect 142 1527 176 1561
rect 210 1527 248 1561
rect 282 1527 320 1561
rect 354 1527 392 1561
rect 426 1527 464 1561
rect 498 1527 536 1561
rect 570 1527 608 1561
rect 642 1527 680 1561
rect 714 1527 752 1561
rect 786 1527 824 1561
rect 858 1527 896 1561
rect 930 1527 968 1561
rect 1002 1527 1040 1561
rect 1074 1527 1112 1561
rect 1146 1527 1184 1561
rect 1218 1527 1256 1561
rect 1290 1527 1328 1561
rect 1362 1527 1400 1561
rect 1434 1527 1472 1561
rect 1506 1527 1544 1561
rect 1578 1527 1616 1561
rect 1650 1527 1688 1561
rect 1722 1527 1760 1561
rect 1794 1527 1832 1561
rect 1866 1527 1904 1561
rect 1938 1527 1976 1561
rect 2010 1527 2048 1561
rect 2082 1527 2120 1561
rect 2154 1527 2192 1561
rect 2226 1527 2264 1561
rect 2298 1527 2336 1561
rect 2370 1527 2408 1561
rect 2442 1527 2480 1561
rect 2514 1527 2552 1561
rect 2586 1527 2624 1561
rect 2658 1527 2696 1561
rect 2730 1527 2768 1561
rect 2802 1527 2840 1561
rect 2874 1527 2912 1561
rect 2946 1527 2984 1561
rect 3018 1527 3056 1561
rect 3090 1527 3128 1561
rect 3162 1527 3200 1561
rect 3234 1527 3272 1561
rect 3306 1527 3344 1561
rect 3378 1527 3416 1561
rect 3450 1527 3488 1561
rect 3522 1527 3560 1561
rect 3594 1527 3632 1561
rect 3666 1527 3704 1561
rect 3738 1527 3776 1561
rect 3810 1527 3848 1561
rect 3882 1527 3920 1561
rect 3954 1527 3992 1561
rect 4026 1527 4064 1561
rect 4098 1527 4136 1561
rect 4170 1527 4208 1561
rect 4242 1527 4280 1561
rect 4314 1527 4352 1561
rect 4386 1527 4424 1561
rect 4458 1527 4496 1561
rect 4530 1527 4568 1561
rect 4602 1527 4640 1561
rect 4674 1527 4712 1561
rect 4746 1527 4784 1561
rect 4818 1527 4856 1561
rect 4890 1527 4928 1561
rect 4962 1527 5000 1561
rect 5034 1527 5072 1561
rect 5106 1527 5144 1561
rect 5178 1527 5216 1561
rect 5250 1527 5288 1561
rect 5322 1527 5360 1561
rect 5394 1527 5432 1561
rect 5466 1527 5504 1561
rect 5538 1527 5576 1561
rect 5610 1527 5648 1561
rect 5682 1527 5720 1561
rect 5754 1527 5792 1561
rect 5826 1527 5864 1561
rect 5898 1527 5936 1561
rect 5970 1527 6008 1561
rect 6042 1527 6080 1561
rect 6114 1527 6152 1561
rect 6186 1527 6224 1561
rect 6258 1527 6296 1561
rect 6330 1527 6368 1561
rect 6402 1527 6440 1561
rect 6474 1527 6512 1561
rect 6546 1527 6584 1561
rect 6618 1527 6656 1561
rect 6690 1527 6728 1561
rect 6762 1527 6800 1561
rect 6834 1527 6872 1561
rect 6906 1527 6944 1561
rect 6978 1527 7016 1561
rect 7050 1527 7088 1561
rect 7122 1527 7160 1561
rect 7194 1527 7228 1561
rect 142 -123 160 -89
rect 194 -123 232 -89
rect 266 -123 304 -89
rect 338 -123 376 -89
rect 410 -123 448 -89
rect 482 -123 520 -89
rect 554 -123 592 -89
rect 626 -123 664 -89
rect 698 -123 736 -89
rect 770 -123 808 -89
rect 842 -123 880 -89
rect 914 -123 952 -89
rect 986 -123 1024 -89
rect 1058 -123 1096 -89
rect 1130 -123 1168 -89
rect 1202 -123 1240 -89
rect 1274 -123 1312 -89
rect 1346 -123 1384 -89
rect 1418 -123 1456 -89
rect 1490 -123 1528 -89
rect 1562 -123 1600 -89
rect 1634 -123 1672 -89
rect 1706 -123 1744 -89
rect 1778 -123 1816 -89
rect 1850 -123 1888 -89
rect 1922 -123 1960 -89
rect 1994 -123 2032 -89
rect 2066 -123 2104 -89
rect 2138 -123 2176 -89
rect 2210 -123 2248 -89
rect 2282 -123 2320 -89
rect 2354 -123 2392 -89
rect 2426 -123 2464 -89
rect 2498 -123 2536 -89
rect 2570 -123 2608 -89
rect 2642 -123 2680 -89
rect 2714 -123 2752 -89
rect 2786 -123 2824 -89
rect 2858 -123 2896 -89
rect 2930 -123 2968 -89
rect 3002 -123 3040 -89
rect 3074 -123 3112 -89
rect 3146 -123 3184 -89
rect 3218 -123 3256 -89
rect 3290 -123 3328 -89
rect 3362 -123 3400 -89
rect 3434 -123 3472 -89
rect 3506 -123 3544 -89
rect 3578 -123 3616 -89
rect 3650 -123 3688 -89
rect 3722 -123 3740 -89
<< viali >>
rect 176 1527 210 1561
rect 248 1527 282 1561
rect 320 1527 354 1561
rect 392 1527 426 1561
rect 464 1527 498 1561
rect 536 1527 570 1561
rect 608 1527 642 1561
rect 680 1527 714 1561
rect 752 1527 786 1561
rect 824 1527 858 1561
rect 896 1527 930 1561
rect 968 1527 1002 1561
rect 1040 1527 1074 1561
rect 1112 1527 1146 1561
rect 1184 1527 1218 1561
rect 1256 1527 1290 1561
rect 1328 1527 1362 1561
rect 1400 1527 1434 1561
rect 1472 1527 1506 1561
rect 1544 1527 1578 1561
rect 1616 1527 1650 1561
rect 1688 1527 1722 1561
rect 1760 1527 1794 1561
rect 1832 1527 1866 1561
rect 1904 1527 1938 1561
rect 1976 1527 2010 1561
rect 2048 1527 2082 1561
rect 2120 1527 2154 1561
rect 2192 1527 2226 1561
rect 2264 1527 2298 1561
rect 2336 1527 2370 1561
rect 2408 1527 2442 1561
rect 2480 1527 2514 1561
rect 2552 1527 2586 1561
rect 2624 1527 2658 1561
rect 2696 1527 2730 1561
rect 2768 1527 2802 1561
rect 2840 1527 2874 1561
rect 2912 1527 2946 1561
rect 2984 1527 3018 1561
rect 3056 1527 3090 1561
rect 3128 1527 3162 1561
rect 3200 1527 3234 1561
rect 3272 1527 3306 1561
rect 3344 1527 3378 1561
rect 3416 1527 3450 1561
rect 3488 1527 3522 1561
rect 3560 1527 3594 1561
rect 3632 1527 3666 1561
rect 3704 1527 3738 1561
rect 3776 1527 3810 1561
rect 3848 1527 3882 1561
rect 3920 1527 3954 1561
rect 3992 1527 4026 1561
rect 4064 1527 4098 1561
rect 4136 1527 4170 1561
rect 4208 1527 4242 1561
rect 4280 1527 4314 1561
rect 4352 1527 4386 1561
rect 4424 1527 4458 1561
rect 4496 1527 4530 1561
rect 4568 1527 4602 1561
rect 4640 1527 4674 1561
rect 4712 1527 4746 1561
rect 4784 1527 4818 1561
rect 4856 1527 4890 1561
rect 4928 1527 4962 1561
rect 5000 1527 5034 1561
rect 5072 1527 5106 1561
rect 5144 1527 5178 1561
rect 5216 1527 5250 1561
rect 5288 1527 5322 1561
rect 5360 1527 5394 1561
rect 5432 1527 5466 1561
rect 5504 1527 5538 1561
rect 5576 1527 5610 1561
rect 5648 1527 5682 1561
rect 5720 1527 5754 1561
rect 5792 1527 5826 1561
rect 5864 1527 5898 1561
rect 5936 1527 5970 1561
rect 6008 1527 6042 1561
rect 6080 1527 6114 1561
rect 6152 1527 6186 1561
rect 6224 1527 6258 1561
rect 6296 1527 6330 1561
rect 6368 1527 6402 1561
rect 6440 1527 6474 1561
rect 6512 1527 6546 1561
rect 6584 1527 6618 1561
rect 6656 1527 6690 1561
rect 6728 1527 6762 1561
rect 6800 1527 6834 1561
rect 6872 1527 6906 1561
rect 6944 1527 6978 1561
rect 7016 1527 7050 1561
rect 7088 1527 7122 1561
rect 7160 1527 7194 1561
rect 160 -123 194 -89
rect 232 -123 266 -89
rect 304 -123 338 -89
rect 376 -123 410 -89
rect 448 -123 482 -89
rect 520 -123 554 -89
rect 592 -123 626 -89
rect 664 -123 698 -89
rect 736 -123 770 -89
rect 808 -123 842 -89
rect 880 -123 914 -89
rect 952 -123 986 -89
rect 1024 -123 1058 -89
rect 1096 -123 1130 -89
rect 1168 -123 1202 -89
rect 1240 -123 1274 -89
rect 1312 -123 1346 -89
rect 1384 -123 1418 -89
rect 1456 -123 1490 -89
rect 1528 -123 1562 -89
rect 1600 -123 1634 -89
rect 1672 -123 1706 -89
rect 1744 -123 1778 -89
rect 1816 -123 1850 -89
rect 1888 -123 1922 -89
rect 1960 -123 1994 -89
rect 2032 -123 2066 -89
rect 2104 -123 2138 -89
rect 2176 -123 2210 -89
rect 2248 -123 2282 -89
rect 2320 -123 2354 -89
rect 2392 -123 2426 -89
rect 2464 -123 2498 -89
rect 2536 -123 2570 -89
rect 2608 -123 2642 -89
rect 2680 -123 2714 -89
rect 2752 -123 2786 -89
rect 2824 -123 2858 -89
rect 2896 -123 2930 -89
rect 2968 -123 3002 -89
rect 3040 -123 3074 -89
rect 3112 -123 3146 -89
rect 3184 -123 3218 -89
rect 3256 -123 3290 -89
rect 3328 -123 3362 -89
rect 3400 -123 3434 -89
rect 3472 -123 3506 -89
rect 3544 -123 3578 -89
rect 3616 -123 3650 -89
rect 3688 -123 3722 -89
<< metal1 >>
rect 106 1561 7264 1597
rect 106 1527 176 1561
rect 210 1527 248 1561
rect 282 1527 320 1561
rect 354 1527 392 1561
rect 426 1527 464 1561
rect 498 1527 536 1561
rect 570 1527 608 1561
rect 642 1527 680 1561
rect 714 1527 752 1561
rect 786 1527 824 1561
rect 858 1527 896 1561
rect 930 1527 968 1561
rect 1002 1527 1040 1561
rect 1074 1527 1112 1561
rect 1146 1527 1184 1561
rect 1218 1527 1256 1561
rect 1290 1527 1328 1561
rect 1362 1527 1400 1561
rect 1434 1527 1472 1561
rect 1506 1527 1544 1561
rect 1578 1527 1616 1561
rect 1650 1527 1688 1561
rect 1722 1527 1760 1561
rect 1794 1527 1832 1561
rect 1866 1527 1904 1561
rect 1938 1527 1976 1561
rect 2010 1527 2048 1561
rect 2082 1527 2120 1561
rect 2154 1527 2192 1561
rect 2226 1527 2264 1561
rect 2298 1527 2336 1561
rect 2370 1527 2408 1561
rect 2442 1527 2480 1561
rect 2514 1527 2552 1561
rect 2586 1527 2624 1561
rect 2658 1527 2696 1561
rect 2730 1527 2768 1561
rect 2802 1527 2840 1561
rect 2874 1527 2912 1561
rect 2946 1527 2984 1561
rect 3018 1527 3056 1561
rect 3090 1527 3128 1561
rect 3162 1527 3200 1561
rect 3234 1527 3272 1561
rect 3306 1527 3344 1561
rect 3378 1527 3416 1561
rect 3450 1527 3488 1561
rect 3522 1527 3560 1561
rect 3594 1527 3632 1561
rect 3666 1527 3704 1561
rect 3738 1527 3776 1561
rect 3810 1527 3848 1561
rect 3882 1527 3920 1561
rect 3954 1527 3992 1561
rect 4026 1527 4064 1561
rect 4098 1527 4136 1561
rect 4170 1527 4208 1561
rect 4242 1527 4280 1561
rect 4314 1527 4352 1561
rect 4386 1527 4424 1561
rect 4458 1527 4496 1561
rect 4530 1527 4568 1561
rect 4602 1527 4640 1561
rect 4674 1527 4712 1561
rect 4746 1527 4784 1561
rect 4818 1527 4856 1561
rect 4890 1527 4928 1561
rect 4962 1527 5000 1561
rect 5034 1527 5072 1561
rect 5106 1527 5144 1561
rect 5178 1527 5216 1561
rect 5250 1527 5288 1561
rect 5322 1527 5360 1561
rect 5394 1527 5432 1561
rect 5466 1527 5504 1561
rect 5538 1527 5576 1561
rect 5610 1527 5648 1561
rect 5682 1527 5720 1561
rect 5754 1527 5792 1561
rect 5826 1527 5864 1561
rect 5898 1527 5936 1561
rect 5970 1527 6008 1561
rect 6042 1527 6080 1561
rect 6114 1527 6152 1561
rect 6186 1527 6224 1561
rect 6258 1527 6296 1561
rect 6330 1527 6368 1561
rect 6402 1527 6440 1561
rect 6474 1527 6512 1561
rect 6546 1527 6584 1561
rect 6618 1527 6656 1561
rect 6690 1527 6728 1561
rect 6762 1527 6800 1561
rect 6834 1527 6872 1561
rect 6906 1527 6944 1561
rect 6978 1527 7016 1561
rect 7050 1527 7088 1561
rect 7122 1527 7160 1561
rect 7194 1527 7264 1561
rect 106 1521 7264 1527
rect 325 1447 7045 1521
rect 106 1377 284 1401
rect 106 1325 176 1377
rect 228 1325 284 1377
rect 106 1301 284 1325
rect 325 1061 7045 1255
rect 106 915 284 1015
rect 106 569 7264 869
rect 106 423 284 523
rect 316 183 3566 377
rect 166 113 284 137
rect 166 61 176 113
rect 228 61 284 113
rect 166 37 284 61
rect 316 -83 3566 -9
rect 106 -89 7264 -83
rect 106 -123 160 -89
rect 194 -123 232 -89
rect 266 -123 304 -89
rect 338 -123 376 -89
rect 410 -123 448 -89
rect 482 -123 520 -89
rect 554 -123 592 -89
rect 626 -123 664 -89
rect 698 -123 736 -89
rect 770 -123 808 -89
rect 842 -123 880 -89
rect 914 -123 952 -89
rect 986 -123 1024 -89
rect 1058 -123 1096 -89
rect 1130 -123 1168 -89
rect 1202 -123 1240 -89
rect 1274 -123 1312 -89
rect 1346 -123 1384 -89
rect 1418 -123 1456 -89
rect 1490 -123 1528 -89
rect 1562 -123 1600 -89
rect 1634 -123 1672 -89
rect 1706 -123 1744 -89
rect 1778 -123 1816 -89
rect 1850 -123 1888 -89
rect 1922 -123 1960 -89
rect 1994 -123 2032 -89
rect 2066 -123 2104 -89
rect 2138 -123 2176 -89
rect 2210 -123 2248 -89
rect 2282 -123 2320 -89
rect 2354 -123 2392 -89
rect 2426 -123 2464 -89
rect 2498 -123 2536 -89
rect 2570 -123 2608 -89
rect 2642 -123 2680 -89
rect 2714 -123 2752 -89
rect 2786 -123 2824 -89
rect 2858 -123 2896 -89
rect 2930 -123 2968 -89
rect 3002 -123 3040 -89
rect 3074 -123 3112 -89
rect 3146 -123 3184 -89
rect 3218 -123 3256 -89
rect 3290 -123 3328 -89
rect 3362 -123 3400 -89
rect 3434 -123 3472 -89
rect 3506 -123 3544 -89
rect 3578 -123 3616 -89
rect 3650 -123 3688 -89
rect 3722 -123 7264 -89
rect 106 -159 7264 -123
<< via1 >>
rect 176 1325 228 1377
rect 176 61 228 113
<< metal2 >>
rect 176 1377 228 1411
rect 176 113 228 1325
rect 176 27 228 61
use sky130_fd_pr__nfet_01v8_K9ZN2D  sky130_fd_pr__nfet_01v8_K9ZN2D_0
timestamp 1750100919
transform 0 1 1941 -1 0 87
box -236 -1825 236 1825
use sky130_fd_pr__pfet_01v8_D9Q5W2  sky130_fd_pr__pfet_01v8_D9Q5W2_0
timestamp 1750100919
transform 0 1 3685 -1 0 965
box -246 -3579 246 3579
use sky130_fd_pr__pfet_01v8_D9Q5W2  XM1
timestamp 1750100919
transform 0 1 3685 -1 0 1351
box -246 -3579 246 3579
use sky130_fd_pr__nfet_01v8_K9ZN2D  XM3
timestamp 1750100919
transform 0 1 1941 -1 0 473
box -236 -1825 236 1825
<< labels >>
flabel metal1 s 122 1555 130 1564 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 119 1343 127 1352 0 FreeSans 500 0 0 0 IN
port 2 nsew
flabel metal1 s 122 959 130 968 0 FreeSans 500 0 0 0 CKB
port 3 nsew
flabel metal1 s 120 466 128 475 0 FreeSans 500 0 0 0 CK
port 4 nsew
flabel metal1 s 123 -126 131 -117 0 FreeSans 500 0 0 0 VSS
port 5 nsew
flabel metal1 s 7220 701 7228 710 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
