magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< dnwell >>
rect -2373 100892 47207 116761
rect -10676 64109 -3707 76121
rect -7184 56281 -3707 64109
rect 50479 58365 56327 62017
rect -10676 44269 -3707 56281
rect 59127 45909 70849 74783
rect -2373 3629 47207 19498
<< nwell >>
rect -2453 116555 47287 116841
rect -2453 101098 -2167 116555
rect 47001 101098 47287 116555
rect -2453 100812 47287 101098
rect -10756 75915 -3627 76201
rect -10756 64315 -10470 75915
rect -10756 64029 -6978 64315
rect -7264 56361 -6978 64029
rect -10756 56075 -6978 56361
rect -10756 44475 -10470 56075
rect -3913 44475 -3627 75915
rect 59047 74577 70929 74863
rect 50399 61811 56407 62097
rect 50399 58571 50685 61811
rect 56121 58571 56407 61811
rect 50399 58285 56407 58571
rect 59047 46115 59333 74577
rect 70643 46115 70929 74577
rect 59047 45829 70929 46115
rect -10756 44189 -3627 44475
rect -2453 19292 47287 19578
rect -2453 3835 -2167 19292
rect 47001 3835 47287 19292
rect -2453 3549 47287 3835
<< nsubdiff >>
rect -2416 116784 47250 116804
rect -2416 116750 -2318 116784
rect -2284 116750 -2250 116784
rect -2216 116750 -2182 116784
rect -2148 116750 -2114 116784
rect -2080 116750 -2046 116784
rect -2012 116750 -1978 116784
rect -1944 116750 -1910 116784
rect -1876 116750 -1842 116784
rect -1808 116750 -1774 116784
rect -1740 116750 -1706 116784
rect -1672 116750 -1638 116784
rect -1604 116750 -1570 116784
rect -1536 116750 -1502 116784
rect -1468 116750 -1434 116784
rect -1400 116750 -1366 116784
rect -1332 116750 -1298 116784
rect -1264 116750 -1230 116784
rect -1196 116750 -1162 116784
rect -1128 116750 -1094 116784
rect -1060 116750 -1026 116784
rect -992 116750 -958 116784
rect -924 116750 -890 116784
rect -856 116750 -822 116784
rect -788 116750 -754 116784
rect -720 116750 -686 116784
rect -652 116750 -618 116784
rect -584 116750 -550 116784
rect -516 116750 -482 116784
rect -448 116750 -414 116784
rect -380 116750 -346 116784
rect -312 116750 -278 116784
rect -244 116750 -210 116784
rect -176 116750 -142 116784
rect -108 116750 -74 116784
rect -40 116750 -6 116784
rect 28 116750 62 116784
rect 96 116750 130 116784
rect 164 116750 198 116784
rect 232 116750 266 116784
rect 300 116750 334 116784
rect 368 116750 402 116784
rect 436 116750 470 116784
rect 504 116750 538 116784
rect 572 116750 606 116784
rect 640 116750 674 116784
rect 708 116750 742 116784
rect 776 116750 810 116784
rect 844 116750 878 116784
rect 912 116750 946 116784
rect 980 116750 1014 116784
rect 1048 116750 1082 116784
rect 1116 116750 1150 116784
rect 1184 116750 1218 116784
rect 1252 116750 1286 116784
rect 1320 116750 1354 116784
rect 1388 116750 1422 116784
rect 1456 116750 1490 116784
rect 1524 116750 1558 116784
rect 1592 116750 1626 116784
rect 1660 116750 1694 116784
rect 1728 116750 1762 116784
rect 1796 116750 1830 116784
rect 1864 116750 1898 116784
rect 1932 116750 1966 116784
rect 2000 116750 2034 116784
rect 2068 116750 2102 116784
rect 2136 116750 2170 116784
rect 2204 116750 2238 116784
rect 2272 116750 2306 116784
rect 2340 116750 2374 116784
rect 2408 116750 2442 116784
rect 2476 116750 2510 116784
rect 2544 116750 2578 116784
rect 2612 116750 2646 116784
rect 2680 116750 2714 116784
rect 2748 116750 2782 116784
rect 2816 116750 2850 116784
rect 2884 116750 2918 116784
rect 2952 116750 2986 116784
rect 3020 116750 3054 116784
rect 3088 116750 3122 116784
rect 3156 116750 3190 116784
rect 3224 116750 3258 116784
rect 3292 116750 3326 116784
rect 3360 116750 3394 116784
rect 3428 116750 3462 116784
rect 3496 116750 3530 116784
rect 3564 116750 3598 116784
rect 3632 116750 3666 116784
rect 3700 116750 3734 116784
rect 3768 116750 3802 116784
rect 3836 116750 3870 116784
rect 3904 116750 3938 116784
rect 3972 116750 4006 116784
rect 4040 116750 4074 116784
rect 4108 116750 4142 116784
rect 4176 116750 4210 116784
rect 4244 116750 4278 116784
rect 4312 116750 4346 116784
rect 4380 116750 4414 116784
rect 4448 116750 4482 116784
rect 4516 116750 4550 116784
rect 4584 116750 4618 116784
rect 4652 116750 4686 116784
rect 4720 116750 4754 116784
rect 4788 116750 4822 116784
rect 4856 116750 4890 116784
rect 4924 116750 4958 116784
rect 4992 116750 5026 116784
rect 5060 116750 5094 116784
rect 5128 116750 5162 116784
rect 5196 116750 5230 116784
rect 5264 116750 5298 116784
rect 5332 116750 5366 116784
rect 5400 116750 5434 116784
rect 5468 116750 5502 116784
rect 5536 116750 5570 116784
rect 5604 116750 5638 116784
rect 5672 116750 5706 116784
rect 5740 116750 5774 116784
rect 5808 116750 5842 116784
rect 5876 116750 5910 116784
rect 5944 116750 5978 116784
rect 6012 116750 6046 116784
rect 6080 116750 6114 116784
rect 6148 116750 6182 116784
rect 6216 116750 6250 116784
rect 6284 116750 6318 116784
rect 6352 116750 6386 116784
rect 6420 116750 6454 116784
rect 6488 116750 6522 116784
rect 6556 116750 6590 116784
rect 6624 116750 6658 116784
rect 6692 116750 6726 116784
rect 6760 116750 6794 116784
rect 6828 116750 6862 116784
rect 6896 116750 6930 116784
rect 6964 116750 6998 116784
rect 7032 116750 7066 116784
rect 7100 116750 7134 116784
rect 7168 116750 7202 116784
rect 7236 116750 7270 116784
rect 7304 116750 7338 116784
rect 7372 116750 7406 116784
rect 7440 116750 7474 116784
rect 7508 116750 7542 116784
rect 7576 116750 7610 116784
rect 7644 116750 7678 116784
rect 7712 116750 7746 116784
rect 7780 116750 7814 116784
rect 7848 116750 7882 116784
rect 7916 116750 7950 116784
rect 7984 116750 8018 116784
rect 8052 116750 8086 116784
rect 8120 116750 8154 116784
rect 8188 116750 8222 116784
rect 8256 116750 8290 116784
rect 8324 116750 8358 116784
rect 8392 116750 8426 116784
rect 8460 116750 8494 116784
rect 8528 116750 8562 116784
rect 8596 116750 8630 116784
rect 8664 116750 8698 116784
rect 8732 116750 8766 116784
rect 8800 116750 8834 116784
rect 8868 116750 8902 116784
rect 8936 116750 8970 116784
rect 9004 116750 9038 116784
rect 9072 116750 9106 116784
rect 9140 116750 9174 116784
rect 9208 116750 9242 116784
rect 9276 116750 9310 116784
rect 9344 116750 9378 116784
rect 9412 116750 9446 116784
rect 9480 116750 9514 116784
rect 9548 116750 9582 116784
rect 9616 116750 9650 116784
rect 9684 116750 9718 116784
rect 9752 116750 9786 116784
rect 9820 116750 9854 116784
rect 9888 116750 9922 116784
rect 9956 116750 9990 116784
rect 10024 116750 10058 116784
rect 10092 116750 10126 116784
rect 10160 116750 10194 116784
rect 10228 116750 10262 116784
rect 10296 116750 10330 116784
rect 10364 116750 10398 116784
rect 10432 116750 10466 116784
rect 10500 116750 10534 116784
rect 10568 116750 10602 116784
rect 10636 116750 10670 116784
rect 10704 116750 10738 116784
rect 10772 116750 10806 116784
rect 10840 116750 10874 116784
rect 10908 116750 10942 116784
rect 10976 116750 11010 116784
rect 11044 116750 11078 116784
rect 11112 116750 11146 116784
rect 11180 116750 11214 116784
rect 11248 116750 11282 116784
rect 11316 116750 11350 116784
rect 11384 116750 11418 116784
rect 11452 116750 11486 116784
rect 11520 116750 11554 116784
rect 11588 116750 11622 116784
rect 11656 116750 11690 116784
rect 11724 116750 11758 116784
rect 11792 116750 11826 116784
rect 11860 116750 11894 116784
rect 11928 116750 11962 116784
rect 11996 116750 12030 116784
rect 12064 116750 12098 116784
rect 12132 116750 12166 116784
rect 12200 116750 12234 116784
rect 12268 116750 12302 116784
rect 12336 116750 12370 116784
rect 12404 116750 12438 116784
rect 12472 116750 12506 116784
rect 12540 116750 12574 116784
rect 12608 116750 12642 116784
rect 12676 116750 12710 116784
rect 12744 116750 12778 116784
rect 12812 116750 12846 116784
rect 12880 116750 12914 116784
rect 12948 116750 12982 116784
rect 13016 116750 13050 116784
rect 13084 116750 13118 116784
rect 13152 116750 13186 116784
rect 13220 116750 13254 116784
rect 13288 116750 13322 116784
rect 13356 116750 13390 116784
rect 13424 116750 13458 116784
rect 13492 116750 13526 116784
rect 13560 116750 13594 116784
rect 13628 116750 13662 116784
rect 13696 116750 13730 116784
rect 13764 116750 13798 116784
rect 13832 116750 13866 116784
rect 13900 116750 13934 116784
rect 13968 116750 14002 116784
rect 14036 116750 14070 116784
rect 14104 116750 14138 116784
rect 14172 116750 14206 116784
rect 14240 116750 14274 116784
rect 14308 116750 14342 116784
rect 14376 116750 14410 116784
rect 14444 116750 14478 116784
rect 14512 116750 14546 116784
rect 14580 116750 14614 116784
rect 14648 116750 14682 116784
rect 14716 116750 14750 116784
rect 14784 116750 14818 116784
rect 14852 116750 14886 116784
rect 14920 116750 14954 116784
rect 14988 116750 15022 116784
rect 15056 116750 15090 116784
rect 15124 116750 15158 116784
rect 15192 116750 15226 116784
rect 15260 116750 15294 116784
rect 15328 116750 15362 116784
rect 15396 116750 15430 116784
rect 15464 116750 15498 116784
rect 15532 116750 15566 116784
rect 15600 116750 15634 116784
rect 15668 116750 15702 116784
rect 15736 116750 15770 116784
rect 15804 116750 15838 116784
rect 15872 116750 15906 116784
rect 15940 116750 15974 116784
rect 16008 116750 16042 116784
rect 16076 116750 16110 116784
rect 16144 116750 16178 116784
rect 16212 116750 16246 116784
rect 16280 116750 16314 116784
rect 16348 116750 16382 116784
rect 16416 116750 16450 116784
rect 16484 116750 16518 116784
rect 16552 116750 16586 116784
rect 16620 116750 16654 116784
rect 16688 116750 16722 116784
rect 16756 116750 16790 116784
rect 16824 116750 16858 116784
rect 16892 116750 16926 116784
rect 16960 116750 16994 116784
rect 17028 116750 17062 116784
rect 17096 116750 17130 116784
rect 17164 116750 17198 116784
rect 17232 116750 17266 116784
rect 17300 116750 17334 116784
rect 17368 116750 17402 116784
rect 17436 116750 17470 116784
rect 17504 116750 17538 116784
rect 17572 116750 17606 116784
rect 17640 116750 17674 116784
rect 17708 116750 17742 116784
rect 17776 116750 17810 116784
rect 17844 116750 17878 116784
rect 17912 116750 17946 116784
rect 17980 116750 18014 116784
rect 18048 116750 18082 116784
rect 18116 116750 18150 116784
rect 18184 116750 18218 116784
rect 18252 116750 18286 116784
rect 18320 116750 18354 116784
rect 18388 116750 18422 116784
rect 18456 116750 18490 116784
rect 18524 116750 18558 116784
rect 18592 116750 18626 116784
rect 18660 116750 18694 116784
rect 18728 116750 18762 116784
rect 18796 116750 18830 116784
rect 18864 116750 18898 116784
rect 18932 116750 18966 116784
rect 19000 116750 19034 116784
rect 19068 116750 19102 116784
rect 19136 116750 19170 116784
rect 19204 116750 19238 116784
rect 19272 116750 19306 116784
rect 19340 116750 19374 116784
rect 19408 116750 19442 116784
rect 19476 116750 19510 116784
rect 19544 116750 19578 116784
rect 19612 116750 19646 116784
rect 19680 116750 19714 116784
rect 19748 116750 19782 116784
rect 19816 116750 19850 116784
rect 19884 116750 19918 116784
rect 19952 116750 19986 116784
rect 20020 116750 20054 116784
rect 20088 116750 20122 116784
rect 20156 116750 20190 116784
rect 20224 116750 20258 116784
rect 20292 116750 20326 116784
rect 20360 116750 20394 116784
rect 20428 116750 20462 116784
rect 20496 116750 20530 116784
rect 20564 116750 20598 116784
rect 20632 116750 20666 116784
rect 20700 116750 20734 116784
rect 20768 116750 20802 116784
rect 20836 116750 20870 116784
rect 20904 116750 20938 116784
rect 20972 116750 21006 116784
rect 21040 116750 21074 116784
rect 21108 116750 21142 116784
rect 21176 116750 21210 116784
rect 21244 116750 21278 116784
rect 21312 116750 21346 116784
rect 21380 116750 21414 116784
rect 21448 116750 21482 116784
rect 21516 116750 21550 116784
rect 21584 116750 21618 116784
rect 21652 116750 21686 116784
rect 21720 116750 21754 116784
rect 21788 116750 21822 116784
rect 21856 116750 21890 116784
rect 21924 116750 21958 116784
rect 21992 116750 22026 116784
rect 22060 116750 22094 116784
rect 22128 116750 22162 116784
rect 22196 116750 22230 116784
rect 22264 116750 22298 116784
rect 22332 116750 22366 116784
rect 22400 116750 22434 116784
rect 22468 116750 22502 116784
rect 22536 116750 22570 116784
rect 22604 116750 22638 116784
rect 22672 116750 22706 116784
rect 22740 116750 22774 116784
rect 22808 116750 22842 116784
rect 22876 116750 22910 116784
rect 22944 116750 22978 116784
rect 23012 116750 23046 116784
rect 23080 116750 23114 116784
rect 23148 116750 23182 116784
rect 23216 116750 23250 116784
rect 23284 116750 23318 116784
rect 23352 116750 23386 116784
rect 23420 116750 23454 116784
rect 23488 116750 23522 116784
rect 23556 116750 23590 116784
rect 23624 116750 23658 116784
rect 23692 116750 23726 116784
rect 23760 116750 23794 116784
rect 23828 116750 23862 116784
rect 23896 116750 23930 116784
rect 23964 116750 23998 116784
rect 24032 116750 24066 116784
rect 24100 116750 24134 116784
rect 24168 116750 24202 116784
rect 24236 116750 24270 116784
rect 24304 116750 24338 116784
rect 24372 116750 24406 116784
rect 24440 116750 24474 116784
rect 24508 116750 24542 116784
rect 24576 116750 24610 116784
rect 24644 116750 24678 116784
rect 24712 116750 24746 116784
rect 24780 116750 24814 116784
rect 24848 116750 24882 116784
rect 24916 116750 24950 116784
rect 24984 116750 25018 116784
rect 25052 116750 25086 116784
rect 25120 116750 25154 116784
rect 25188 116750 25222 116784
rect 25256 116750 25290 116784
rect 25324 116750 25358 116784
rect 25392 116750 25426 116784
rect 25460 116750 25494 116784
rect 25528 116750 25562 116784
rect 25596 116750 25630 116784
rect 25664 116750 25698 116784
rect 25732 116750 25766 116784
rect 25800 116750 25834 116784
rect 25868 116750 25902 116784
rect 25936 116750 25970 116784
rect 26004 116750 26038 116784
rect 26072 116750 26106 116784
rect 26140 116750 26174 116784
rect 26208 116750 26242 116784
rect 26276 116750 26310 116784
rect 26344 116750 26378 116784
rect 26412 116750 26446 116784
rect 26480 116750 26514 116784
rect 26548 116750 26582 116784
rect 26616 116750 26650 116784
rect 26684 116750 26718 116784
rect 26752 116750 26786 116784
rect 26820 116750 26854 116784
rect 26888 116750 26922 116784
rect 26956 116750 26990 116784
rect 27024 116750 27058 116784
rect 27092 116750 27126 116784
rect 27160 116750 27194 116784
rect 27228 116750 27262 116784
rect 27296 116750 27330 116784
rect 27364 116750 27398 116784
rect 27432 116750 27466 116784
rect 27500 116750 27534 116784
rect 27568 116750 27602 116784
rect 27636 116750 27670 116784
rect 27704 116750 27738 116784
rect 27772 116750 27806 116784
rect 27840 116750 27874 116784
rect 27908 116750 27942 116784
rect 27976 116750 28010 116784
rect 28044 116750 28078 116784
rect 28112 116750 28146 116784
rect 28180 116750 28214 116784
rect 28248 116750 28282 116784
rect 28316 116750 28350 116784
rect 28384 116750 28418 116784
rect 28452 116750 28486 116784
rect 28520 116750 28554 116784
rect 28588 116750 28622 116784
rect 28656 116750 28690 116784
rect 28724 116750 28758 116784
rect 28792 116750 28826 116784
rect 28860 116750 28894 116784
rect 28928 116750 28962 116784
rect 28996 116750 29030 116784
rect 29064 116750 29098 116784
rect 29132 116750 29166 116784
rect 29200 116750 29234 116784
rect 29268 116750 29302 116784
rect 29336 116750 29370 116784
rect 29404 116750 29438 116784
rect 29472 116750 29506 116784
rect 29540 116750 29574 116784
rect 29608 116750 29642 116784
rect 29676 116750 29710 116784
rect 29744 116750 29778 116784
rect 29812 116750 29846 116784
rect 29880 116750 29914 116784
rect 29948 116750 29982 116784
rect 30016 116750 30050 116784
rect 30084 116750 30118 116784
rect 30152 116750 30186 116784
rect 30220 116750 30254 116784
rect 30288 116750 30322 116784
rect 30356 116750 30390 116784
rect 30424 116750 30458 116784
rect 30492 116750 30526 116784
rect 30560 116750 30594 116784
rect 30628 116750 30662 116784
rect 30696 116750 30730 116784
rect 30764 116750 30798 116784
rect 30832 116750 30866 116784
rect 30900 116750 30934 116784
rect 30968 116750 31002 116784
rect 31036 116750 31070 116784
rect 31104 116750 31138 116784
rect 31172 116750 31206 116784
rect 31240 116750 31274 116784
rect 31308 116750 31342 116784
rect 31376 116750 31410 116784
rect 31444 116750 31478 116784
rect 31512 116750 31546 116784
rect 31580 116750 31614 116784
rect 31648 116750 31682 116784
rect 31716 116750 31750 116784
rect 31784 116750 31818 116784
rect 31852 116750 31886 116784
rect 31920 116750 31954 116784
rect 31988 116750 32022 116784
rect 32056 116750 32090 116784
rect 32124 116750 32158 116784
rect 32192 116750 32226 116784
rect 32260 116750 32294 116784
rect 32328 116750 32362 116784
rect 32396 116750 32430 116784
rect 32464 116750 32498 116784
rect 32532 116750 32566 116784
rect 32600 116750 32634 116784
rect 32668 116750 32702 116784
rect 32736 116750 32770 116784
rect 32804 116750 32838 116784
rect 32872 116750 32906 116784
rect 32940 116750 32974 116784
rect 33008 116750 33042 116784
rect 33076 116750 33110 116784
rect 33144 116750 33178 116784
rect 33212 116750 33246 116784
rect 33280 116750 33314 116784
rect 33348 116750 33382 116784
rect 33416 116750 33450 116784
rect 33484 116750 33518 116784
rect 33552 116750 33586 116784
rect 33620 116750 33654 116784
rect 33688 116750 33722 116784
rect 33756 116750 33790 116784
rect 33824 116750 33858 116784
rect 33892 116750 33926 116784
rect 33960 116750 33994 116784
rect 34028 116750 34062 116784
rect 34096 116750 34130 116784
rect 34164 116750 34198 116784
rect 34232 116750 34266 116784
rect 34300 116750 34334 116784
rect 34368 116750 34402 116784
rect 34436 116750 34470 116784
rect 34504 116750 34538 116784
rect 34572 116750 34606 116784
rect 34640 116750 34674 116784
rect 34708 116750 34742 116784
rect 34776 116750 34810 116784
rect 34844 116750 34878 116784
rect 34912 116750 34946 116784
rect 34980 116750 35014 116784
rect 35048 116750 35082 116784
rect 35116 116750 35150 116784
rect 35184 116750 35218 116784
rect 35252 116750 35286 116784
rect 35320 116750 35354 116784
rect 35388 116750 35422 116784
rect 35456 116750 35490 116784
rect 35524 116750 35558 116784
rect 35592 116750 35626 116784
rect 35660 116750 35694 116784
rect 35728 116750 35762 116784
rect 35796 116750 35830 116784
rect 35864 116750 35898 116784
rect 35932 116750 35966 116784
rect 36000 116750 36034 116784
rect 36068 116750 36102 116784
rect 36136 116750 36170 116784
rect 36204 116750 36238 116784
rect 36272 116750 36306 116784
rect 36340 116750 36374 116784
rect 36408 116750 36442 116784
rect 36476 116750 36510 116784
rect 36544 116750 36578 116784
rect 36612 116750 36646 116784
rect 36680 116750 36714 116784
rect 36748 116750 36782 116784
rect 36816 116750 36850 116784
rect 36884 116750 36918 116784
rect 36952 116750 36986 116784
rect 37020 116750 37054 116784
rect 37088 116750 37122 116784
rect 37156 116750 37190 116784
rect 37224 116750 37258 116784
rect 37292 116750 37326 116784
rect 37360 116750 37394 116784
rect 37428 116750 37462 116784
rect 37496 116750 37530 116784
rect 37564 116750 37598 116784
rect 37632 116750 37666 116784
rect 37700 116750 37734 116784
rect 37768 116750 37802 116784
rect 37836 116750 37870 116784
rect 37904 116750 37938 116784
rect 37972 116750 38006 116784
rect 38040 116750 38074 116784
rect 38108 116750 38142 116784
rect 38176 116750 38210 116784
rect 38244 116750 38278 116784
rect 38312 116750 38346 116784
rect 38380 116750 38414 116784
rect 38448 116750 38482 116784
rect 38516 116750 38550 116784
rect 38584 116750 38618 116784
rect 38652 116750 38686 116784
rect 38720 116750 38754 116784
rect 38788 116750 38822 116784
rect 38856 116750 38890 116784
rect 38924 116750 38958 116784
rect 38992 116750 39026 116784
rect 39060 116750 39094 116784
rect 39128 116750 39162 116784
rect 39196 116750 39230 116784
rect 39264 116750 39298 116784
rect 39332 116750 39366 116784
rect 39400 116750 39434 116784
rect 39468 116750 39502 116784
rect 39536 116750 39570 116784
rect 39604 116750 39638 116784
rect 39672 116750 39706 116784
rect 39740 116750 39774 116784
rect 39808 116750 39842 116784
rect 39876 116750 39910 116784
rect 39944 116750 39978 116784
rect 40012 116750 40046 116784
rect 40080 116750 40114 116784
rect 40148 116750 40182 116784
rect 40216 116750 40250 116784
rect 40284 116750 40318 116784
rect 40352 116750 40386 116784
rect 40420 116750 40454 116784
rect 40488 116750 40522 116784
rect 40556 116750 40590 116784
rect 40624 116750 40658 116784
rect 40692 116750 40726 116784
rect 40760 116750 40794 116784
rect 40828 116750 40862 116784
rect 40896 116750 40930 116784
rect 40964 116750 40998 116784
rect 41032 116750 41066 116784
rect 41100 116750 41134 116784
rect 41168 116750 41202 116784
rect 41236 116750 41270 116784
rect 41304 116750 41338 116784
rect 41372 116750 41406 116784
rect 41440 116750 41474 116784
rect 41508 116750 41542 116784
rect 41576 116750 41610 116784
rect 41644 116750 41678 116784
rect 41712 116750 41746 116784
rect 41780 116750 41814 116784
rect 41848 116750 41882 116784
rect 41916 116750 41950 116784
rect 41984 116750 42018 116784
rect 42052 116750 42086 116784
rect 42120 116750 42154 116784
rect 42188 116750 42222 116784
rect 42256 116750 42290 116784
rect 42324 116750 42358 116784
rect 42392 116750 42426 116784
rect 42460 116750 42494 116784
rect 42528 116750 42562 116784
rect 42596 116750 42630 116784
rect 42664 116750 42698 116784
rect 42732 116750 42766 116784
rect 42800 116750 42834 116784
rect 42868 116750 42902 116784
rect 42936 116750 42970 116784
rect 43004 116750 43038 116784
rect 43072 116750 43106 116784
rect 43140 116750 43174 116784
rect 43208 116750 43242 116784
rect 43276 116750 43310 116784
rect 43344 116750 43378 116784
rect 43412 116750 43446 116784
rect 43480 116750 43514 116784
rect 43548 116750 43582 116784
rect 43616 116750 43650 116784
rect 43684 116750 43718 116784
rect 43752 116750 43786 116784
rect 43820 116750 43854 116784
rect 43888 116750 43922 116784
rect 43956 116750 43990 116784
rect 44024 116750 44058 116784
rect 44092 116750 44126 116784
rect 44160 116750 44194 116784
rect 44228 116750 44262 116784
rect 44296 116750 44330 116784
rect 44364 116750 44398 116784
rect 44432 116750 44466 116784
rect 44500 116750 44534 116784
rect 44568 116750 44602 116784
rect 44636 116750 44670 116784
rect 44704 116750 44738 116784
rect 44772 116750 44806 116784
rect 44840 116750 44874 116784
rect 44908 116750 44942 116784
rect 44976 116750 45010 116784
rect 45044 116750 45078 116784
rect 45112 116750 45146 116784
rect 45180 116750 45214 116784
rect 45248 116750 45282 116784
rect 45316 116750 45350 116784
rect 45384 116750 45418 116784
rect 45452 116750 45486 116784
rect 45520 116750 45554 116784
rect 45588 116750 45622 116784
rect 45656 116750 45690 116784
rect 45724 116750 45758 116784
rect 45792 116750 45826 116784
rect 45860 116750 45894 116784
rect 45928 116750 45962 116784
rect 45996 116750 46030 116784
rect 46064 116750 46098 116784
rect 46132 116750 46166 116784
rect 46200 116750 46234 116784
rect 46268 116750 46302 116784
rect 46336 116750 46370 116784
rect 46404 116750 46438 116784
rect 46472 116750 46506 116784
rect 46540 116750 46574 116784
rect 46608 116750 46642 116784
rect 46676 116750 46710 116784
rect 46744 116750 46778 116784
rect 46812 116750 46846 116784
rect 46880 116750 46914 116784
rect 46948 116750 46982 116784
rect 47016 116750 47050 116784
rect 47084 116750 47118 116784
rect 47152 116750 47250 116784
rect -2416 116730 47250 116750
rect -2416 116697 -2342 116730
rect -2416 116663 -2396 116697
rect -2362 116663 -2342 116697
rect -2416 116629 -2342 116663
rect -2416 116595 -2396 116629
rect -2362 116595 -2342 116629
rect -2416 116561 -2342 116595
rect -2416 116527 -2396 116561
rect -2362 116527 -2342 116561
rect -2416 116493 -2342 116527
rect -2416 116459 -2396 116493
rect -2362 116459 -2342 116493
rect -2416 116425 -2342 116459
rect -2416 116391 -2396 116425
rect -2362 116391 -2342 116425
rect -2416 116357 -2342 116391
rect -2416 116323 -2396 116357
rect -2362 116323 -2342 116357
rect -2416 116289 -2342 116323
rect -2416 116255 -2396 116289
rect -2362 116255 -2342 116289
rect -2416 116221 -2342 116255
rect -2416 116187 -2396 116221
rect -2362 116187 -2342 116221
rect -2416 116153 -2342 116187
rect -2416 116119 -2396 116153
rect -2362 116119 -2342 116153
rect -2416 116085 -2342 116119
rect -2416 116051 -2396 116085
rect -2362 116051 -2342 116085
rect -2416 116017 -2342 116051
rect -2416 115983 -2396 116017
rect -2362 115983 -2342 116017
rect -2416 115949 -2342 115983
rect -2416 115915 -2396 115949
rect -2362 115915 -2342 115949
rect -2416 115881 -2342 115915
rect -2416 115847 -2396 115881
rect -2362 115847 -2342 115881
rect -2416 115813 -2342 115847
rect -2416 115779 -2396 115813
rect -2362 115779 -2342 115813
rect -2416 115745 -2342 115779
rect -2416 115711 -2396 115745
rect -2362 115711 -2342 115745
rect -2416 115677 -2342 115711
rect -2416 115643 -2396 115677
rect -2362 115643 -2342 115677
rect -2416 115609 -2342 115643
rect -2416 115575 -2396 115609
rect -2362 115575 -2342 115609
rect -2416 115541 -2342 115575
rect -2416 115507 -2396 115541
rect -2362 115507 -2342 115541
rect -2416 115473 -2342 115507
rect -2416 115439 -2396 115473
rect -2362 115439 -2342 115473
rect -2416 115405 -2342 115439
rect -2416 115371 -2396 115405
rect -2362 115371 -2342 115405
rect -2416 115337 -2342 115371
rect -2416 115303 -2396 115337
rect -2362 115303 -2342 115337
rect -2416 115269 -2342 115303
rect -2416 115235 -2396 115269
rect -2362 115235 -2342 115269
rect -2416 115201 -2342 115235
rect -2416 115167 -2396 115201
rect -2362 115167 -2342 115201
rect -2416 115133 -2342 115167
rect -2416 115099 -2396 115133
rect -2362 115099 -2342 115133
rect -2416 115065 -2342 115099
rect -2416 115031 -2396 115065
rect -2362 115031 -2342 115065
rect -2416 114997 -2342 115031
rect -2416 114963 -2396 114997
rect -2362 114963 -2342 114997
rect -2416 114929 -2342 114963
rect -2416 114895 -2396 114929
rect -2362 114895 -2342 114929
rect -2416 114861 -2342 114895
rect -2416 114827 -2396 114861
rect -2362 114827 -2342 114861
rect -2416 114793 -2342 114827
rect -2416 114759 -2396 114793
rect -2362 114759 -2342 114793
rect -2416 114725 -2342 114759
rect -2416 114691 -2396 114725
rect -2362 114691 -2342 114725
rect -2416 114657 -2342 114691
rect -2416 114623 -2396 114657
rect -2362 114623 -2342 114657
rect -2416 114589 -2342 114623
rect -2416 114555 -2396 114589
rect -2362 114555 -2342 114589
rect -2416 114521 -2342 114555
rect -2416 114487 -2396 114521
rect -2362 114487 -2342 114521
rect -2416 114453 -2342 114487
rect -2416 114419 -2396 114453
rect -2362 114419 -2342 114453
rect -2416 114385 -2342 114419
rect -2416 114351 -2396 114385
rect -2362 114351 -2342 114385
rect -2416 114317 -2342 114351
rect -2416 114283 -2396 114317
rect -2362 114283 -2342 114317
rect -2416 114249 -2342 114283
rect -2416 114215 -2396 114249
rect -2362 114215 -2342 114249
rect -2416 114181 -2342 114215
rect -2416 114147 -2396 114181
rect -2362 114147 -2342 114181
rect -2416 114113 -2342 114147
rect -2416 114079 -2396 114113
rect -2362 114079 -2342 114113
rect -2416 114045 -2342 114079
rect -2416 114011 -2396 114045
rect -2362 114011 -2342 114045
rect -2416 113977 -2342 114011
rect -2416 113943 -2396 113977
rect -2362 113943 -2342 113977
rect -2416 113909 -2342 113943
rect -2416 113875 -2396 113909
rect -2362 113875 -2342 113909
rect -2416 113841 -2342 113875
rect -2416 113807 -2396 113841
rect -2362 113807 -2342 113841
rect -2416 113773 -2342 113807
rect -2416 113739 -2396 113773
rect -2362 113739 -2342 113773
rect -2416 113705 -2342 113739
rect -2416 113671 -2396 113705
rect -2362 113671 -2342 113705
rect -2416 113637 -2342 113671
rect -2416 113603 -2396 113637
rect -2362 113603 -2342 113637
rect -2416 113569 -2342 113603
rect -2416 113535 -2396 113569
rect -2362 113535 -2342 113569
rect -2416 113501 -2342 113535
rect -2416 113467 -2396 113501
rect -2362 113467 -2342 113501
rect -2416 113433 -2342 113467
rect -2416 113399 -2396 113433
rect -2362 113399 -2342 113433
rect -2416 113365 -2342 113399
rect -2416 113331 -2396 113365
rect -2362 113331 -2342 113365
rect -2416 113297 -2342 113331
rect -2416 113263 -2396 113297
rect -2362 113263 -2342 113297
rect -2416 113229 -2342 113263
rect -2416 113195 -2396 113229
rect -2362 113195 -2342 113229
rect -2416 113161 -2342 113195
rect -2416 113127 -2396 113161
rect -2362 113127 -2342 113161
rect -2416 113093 -2342 113127
rect -2416 113059 -2396 113093
rect -2362 113059 -2342 113093
rect -2416 113025 -2342 113059
rect -2416 112991 -2396 113025
rect -2362 112991 -2342 113025
rect -2416 112957 -2342 112991
rect -2416 112923 -2396 112957
rect -2362 112923 -2342 112957
rect -2416 112889 -2342 112923
rect -2416 112855 -2396 112889
rect -2362 112855 -2342 112889
rect -2416 112821 -2342 112855
rect -2416 112787 -2396 112821
rect -2362 112787 -2342 112821
rect -2416 112753 -2342 112787
rect -2416 112719 -2396 112753
rect -2362 112719 -2342 112753
rect -2416 112685 -2342 112719
rect -2416 112651 -2396 112685
rect -2362 112651 -2342 112685
rect -2416 112617 -2342 112651
rect -2416 112583 -2396 112617
rect -2362 112583 -2342 112617
rect -2416 112549 -2342 112583
rect -2416 112515 -2396 112549
rect -2362 112515 -2342 112549
rect -2416 112481 -2342 112515
rect -2416 112447 -2396 112481
rect -2362 112447 -2342 112481
rect -2416 112413 -2342 112447
rect -2416 112379 -2396 112413
rect -2362 112379 -2342 112413
rect -2416 112345 -2342 112379
rect -2416 112311 -2396 112345
rect -2362 112311 -2342 112345
rect -2416 112277 -2342 112311
rect -2416 112243 -2396 112277
rect -2362 112243 -2342 112277
rect -2416 112209 -2342 112243
rect -2416 112175 -2396 112209
rect -2362 112175 -2342 112209
rect -2416 112141 -2342 112175
rect -2416 112107 -2396 112141
rect -2362 112107 -2342 112141
rect -2416 112073 -2342 112107
rect -2416 112039 -2396 112073
rect -2362 112039 -2342 112073
rect -2416 112005 -2342 112039
rect -2416 111971 -2396 112005
rect -2362 111971 -2342 112005
rect -2416 111937 -2342 111971
rect -2416 111903 -2396 111937
rect -2362 111903 -2342 111937
rect -2416 111869 -2342 111903
rect -2416 111835 -2396 111869
rect -2362 111835 -2342 111869
rect -2416 111801 -2342 111835
rect -2416 111767 -2396 111801
rect -2362 111767 -2342 111801
rect -2416 111733 -2342 111767
rect -2416 111699 -2396 111733
rect -2362 111699 -2342 111733
rect -2416 111665 -2342 111699
rect -2416 111631 -2396 111665
rect -2362 111631 -2342 111665
rect -2416 111597 -2342 111631
rect -2416 111563 -2396 111597
rect -2362 111563 -2342 111597
rect -2416 111529 -2342 111563
rect -2416 111495 -2396 111529
rect -2362 111495 -2342 111529
rect -2416 111461 -2342 111495
rect -2416 111427 -2396 111461
rect -2362 111427 -2342 111461
rect -2416 111393 -2342 111427
rect -2416 111359 -2396 111393
rect -2362 111359 -2342 111393
rect -2416 111325 -2342 111359
rect -2416 111291 -2396 111325
rect -2362 111291 -2342 111325
rect -2416 111257 -2342 111291
rect -2416 111223 -2396 111257
rect -2362 111223 -2342 111257
rect -2416 111189 -2342 111223
rect -2416 111155 -2396 111189
rect -2362 111155 -2342 111189
rect -2416 111121 -2342 111155
rect -2416 111087 -2396 111121
rect -2362 111087 -2342 111121
rect -2416 111053 -2342 111087
rect -2416 111019 -2396 111053
rect -2362 111019 -2342 111053
rect -2416 110985 -2342 111019
rect -2416 110951 -2396 110985
rect -2362 110951 -2342 110985
rect -2416 110917 -2342 110951
rect -2416 110883 -2396 110917
rect -2362 110883 -2342 110917
rect -2416 110849 -2342 110883
rect -2416 110815 -2396 110849
rect -2362 110815 -2342 110849
rect -2416 110781 -2342 110815
rect -2416 110747 -2396 110781
rect -2362 110747 -2342 110781
rect -2416 110713 -2342 110747
rect -2416 110679 -2396 110713
rect -2362 110679 -2342 110713
rect -2416 110645 -2342 110679
rect -2416 110611 -2396 110645
rect -2362 110611 -2342 110645
rect -2416 110577 -2342 110611
rect -2416 110543 -2396 110577
rect -2362 110543 -2342 110577
rect -2416 110509 -2342 110543
rect -2416 110475 -2396 110509
rect -2362 110475 -2342 110509
rect -2416 110441 -2342 110475
rect -2416 110407 -2396 110441
rect -2362 110407 -2342 110441
rect -2416 110373 -2342 110407
rect -2416 110339 -2396 110373
rect -2362 110339 -2342 110373
rect -2416 110305 -2342 110339
rect -2416 110271 -2396 110305
rect -2362 110271 -2342 110305
rect -2416 110237 -2342 110271
rect -2416 110203 -2396 110237
rect -2362 110203 -2342 110237
rect -2416 110169 -2342 110203
rect -2416 110135 -2396 110169
rect -2362 110135 -2342 110169
rect -2416 110101 -2342 110135
rect -2416 110067 -2396 110101
rect -2362 110067 -2342 110101
rect -2416 110033 -2342 110067
rect -2416 109999 -2396 110033
rect -2362 109999 -2342 110033
rect -2416 109965 -2342 109999
rect -2416 109931 -2396 109965
rect -2362 109931 -2342 109965
rect -2416 109897 -2342 109931
rect -2416 109863 -2396 109897
rect -2362 109863 -2342 109897
rect -2416 109829 -2342 109863
rect -2416 109795 -2396 109829
rect -2362 109795 -2342 109829
rect -2416 109761 -2342 109795
rect -2416 109727 -2396 109761
rect -2362 109727 -2342 109761
rect -2416 109693 -2342 109727
rect -2416 109659 -2396 109693
rect -2362 109659 -2342 109693
rect -2416 109625 -2342 109659
rect -2416 109591 -2396 109625
rect -2362 109591 -2342 109625
rect -2416 109557 -2342 109591
rect -2416 109523 -2396 109557
rect -2362 109523 -2342 109557
rect -2416 109489 -2342 109523
rect -2416 109455 -2396 109489
rect -2362 109455 -2342 109489
rect -2416 109421 -2342 109455
rect -2416 109387 -2396 109421
rect -2362 109387 -2342 109421
rect -2416 109353 -2342 109387
rect -2416 109319 -2396 109353
rect -2362 109319 -2342 109353
rect -2416 109285 -2342 109319
rect -2416 109251 -2396 109285
rect -2362 109251 -2342 109285
rect -2416 109217 -2342 109251
rect -2416 109183 -2396 109217
rect -2362 109183 -2342 109217
rect -2416 109149 -2342 109183
rect -2416 109115 -2396 109149
rect -2362 109115 -2342 109149
rect -2416 109081 -2342 109115
rect -2416 109047 -2396 109081
rect -2362 109047 -2342 109081
rect -2416 109013 -2342 109047
rect -2416 108979 -2396 109013
rect -2362 108979 -2342 109013
rect -2416 108945 -2342 108979
rect -2416 108911 -2396 108945
rect -2362 108911 -2342 108945
rect -2416 108877 -2342 108911
rect -2416 108843 -2396 108877
rect -2362 108843 -2342 108877
rect -2416 108809 -2342 108843
rect -2416 108775 -2396 108809
rect -2362 108775 -2342 108809
rect -2416 108741 -2342 108775
rect -2416 108707 -2396 108741
rect -2362 108707 -2342 108741
rect -2416 108673 -2342 108707
rect -2416 108639 -2396 108673
rect -2362 108639 -2342 108673
rect -2416 108605 -2342 108639
rect -2416 108571 -2396 108605
rect -2362 108571 -2342 108605
rect -2416 108537 -2342 108571
rect -2416 108503 -2396 108537
rect -2362 108503 -2342 108537
rect -2416 108469 -2342 108503
rect -2416 108435 -2396 108469
rect -2362 108435 -2342 108469
rect -2416 108401 -2342 108435
rect -2416 108367 -2396 108401
rect -2362 108367 -2342 108401
rect -2416 108333 -2342 108367
rect -2416 108299 -2396 108333
rect -2362 108299 -2342 108333
rect -2416 108265 -2342 108299
rect -2416 108231 -2396 108265
rect -2362 108231 -2342 108265
rect -2416 108197 -2342 108231
rect -2416 108163 -2396 108197
rect -2362 108163 -2342 108197
rect -2416 108129 -2342 108163
rect -2416 108095 -2396 108129
rect -2362 108095 -2342 108129
rect -2416 108061 -2342 108095
rect -2416 108027 -2396 108061
rect -2362 108027 -2342 108061
rect -2416 107993 -2342 108027
rect -2416 107959 -2396 107993
rect -2362 107959 -2342 107993
rect -2416 107925 -2342 107959
rect -2416 107891 -2396 107925
rect -2362 107891 -2342 107925
rect -2416 107857 -2342 107891
rect -2416 107823 -2396 107857
rect -2362 107823 -2342 107857
rect -2416 107789 -2342 107823
rect -2416 107755 -2396 107789
rect -2362 107755 -2342 107789
rect -2416 107721 -2342 107755
rect -2416 107687 -2396 107721
rect -2362 107687 -2342 107721
rect -2416 107653 -2342 107687
rect -2416 107619 -2396 107653
rect -2362 107619 -2342 107653
rect -2416 107585 -2342 107619
rect -2416 107551 -2396 107585
rect -2362 107551 -2342 107585
rect -2416 107517 -2342 107551
rect -2416 107483 -2396 107517
rect -2362 107483 -2342 107517
rect -2416 107449 -2342 107483
rect -2416 107415 -2396 107449
rect -2362 107415 -2342 107449
rect -2416 107381 -2342 107415
rect -2416 107347 -2396 107381
rect -2362 107347 -2342 107381
rect -2416 107313 -2342 107347
rect -2416 107279 -2396 107313
rect -2362 107279 -2342 107313
rect -2416 107245 -2342 107279
rect -2416 107211 -2396 107245
rect -2362 107211 -2342 107245
rect -2416 107177 -2342 107211
rect -2416 107143 -2396 107177
rect -2362 107143 -2342 107177
rect -2416 107109 -2342 107143
rect -2416 107075 -2396 107109
rect -2362 107075 -2342 107109
rect -2416 107041 -2342 107075
rect -2416 107007 -2396 107041
rect -2362 107007 -2342 107041
rect -2416 106973 -2342 107007
rect -2416 106939 -2396 106973
rect -2362 106939 -2342 106973
rect -2416 106905 -2342 106939
rect -2416 106871 -2396 106905
rect -2362 106871 -2342 106905
rect -2416 106837 -2342 106871
rect -2416 106803 -2396 106837
rect -2362 106803 -2342 106837
rect -2416 106769 -2342 106803
rect -2416 106735 -2396 106769
rect -2362 106735 -2342 106769
rect -2416 106701 -2342 106735
rect -2416 106667 -2396 106701
rect -2362 106667 -2342 106701
rect -2416 106633 -2342 106667
rect -2416 106599 -2396 106633
rect -2362 106599 -2342 106633
rect -2416 106565 -2342 106599
rect -2416 106531 -2396 106565
rect -2362 106531 -2342 106565
rect -2416 106497 -2342 106531
rect -2416 106463 -2396 106497
rect -2362 106463 -2342 106497
rect -2416 106429 -2342 106463
rect -2416 106395 -2396 106429
rect -2362 106395 -2342 106429
rect -2416 106361 -2342 106395
rect -2416 106327 -2396 106361
rect -2362 106327 -2342 106361
rect -2416 106293 -2342 106327
rect -2416 106259 -2396 106293
rect -2362 106259 -2342 106293
rect -2416 106225 -2342 106259
rect -2416 106191 -2396 106225
rect -2362 106191 -2342 106225
rect -2416 106157 -2342 106191
rect -2416 106123 -2396 106157
rect -2362 106123 -2342 106157
rect -2416 106089 -2342 106123
rect -2416 106055 -2396 106089
rect -2362 106055 -2342 106089
rect -2416 106021 -2342 106055
rect -2416 105987 -2396 106021
rect -2362 105987 -2342 106021
rect -2416 105953 -2342 105987
rect -2416 105919 -2396 105953
rect -2362 105919 -2342 105953
rect -2416 105885 -2342 105919
rect -2416 105851 -2396 105885
rect -2362 105851 -2342 105885
rect -2416 105817 -2342 105851
rect -2416 105783 -2396 105817
rect -2362 105783 -2342 105817
rect -2416 105749 -2342 105783
rect -2416 105715 -2396 105749
rect -2362 105715 -2342 105749
rect -2416 105681 -2342 105715
rect -2416 105647 -2396 105681
rect -2362 105647 -2342 105681
rect -2416 105613 -2342 105647
rect -2416 105579 -2396 105613
rect -2362 105579 -2342 105613
rect -2416 105545 -2342 105579
rect -2416 105511 -2396 105545
rect -2362 105511 -2342 105545
rect -2416 105477 -2342 105511
rect -2416 105443 -2396 105477
rect -2362 105443 -2342 105477
rect -2416 105409 -2342 105443
rect -2416 105375 -2396 105409
rect -2362 105375 -2342 105409
rect -2416 105341 -2342 105375
rect -2416 105307 -2396 105341
rect -2362 105307 -2342 105341
rect -2416 105273 -2342 105307
rect -2416 105239 -2396 105273
rect -2362 105239 -2342 105273
rect -2416 105205 -2342 105239
rect -2416 105171 -2396 105205
rect -2362 105171 -2342 105205
rect -2416 105137 -2342 105171
rect -2416 105103 -2396 105137
rect -2362 105103 -2342 105137
rect -2416 105069 -2342 105103
rect -2416 105035 -2396 105069
rect -2362 105035 -2342 105069
rect -2416 105001 -2342 105035
rect -2416 104967 -2396 105001
rect -2362 104967 -2342 105001
rect -2416 104933 -2342 104967
rect -2416 104899 -2396 104933
rect -2362 104899 -2342 104933
rect -2416 104865 -2342 104899
rect -2416 104831 -2396 104865
rect -2362 104831 -2342 104865
rect -2416 104797 -2342 104831
rect -2416 104763 -2396 104797
rect -2362 104763 -2342 104797
rect -2416 104729 -2342 104763
rect -2416 104695 -2396 104729
rect -2362 104695 -2342 104729
rect -2416 104661 -2342 104695
rect -2416 104627 -2396 104661
rect -2362 104627 -2342 104661
rect -2416 104593 -2342 104627
rect -2416 104559 -2396 104593
rect -2362 104559 -2342 104593
rect -2416 104525 -2342 104559
rect -2416 104491 -2396 104525
rect -2362 104491 -2342 104525
rect -2416 104457 -2342 104491
rect -2416 104423 -2396 104457
rect -2362 104423 -2342 104457
rect -2416 104389 -2342 104423
rect -2416 104355 -2396 104389
rect -2362 104355 -2342 104389
rect -2416 104321 -2342 104355
rect -2416 104287 -2396 104321
rect -2362 104287 -2342 104321
rect -2416 104253 -2342 104287
rect -2416 104219 -2396 104253
rect -2362 104219 -2342 104253
rect -2416 104185 -2342 104219
rect -2416 104151 -2396 104185
rect -2362 104151 -2342 104185
rect -2416 104117 -2342 104151
rect -2416 104083 -2396 104117
rect -2362 104083 -2342 104117
rect -2416 104049 -2342 104083
rect -2416 104015 -2396 104049
rect -2362 104015 -2342 104049
rect -2416 103981 -2342 104015
rect -2416 103947 -2396 103981
rect -2362 103947 -2342 103981
rect -2416 103913 -2342 103947
rect -2416 103879 -2396 103913
rect -2362 103879 -2342 103913
rect -2416 103845 -2342 103879
rect -2416 103811 -2396 103845
rect -2362 103811 -2342 103845
rect -2416 103777 -2342 103811
rect -2416 103743 -2396 103777
rect -2362 103743 -2342 103777
rect -2416 103709 -2342 103743
rect -2416 103675 -2396 103709
rect -2362 103675 -2342 103709
rect -2416 103641 -2342 103675
rect -2416 103607 -2396 103641
rect -2362 103607 -2342 103641
rect -2416 103573 -2342 103607
rect -2416 103539 -2396 103573
rect -2362 103539 -2342 103573
rect -2416 103505 -2342 103539
rect -2416 103471 -2396 103505
rect -2362 103471 -2342 103505
rect -2416 103437 -2342 103471
rect -2416 103403 -2396 103437
rect -2362 103403 -2342 103437
rect -2416 103369 -2342 103403
rect -2416 103335 -2396 103369
rect -2362 103335 -2342 103369
rect -2416 103301 -2342 103335
rect -2416 103267 -2396 103301
rect -2362 103267 -2342 103301
rect -2416 103233 -2342 103267
rect -2416 103199 -2396 103233
rect -2362 103199 -2342 103233
rect -2416 103165 -2342 103199
rect -2416 103131 -2396 103165
rect -2362 103131 -2342 103165
rect -2416 103097 -2342 103131
rect -2416 103063 -2396 103097
rect -2362 103063 -2342 103097
rect -2416 103029 -2342 103063
rect -2416 102995 -2396 103029
rect -2362 102995 -2342 103029
rect -2416 102961 -2342 102995
rect -2416 102927 -2396 102961
rect -2362 102927 -2342 102961
rect -2416 102893 -2342 102927
rect -2416 102859 -2396 102893
rect -2362 102859 -2342 102893
rect -2416 102825 -2342 102859
rect -2416 102791 -2396 102825
rect -2362 102791 -2342 102825
rect -2416 102757 -2342 102791
rect -2416 102723 -2396 102757
rect -2362 102723 -2342 102757
rect -2416 102689 -2342 102723
rect -2416 102655 -2396 102689
rect -2362 102655 -2342 102689
rect -2416 102621 -2342 102655
rect -2416 102587 -2396 102621
rect -2362 102587 -2342 102621
rect -2416 102553 -2342 102587
rect -2416 102519 -2396 102553
rect -2362 102519 -2342 102553
rect -2416 102485 -2342 102519
rect -2416 102451 -2396 102485
rect -2362 102451 -2342 102485
rect -2416 102417 -2342 102451
rect -2416 102383 -2396 102417
rect -2362 102383 -2342 102417
rect -2416 102349 -2342 102383
rect -2416 102315 -2396 102349
rect -2362 102315 -2342 102349
rect -2416 102281 -2342 102315
rect -2416 102247 -2396 102281
rect -2362 102247 -2342 102281
rect -2416 102213 -2342 102247
rect -2416 102179 -2396 102213
rect -2362 102179 -2342 102213
rect -2416 102145 -2342 102179
rect -2416 102111 -2396 102145
rect -2362 102111 -2342 102145
rect -2416 102077 -2342 102111
rect -2416 102043 -2396 102077
rect -2362 102043 -2342 102077
rect -2416 102009 -2342 102043
rect -2416 101975 -2396 102009
rect -2362 101975 -2342 102009
rect -2416 101941 -2342 101975
rect -2416 101907 -2396 101941
rect -2362 101907 -2342 101941
rect -2416 101873 -2342 101907
rect -2416 101839 -2396 101873
rect -2362 101839 -2342 101873
rect -2416 101805 -2342 101839
rect -2416 101771 -2396 101805
rect -2362 101771 -2342 101805
rect -2416 101737 -2342 101771
rect -2416 101703 -2396 101737
rect -2362 101703 -2342 101737
rect -2416 101669 -2342 101703
rect -2416 101635 -2396 101669
rect -2362 101635 -2342 101669
rect -2416 101601 -2342 101635
rect -2416 101567 -2396 101601
rect -2362 101567 -2342 101601
rect -2416 101533 -2342 101567
rect -2416 101499 -2396 101533
rect -2362 101499 -2342 101533
rect -2416 101465 -2342 101499
rect -2416 101431 -2396 101465
rect -2362 101431 -2342 101465
rect -2416 101397 -2342 101431
rect -2416 101363 -2396 101397
rect -2362 101363 -2342 101397
rect -2416 101329 -2342 101363
rect -2416 101295 -2396 101329
rect -2362 101295 -2342 101329
rect -2416 101261 -2342 101295
rect -2416 101227 -2396 101261
rect -2362 101227 -2342 101261
rect -2416 101193 -2342 101227
rect -2416 101159 -2396 101193
rect -2362 101159 -2342 101193
rect -2416 101125 -2342 101159
rect -2416 101091 -2396 101125
rect -2362 101091 -2342 101125
rect -2416 101057 -2342 101091
rect -2416 101023 -2396 101057
rect -2362 101023 -2342 101057
rect -2416 100989 -2342 101023
rect -2416 100955 -2396 100989
rect -2362 100955 -2342 100989
rect -2416 100923 -2342 100955
rect 47176 116697 47250 116730
rect 47176 116663 47196 116697
rect 47230 116663 47250 116697
rect 47176 116629 47250 116663
rect 47176 116595 47196 116629
rect 47230 116595 47250 116629
rect 47176 116561 47250 116595
rect 47176 116527 47196 116561
rect 47230 116527 47250 116561
rect 47176 116493 47250 116527
rect 47176 116459 47196 116493
rect 47230 116459 47250 116493
rect 47176 116425 47250 116459
rect 47176 116391 47196 116425
rect 47230 116391 47250 116425
rect 47176 116357 47250 116391
rect 47176 116323 47196 116357
rect 47230 116323 47250 116357
rect 47176 116289 47250 116323
rect 47176 116255 47196 116289
rect 47230 116255 47250 116289
rect 47176 116221 47250 116255
rect 47176 116187 47196 116221
rect 47230 116187 47250 116221
rect 47176 116153 47250 116187
rect 47176 116119 47196 116153
rect 47230 116119 47250 116153
rect 47176 116085 47250 116119
rect 47176 116051 47196 116085
rect 47230 116051 47250 116085
rect 47176 116017 47250 116051
rect 47176 115983 47196 116017
rect 47230 115983 47250 116017
rect 47176 115949 47250 115983
rect 47176 115915 47196 115949
rect 47230 115915 47250 115949
rect 47176 115881 47250 115915
rect 47176 115847 47196 115881
rect 47230 115847 47250 115881
rect 47176 115813 47250 115847
rect 47176 115779 47196 115813
rect 47230 115779 47250 115813
rect 47176 115745 47250 115779
rect 47176 115711 47196 115745
rect 47230 115711 47250 115745
rect 47176 115677 47250 115711
rect 47176 115643 47196 115677
rect 47230 115643 47250 115677
rect 47176 115609 47250 115643
rect 47176 115575 47196 115609
rect 47230 115575 47250 115609
rect 47176 115541 47250 115575
rect 47176 115507 47196 115541
rect 47230 115507 47250 115541
rect 47176 115473 47250 115507
rect 47176 115439 47196 115473
rect 47230 115439 47250 115473
rect 47176 115405 47250 115439
rect 47176 115371 47196 115405
rect 47230 115371 47250 115405
rect 47176 115337 47250 115371
rect 47176 115303 47196 115337
rect 47230 115303 47250 115337
rect 47176 115269 47250 115303
rect 47176 115235 47196 115269
rect 47230 115235 47250 115269
rect 47176 115201 47250 115235
rect 47176 115167 47196 115201
rect 47230 115167 47250 115201
rect 47176 115133 47250 115167
rect 47176 115099 47196 115133
rect 47230 115099 47250 115133
rect 47176 115065 47250 115099
rect 47176 115031 47196 115065
rect 47230 115031 47250 115065
rect 47176 114997 47250 115031
rect 47176 114963 47196 114997
rect 47230 114963 47250 114997
rect 47176 114929 47250 114963
rect 47176 114895 47196 114929
rect 47230 114895 47250 114929
rect 47176 114861 47250 114895
rect 47176 114827 47196 114861
rect 47230 114827 47250 114861
rect 47176 114793 47250 114827
rect 47176 114759 47196 114793
rect 47230 114759 47250 114793
rect 47176 114725 47250 114759
rect 47176 114691 47196 114725
rect 47230 114691 47250 114725
rect 47176 114657 47250 114691
rect 47176 114623 47196 114657
rect 47230 114623 47250 114657
rect 47176 114589 47250 114623
rect 47176 114555 47196 114589
rect 47230 114555 47250 114589
rect 47176 114521 47250 114555
rect 47176 114487 47196 114521
rect 47230 114487 47250 114521
rect 47176 114453 47250 114487
rect 47176 114419 47196 114453
rect 47230 114419 47250 114453
rect 47176 114385 47250 114419
rect 47176 114351 47196 114385
rect 47230 114351 47250 114385
rect 47176 114317 47250 114351
rect 47176 114283 47196 114317
rect 47230 114283 47250 114317
rect 47176 114249 47250 114283
rect 47176 114215 47196 114249
rect 47230 114215 47250 114249
rect 47176 114181 47250 114215
rect 47176 114147 47196 114181
rect 47230 114147 47250 114181
rect 47176 114113 47250 114147
rect 47176 114079 47196 114113
rect 47230 114079 47250 114113
rect 47176 114045 47250 114079
rect 47176 114011 47196 114045
rect 47230 114011 47250 114045
rect 47176 113977 47250 114011
rect 47176 113943 47196 113977
rect 47230 113943 47250 113977
rect 47176 113909 47250 113943
rect 47176 113875 47196 113909
rect 47230 113875 47250 113909
rect 47176 113841 47250 113875
rect 47176 113807 47196 113841
rect 47230 113807 47250 113841
rect 47176 113773 47250 113807
rect 47176 113739 47196 113773
rect 47230 113739 47250 113773
rect 47176 113705 47250 113739
rect 47176 113671 47196 113705
rect 47230 113671 47250 113705
rect 47176 113637 47250 113671
rect 47176 113603 47196 113637
rect 47230 113603 47250 113637
rect 47176 113569 47250 113603
rect 47176 113535 47196 113569
rect 47230 113535 47250 113569
rect 47176 113501 47250 113535
rect 47176 113467 47196 113501
rect 47230 113467 47250 113501
rect 47176 113433 47250 113467
rect 47176 113399 47196 113433
rect 47230 113399 47250 113433
rect 47176 113365 47250 113399
rect 47176 113331 47196 113365
rect 47230 113331 47250 113365
rect 47176 113297 47250 113331
rect 47176 113263 47196 113297
rect 47230 113263 47250 113297
rect 47176 113229 47250 113263
rect 47176 113195 47196 113229
rect 47230 113195 47250 113229
rect 47176 113161 47250 113195
rect 47176 113127 47196 113161
rect 47230 113127 47250 113161
rect 47176 113093 47250 113127
rect 47176 113059 47196 113093
rect 47230 113059 47250 113093
rect 47176 113025 47250 113059
rect 47176 112991 47196 113025
rect 47230 112991 47250 113025
rect 47176 112957 47250 112991
rect 47176 112923 47196 112957
rect 47230 112923 47250 112957
rect 47176 112889 47250 112923
rect 47176 112855 47196 112889
rect 47230 112855 47250 112889
rect 47176 112821 47250 112855
rect 47176 112787 47196 112821
rect 47230 112787 47250 112821
rect 47176 112753 47250 112787
rect 47176 112719 47196 112753
rect 47230 112719 47250 112753
rect 47176 112685 47250 112719
rect 47176 112651 47196 112685
rect 47230 112651 47250 112685
rect 47176 112617 47250 112651
rect 47176 112583 47196 112617
rect 47230 112583 47250 112617
rect 47176 112549 47250 112583
rect 47176 112515 47196 112549
rect 47230 112515 47250 112549
rect 47176 112481 47250 112515
rect 47176 112447 47196 112481
rect 47230 112447 47250 112481
rect 47176 112413 47250 112447
rect 47176 112379 47196 112413
rect 47230 112379 47250 112413
rect 47176 112345 47250 112379
rect 47176 112311 47196 112345
rect 47230 112311 47250 112345
rect 47176 112277 47250 112311
rect 47176 112243 47196 112277
rect 47230 112243 47250 112277
rect 47176 112209 47250 112243
rect 47176 112175 47196 112209
rect 47230 112175 47250 112209
rect 47176 112141 47250 112175
rect 47176 112107 47196 112141
rect 47230 112107 47250 112141
rect 47176 112073 47250 112107
rect 47176 112039 47196 112073
rect 47230 112039 47250 112073
rect 47176 112005 47250 112039
rect 47176 111971 47196 112005
rect 47230 111971 47250 112005
rect 47176 111937 47250 111971
rect 47176 111903 47196 111937
rect 47230 111903 47250 111937
rect 47176 111869 47250 111903
rect 47176 111835 47196 111869
rect 47230 111835 47250 111869
rect 47176 111801 47250 111835
rect 47176 111767 47196 111801
rect 47230 111767 47250 111801
rect 47176 111733 47250 111767
rect 47176 111699 47196 111733
rect 47230 111699 47250 111733
rect 47176 111665 47250 111699
rect 47176 111631 47196 111665
rect 47230 111631 47250 111665
rect 47176 111597 47250 111631
rect 47176 111563 47196 111597
rect 47230 111563 47250 111597
rect 47176 111529 47250 111563
rect 47176 111495 47196 111529
rect 47230 111495 47250 111529
rect 47176 111461 47250 111495
rect 47176 111427 47196 111461
rect 47230 111427 47250 111461
rect 47176 111393 47250 111427
rect 47176 111359 47196 111393
rect 47230 111359 47250 111393
rect 47176 111325 47250 111359
rect 47176 111291 47196 111325
rect 47230 111291 47250 111325
rect 47176 111257 47250 111291
rect 47176 111223 47196 111257
rect 47230 111223 47250 111257
rect 47176 111189 47250 111223
rect 47176 111155 47196 111189
rect 47230 111155 47250 111189
rect 47176 111121 47250 111155
rect 47176 111087 47196 111121
rect 47230 111087 47250 111121
rect 47176 111053 47250 111087
rect 47176 111019 47196 111053
rect 47230 111019 47250 111053
rect 47176 110985 47250 111019
rect 47176 110951 47196 110985
rect 47230 110951 47250 110985
rect 47176 110917 47250 110951
rect 47176 110883 47196 110917
rect 47230 110883 47250 110917
rect 47176 110849 47250 110883
rect 47176 110815 47196 110849
rect 47230 110815 47250 110849
rect 47176 110781 47250 110815
rect 47176 110747 47196 110781
rect 47230 110747 47250 110781
rect 47176 110713 47250 110747
rect 47176 110679 47196 110713
rect 47230 110679 47250 110713
rect 47176 110645 47250 110679
rect 47176 110611 47196 110645
rect 47230 110611 47250 110645
rect 47176 110577 47250 110611
rect 47176 110543 47196 110577
rect 47230 110543 47250 110577
rect 47176 110509 47250 110543
rect 47176 110475 47196 110509
rect 47230 110475 47250 110509
rect 47176 110441 47250 110475
rect 47176 110407 47196 110441
rect 47230 110407 47250 110441
rect 47176 110373 47250 110407
rect 47176 110339 47196 110373
rect 47230 110339 47250 110373
rect 47176 110305 47250 110339
rect 47176 110271 47196 110305
rect 47230 110271 47250 110305
rect 47176 110237 47250 110271
rect 47176 110203 47196 110237
rect 47230 110203 47250 110237
rect 47176 110169 47250 110203
rect 47176 110135 47196 110169
rect 47230 110135 47250 110169
rect 47176 110101 47250 110135
rect 47176 110067 47196 110101
rect 47230 110067 47250 110101
rect 47176 110033 47250 110067
rect 47176 109999 47196 110033
rect 47230 109999 47250 110033
rect 47176 109965 47250 109999
rect 47176 109931 47196 109965
rect 47230 109931 47250 109965
rect 47176 109897 47250 109931
rect 47176 109863 47196 109897
rect 47230 109863 47250 109897
rect 47176 109829 47250 109863
rect 47176 109795 47196 109829
rect 47230 109795 47250 109829
rect 47176 109761 47250 109795
rect 47176 109727 47196 109761
rect 47230 109727 47250 109761
rect 47176 109693 47250 109727
rect 47176 109659 47196 109693
rect 47230 109659 47250 109693
rect 47176 109625 47250 109659
rect 47176 109591 47196 109625
rect 47230 109591 47250 109625
rect 47176 109557 47250 109591
rect 47176 109523 47196 109557
rect 47230 109523 47250 109557
rect 47176 109489 47250 109523
rect 47176 109455 47196 109489
rect 47230 109455 47250 109489
rect 47176 109421 47250 109455
rect 47176 109387 47196 109421
rect 47230 109387 47250 109421
rect 47176 109353 47250 109387
rect 47176 109319 47196 109353
rect 47230 109319 47250 109353
rect 47176 109285 47250 109319
rect 47176 109251 47196 109285
rect 47230 109251 47250 109285
rect 47176 109217 47250 109251
rect 47176 109183 47196 109217
rect 47230 109183 47250 109217
rect 47176 109149 47250 109183
rect 47176 109115 47196 109149
rect 47230 109115 47250 109149
rect 47176 109081 47250 109115
rect 47176 109047 47196 109081
rect 47230 109047 47250 109081
rect 47176 109013 47250 109047
rect 47176 108979 47196 109013
rect 47230 108979 47250 109013
rect 47176 108945 47250 108979
rect 47176 108911 47196 108945
rect 47230 108911 47250 108945
rect 47176 108877 47250 108911
rect 47176 108843 47196 108877
rect 47230 108843 47250 108877
rect 47176 108809 47250 108843
rect 47176 108775 47196 108809
rect 47230 108775 47250 108809
rect 47176 108741 47250 108775
rect 47176 108707 47196 108741
rect 47230 108707 47250 108741
rect 47176 108673 47250 108707
rect 47176 108639 47196 108673
rect 47230 108639 47250 108673
rect 47176 108605 47250 108639
rect 47176 108571 47196 108605
rect 47230 108571 47250 108605
rect 47176 108537 47250 108571
rect 47176 108503 47196 108537
rect 47230 108503 47250 108537
rect 47176 108469 47250 108503
rect 47176 108435 47196 108469
rect 47230 108435 47250 108469
rect 47176 108401 47250 108435
rect 47176 108367 47196 108401
rect 47230 108367 47250 108401
rect 47176 108333 47250 108367
rect 47176 108299 47196 108333
rect 47230 108299 47250 108333
rect 47176 108265 47250 108299
rect 47176 108231 47196 108265
rect 47230 108231 47250 108265
rect 47176 108197 47250 108231
rect 47176 108163 47196 108197
rect 47230 108163 47250 108197
rect 47176 108129 47250 108163
rect 47176 108095 47196 108129
rect 47230 108095 47250 108129
rect 47176 108061 47250 108095
rect 47176 108027 47196 108061
rect 47230 108027 47250 108061
rect 47176 107993 47250 108027
rect 47176 107959 47196 107993
rect 47230 107959 47250 107993
rect 47176 107925 47250 107959
rect 47176 107891 47196 107925
rect 47230 107891 47250 107925
rect 47176 107857 47250 107891
rect 47176 107823 47196 107857
rect 47230 107823 47250 107857
rect 47176 107789 47250 107823
rect 47176 107755 47196 107789
rect 47230 107755 47250 107789
rect 47176 107721 47250 107755
rect 47176 107687 47196 107721
rect 47230 107687 47250 107721
rect 47176 107653 47250 107687
rect 47176 107619 47196 107653
rect 47230 107619 47250 107653
rect 47176 107585 47250 107619
rect 47176 107551 47196 107585
rect 47230 107551 47250 107585
rect 47176 107517 47250 107551
rect 47176 107483 47196 107517
rect 47230 107483 47250 107517
rect 47176 107449 47250 107483
rect 47176 107415 47196 107449
rect 47230 107415 47250 107449
rect 47176 107381 47250 107415
rect 47176 107347 47196 107381
rect 47230 107347 47250 107381
rect 47176 107313 47250 107347
rect 47176 107279 47196 107313
rect 47230 107279 47250 107313
rect 47176 107245 47250 107279
rect 47176 107211 47196 107245
rect 47230 107211 47250 107245
rect 47176 107177 47250 107211
rect 47176 107143 47196 107177
rect 47230 107143 47250 107177
rect 47176 107109 47250 107143
rect 47176 107075 47196 107109
rect 47230 107075 47250 107109
rect 47176 107041 47250 107075
rect 47176 107007 47196 107041
rect 47230 107007 47250 107041
rect 47176 106973 47250 107007
rect 47176 106939 47196 106973
rect 47230 106939 47250 106973
rect 47176 106905 47250 106939
rect 47176 106871 47196 106905
rect 47230 106871 47250 106905
rect 47176 106837 47250 106871
rect 47176 106803 47196 106837
rect 47230 106803 47250 106837
rect 47176 106769 47250 106803
rect 47176 106735 47196 106769
rect 47230 106735 47250 106769
rect 47176 106701 47250 106735
rect 47176 106667 47196 106701
rect 47230 106667 47250 106701
rect 47176 106633 47250 106667
rect 47176 106599 47196 106633
rect 47230 106599 47250 106633
rect 47176 106565 47250 106599
rect 47176 106531 47196 106565
rect 47230 106531 47250 106565
rect 47176 106497 47250 106531
rect 47176 106463 47196 106497
rect 47230 106463 47250 106497
rect 47176 106429 47250 106463
rect 47176 106395 47196 106429
rect 47230 106395 47250 106429
rect 47176 106361 47250 106395
rect 47176 106327 47196 106361
rect 47230 106327 47250 106361
rect 47176 106293 47250 106327
rect 47176 106259 47196 106293
rect 47230 106259 47250 106293
rect 47176 106225 47250 106259
rect 47176 106191 47196 106225
rect 47230 106191 47250 106225
rect 47176 106157 47250 106191
rect 47176 106123 47196 106157
rect 47230 106123 47250 106157
rect 47176 106089 47250 106123
rect 47176 106055 47196 106089
rect 47230 106055 47250 106089
rect 47176 106021 47250 106055
rect 47176 105987 47196 106021
rect 47230 105987 47250 106021
rect 47176 105953 47250 105987
rect 47176 105919 47196 105953
rect 47230 105919 47250 105953
rect 47176 105885 47250 105919
rect 47176 105851 47196 105885
rect 47230 105851 47250 105885
rect 47176 105817 47250 105851
rect 47176 105783 47196 105817
rect 47230 105783 47250 105817
rect 47176 105749 47250 105783
rect 47176 105715 47196 105749
rect 47230 105715 47250 105749
rect 47176 105681 47250 105715
rect 47176 105647 47196 105681
rect 47230 105647 47250 105681
rect 47176 105613 47250 105647
rect 47176 105579 47196 105613
rect 47230 105579 47250 105613
rect 47176 105545 47250 105579
rect 47176 105511 47196 105545
rect 47230 105511 47250 105545
rect 47176 105477 47250 105511
rect 47176 105443 47196 105477
rect 47230 105443 47250 105477
rect 47176 105409 47250 105443
rect 47176 105375 47196 105409
rect 47230 105375 47250 105409
rect 47176 105341 47250 105375
rect 47176 105307 47196 105341
rect 47230 105307 47250 105341
rect 47176 105273 47250 105307
rect 47176 105239 47196 105273
rect 47230 105239 47250 105273
rect 47176 105205 47250 105239
rect 47176 105171 47196 105205
rect 47230 105171 47250 105205
rect 47176 105137 47250 105171
rect 47176 105103 47196 105137
rect 47230 105103 47250 105137
rect 47176 105069 47250 105103
rect 47176 105035 47196 105069
rect 47230 105035 47250 105069
rect 47176 105001 47250 105035
rect 47176 104967 47196 105001
rect 47230 104967 47250 105001
rect 47176 104933 47250 104967
rect 47176 104899 47196 104933
rect 47230 104899 47250 104933
rect 47176 104865 47250 104899
rect 47176 104831 47196 104865
rect 47230 104831 47250 104865
rect 47176 104797 47250 104831
rect 47176 104763 47196 104797
rect 47230 104763 47250 104797
rect 47176 104729 47250 104763
rect 47176 104695 47196 104729
rect 47230 104695 47250 104729
rect 47176 104661 47250 104695
rect 47176 104627 47196 104661
rect 47230 104627 47250 104661
rect 47176 104593 47250 104627
rect 47176 104559 47196 104593
rect 47230 104559 47250 104593
rect 47176 104525 47250 104559
rect 47176 104491 47196 104525
rect 47230 104491 47250 104525
rect 47176 104457 47250 104491
rect 47176 104423 47196 104457
rect 47230 104423 47250 104457
rect 47176 104389 47250 104423
rect 47176 104355 47196 104389
rect 47230 104355 47250 104389
rect 47176 104321 47250 104355
rect 47176 104287 47196 104321
rect 47230 104287 47250 104321
rect 47176 104253 47250 104287
rect 47176 104219 47196 104253
rect 47230 104219 47250 104253
rect 47176 104185 47250 104219
rect 47176 104151 47196 104185
rect 47230 104151 47250 104185
rect 47176 104117 47250 104151
rect 47176 104083 47196 104117
rect 47230 104083 47250 104117
rect 47176 104049 47250 104083
rect 47176 104015 47196 104049
rect 47230 104015 47250 104049
rect 47176 103981 47250 104015
rect 47176 103947 47196 103981
rect 47230 103947 47250 103981
rect 47176 103913 47250 103947
rect 47176 103879 47196 103913
rect 47230 103879 47250 103913
rect 47176 103845 47250 103879
rect 47176 103811 47196 103845
rect 47230 103811 47250 103845
rect 47176 103777 47250 103811
rect 47176 103743 47196 103777
rect 47230 103743 47250 103777
rect 47176 103709 47250 103743
rect 47176 103675 47196 103709
rect 47230 103675 47250 103709
rect 47176 103641 47250 103675
rect 47176 103607 47196 103641
rect 47230 103607 47250 103641
rect 47176 103573 47250 103607
rect 47176 103539 47196 103573
rect 47230 103539 47250 103573
rect 47176 103505 47250 103539
rect 47176 103471 47196 103505
rect 47230 103471 47250 103505
rect 47176 103437 47250 103471
rect 47176 103403 47196 103437
rect 47230 103403 47250 103437
rect 47176 103369 47250 103403
rect 47176 103335 47196 103369
rect 47230 103335 47250 103369
rect 47176 103301 47250 103335
rect 47176 103267 47196 103301
rect 47230 103267 47250 103301
rect 47176 103233 47250 103267
rect 47176 103199 47196 103233
rect 47230 103199 47250 103233
rect 47176 103165 47250 103199
rect 47176 103131 47196 103165
rect 47230 103131 47250 103165
rect 47176 103097 47250 103131
rect 47176 103063 47196 103097
rect 47230 103063 47250 103097
rect 47176 103029 47250 103063
rect 47176 102995 47196 103029
rect 47230 102995 47250 103029
rect 47176 102961 47250 102995
rect 47176 102927 47196 102961
rect 47230 102927 47250 102961
rect 47176 102893 47250 102927
rect 47176 102859 47196 102893
rect 47230 102859 47250 102893
rect 47176 102825 47250 102859
rect 47176 102791 47196 102825
rect 47230 102791 47250 102825
rect 47176 102757 47250 102791
rect 47176 102723 47196 102757
rect 47230 102723 47250 102757
rect 47176 102689 47250 102723
rect 47176 102655 47196 102689
rect 47230 102655 47250 102689
rect 47176 102621 47250 102655
rect 47176 102587 47196 102621
rect 47230 102587 47250 102621
rect 47176 102553 47250 102587
rect 47176 102519 47196 102553
rect 47230 102519 47250 102553
rect 47176 102485 47250 102519
rect 47176 102451 47196 102485
rect 47230 102451 47250 102485
rect 47176 102417 47250 102451
rect 47176 102383 47196 102417
rect 47230 102383 47250 102417
rect 47176 102349 47250 102383
rect 47176 102315 47196 102349
rect 47230 102315 47250 102349
rect 47176 102281 47250 102315
rect 47176 102247 47196 102281
rect 47230 102247 47250 102281
rect 47176 102213 47250 102247
rect 47176 102179 47196 102213
rect 47230 102179 47250 102213
rect 47176 102145 47250 102179
rect 47176 102111 47196 102145
rect 47230 102111 47250 102145
rect 47176 102077 47250 102111
rect 47176 102043 47196 102077
rect 47230 102043 47250 102077
rect 47176 102009 47250 102043
rect 47176 101975 47196 102009
rect 47230 101975 47250 102009
rect 47176 101941 47250 101975
rect 47176 101907 47196 101941
rect 47230 101907 47250 101941
rect 47176 101873 47250 101907
rect 47176 101839 47196 101873
rect 47230 101839 47250 101873
rect 47176 101805 47250 101839
rect 47176 101771 47196 101805
rect 47230 101771 47250 101805
rect 47176 101737 47250 101771
rect 47176 101703 47196 101737
rect 47230 101703 47250 101737
rect 47176 101669 47250 101703
rect 47176 101635 47196 101669
rect 47230 101635 47250 101669
rect 47176 101601 47250 101635
rect 47176 101567 47196 101601
rect 47230 101567 47250 101601
rect 47176 101533 47250 101567
rect 47176 101499 47196 101533
rect 47230 101499 47250 101533
rect 47176 101465 47250 101499
rect 47176 101431 47196 101465
rect 47230 101431 47250 101465
rect 47176 101397 47250 101431
rect 47176 101363 47196 101397
rect 47230 101363 47250 101397
rect 47176 101329 47250 101363
rect 47176 101295 47196 101329
rect 47230 101295 47250 101329
rect 47176 101261 47250 101295
rect 47176 101227 47196 101261
rect 47230 101227 47250 101261
rect 47176 101193 47250 101227
rect 47176 101159 47196 101193
rect 47230 101159 47250 101193
rect 47176 101125 47250 101159
rect 47176 101091 47196 101125
rect 47230 101091 47250 101125
rect 47176 101057 47250 101091
rect 47176 101023 47196 101057
rect 47230 101023 47250 101057
rect 47176 100989 47250 101023
rect 47176 100955 47196 100989
rect 47230 100955 47250 100989
rect 47176 100923 47250 100955
rect -2416 100903 47250 100923
rect -2416 100869 -2318 100903
rect -2284 100869 -2250 100903
rect -2216 100869 -2182 100903
rect -2148 100869 -2114 100903
rect -2080 100869 -2046 100903
rect -2012 100869 -1978 100903
rect -1944 100869 -1910 100903
rect -1876 100869 -1842 100903
rect -1808 100869 -1774 100903
rect -1740 100869 -1706 100903
rect -1672 100869 -1638 100903
rect -1604 100869 -1570 100903
rect -1536 100869 -1502 100903
rect -1468 100869 -1434 100903
rect -1400 100869 -1366 100903
rect -1332 100869 -1298 100903
rect -1264 100869 -1230 100903
rect -1196 100869 -1162 100903
rect -1128 100869 -1094 100903
rect -1060 100869 -1026 100903
rect -992 100869 -958 100903
rect -924 100869 -890 100903
rect -856 100869 -822 100903
rect -788 100869 -754 100903
rect -720 100869 -686 100903
rect -652 100869 -618 100903
rect -584 100869 -550 100903
rect -516 100869 -482 100903
rect -448 100869 -414 100903
rect -380 100869 -346 100903
rect -312 100869 -278 100903
rect -244 100869 -210 100903
rect -176 100869 -142 100903
rect -108 100869 -74 100903
rect -40 100869 -6 100903
rect 28 100869 62 100903
rect 96 100869 130 100903
rect 164 100869 198 100903
rect 232 100869 266 100903
rect 300 100869 334 100903
rect 368 100869 402 100903
rect 436 100869 470 100903
rect 504 100869 538 100903
rect 572 100869 606 100903
rect 640 100869 674 100903
rect 708 100869 742 100903
rect 776 100869 810 100903
rect 844 100869 878 100903
rect 912 100869 946 100903
rect 980 100869 1014 100903
rect 1048 100869 1082 100903
rect 1116 100869 1150 100903
rect 1184 100869 1218 100903
rect 1252 100869 1286 100903
rect 1320 100869 1354 100903
rect 1388 100869 1422 100903
rect 1456 100869 1490 100903
rect 1524 100869 1558 100903
rect 1592 100869 1626 100903
rect 1660 100869 1694 100903
rect 1728 100869 1762 100903
rect 1796 100869 1830 100903
rect 1864 100869 1898 100903
rect 1932 100869 1966 100903
rect 2000 100869 2034 100903
rect 2068 100869 2102 100903
rect 2136 100869 2170 100903
rect 2204 100869 2238 100903
rect 2272 100869 2306 100903
rect 2340 100869 2374 100903
rect 2408 100869 2442 100903
rect 2476 100869 2510 100903
rect 2544 100869 2578 100903
rect 2612 100869 2646 100903
rect 2680 100869 2714 100903
rect 2748 100869 2782 100903
rect 2816 100869 2850 100903
rect 2884 100869 2918 100903
rect 2952 100869 2986 100903
rect 3020 100869 3054 100903
rect 3088 100869 3122 100903
rect 3156 100869 3190 100903
rect 3224 100869 3258 100903
rect 3292 100869 3326 100903
rect 3360 100869 3394 100903
rect 3428 100869 3462 100903
rect 3496 100869 3530 100903
rect 3564 100869 3598 100903
rect 3632 100869 3666 100903
rect 3700 100869 3734 100903
rect 3768 100869 3802 100903
rect 3836 100869 3870 100903
rect 3904 100869 3938 100903
rect 3972 100869 4006 100903
rect 4040 100869 4074 100903
rect 4108 100869 4142 100903
rect 4176 100869 4210 100903
rect 4244 100869 4278 100903
rect 4312 100869 4346 100903
rect 4380 100869 4414 100903
rect 4448 100869 4482 100903
rect 4516 100869 4550 100903
rect 4584 100869 4618 100903
rect 4652 100869 4686 100903
rect 4720 100869 4754 100903
rect 4788 100869 4822 100903
rect 4856 100869 4890 100903
rect 4924 100869 4958 100903
rect 4992 100869 5026 100903
rect 5060 100869 5094 100903
rect 5128 100869 5162 100903
rect 5196 100869 5230 100903
rect 5264 100869 5298 100903
rect 5332 100869 5366 100903
rect 5400 100869 5434 100903
rect 5468 100869 5502 100903
rect 5536 100869 5570 100903
rect 5604 100869 5638 100903
rect 5672 100869 5706 100903
rect 5740 100869 5774 100903
rect 5808 100869 5842 100903
rect 5876 100869 5910 100903
rect 5944 100869 5978 100903
rect 6012 100869 6046 100903
rect 6080 100869 6114 100903
rect 6148 100869 6182 100903
rect 6216 100869 6250 100903
rect 6284 100869 6318 100903
rect 6352 100869 6386 100903
rect 6420 100869 6454 100903
rect 6488 100869 6522 100903
rect 6556 100869 6590 100903
rect 6624 100869 6658 100903
rect 6692 100869 6726 100903
rect 6760 100869 6794 100903
rect 6828 100869 6862 100903
rect 6896 100869 6930 100903
rect 6964 100869 6998 100903
rect 7032 100869 7066 100903
rect 7100 100869 7134 100903
rect 7168 100869 7202 100903
rect 7236 100869 7270 100903
rect 7304 100869 7338 100903
rect 7372 100869 7406 100903
rect 7440 100869 7474 100903
rect 7508 100869 7542 100903
rect 7576 100869 7610 100903
rect 7644 100869 7678 100903
rect 7712 100869 7746 100903
rect 7780 100869 7814 100903
rect 7848 100869 7882 100903
rect 7916 100869 7950 100903
rect 7984 100869 8018 100903
rect 8052 100869 8086 100903
rect 8120 100869 8154 100903
rect 8188 100869 8222 100903
rect 8256 100869 8290 100903
rect 8324 100869 8358 100903
rect 8392 100869 8426 100903
rect 8460 100869 8494 100903
rect 8528 100869 8562 100903
rect 8596 100869 8630 100903
rect 8664 100869 8698 100903
rect 8732 100869 8766 100903
rect 8800 100869 8834 100903
rect 8868 100869 8902 100903
rect 8936 100869 8970 100903
rect 9004 100869 9038 100903
rect 9072 100869 9106 100903
rect 9140 100869 9174 100903
rect 9208 100869 9242 100903
rect 9276 100869 9310 100903
rect 9344 100869 9378 100903
rect 9412 100869 9446 100903
rect 9480 100869 9514 100903
rect 9548 100869 9582 100903
rect 9616 100869 9650 100903
rect 9684 100869 9718 100903
rect 9752 100869 9786 100903
rect 9820 100869 9854 100903
rect 9888 100869 9922 100903
rect 9956 100869 9990 100903
rect 10024 100869 10058 100903
rect 10092 100869 10126 100903
rect 10160 100869 10194 100903
rect 10228 100869 10262 100903
rect 10296 100869 10330 100903
rect 10364 100869 10398 100903
rect 10432 100869 10466 100903
rect 10500 100869 10534 100903
rect 10568 100869 10602 100903
rect 10636 100869 10670 100903
rect 10704 100869 10738 100903
rect 10772 100869 10806 100903
rect 10840 100869 10874 100903
rect 10908 100869 10942 100903
rect 10976 100869 11010 100903
rect 11044 100869 11078 100903
rect 11112 100869 11146 100903
rect 11180 100869 11214 100903
rect 11248 100869 11282 100903
rect 11316 100869 11350 100903
rect 11384 100869 11418 100903
rect 11452 100869 11486 100903
rect 11520 100869 11554 100903
rect 11588 100869 11622 100903
rect 11656 100869 11690 100903
rect 11724 100869 11758 100903
rect 11792 100869 11826 100903
rect 11860 100869 11894 100903
rect 11928 100869 11962 100903
rect 11996 100869 12030 100903
rect 12064 100869 12098 100903
rect 12132 100869 12166 100903
rect 12200 100869 12234 100903
rect 12268 100869 12302 100903
rect 12336 100869 12370 100903
rect 12404 100869 12438 100903
rect 12472 100869 12506 100903
rect 12540 100869 12574 100903
rect 12608 100869 12642 100903
rect 12676 100869 12710 100903
rect 12744 100869 12778 100903
rect 12812 100869 12846 100903
rect 12880 100869 12914 100903
rect 12948 100869 12982 100903
rect 13016 100869 13050 100903
rect 13084 100869 13118 100903
rect 13152 100869 13186 100903
rect 13220 100869 13254 100903
rect 13288 100869 13322 100903
rect 13356 100869 13390 100903
rect 13424 100869 13458 100903
rect 13492 100869 13526 100903
rect 13560 100869 13594 100903
rect 13628 100869 13662 100903
rect 13696 100869 13730 100903
rect 13764 100869 13798 100903
rect 13832 100869 13866 100903
rect 13900 100869 13934 100903
rect 13968 100869 14002 100903
rect 14036 100869 14070 100903
rect 14104 100869 14138 100903
rect 14172 100869 14206 100903
rect 14240 100869 14274 100903
rect 14308 100869 14342 100903
rect 14376 100869 14410 100903
rect 14444 100869 14478 100903
rect 14512 100869 14546 100903
rect 14580 100869 14614 100903
rect 14648 100869 14682 100903
rect 14716 100869 14750 100903
rect 14784 100869 14818 100903
rect 14852 100869 14886 100903
rect 14920 100869 14954 100903
rect 14988 100869 15022 100903
rect 15056 100869 15090 100903
rect 15124 100869 15158 100903
rect 15192 100869 15226 100903
rect 15260 100869 15294 100903
rect 15328 100869 15362 100903
rect 15396 100869 15430 100903
rect 15464 100869 15498 100903
rect 15532 100869 15566 100903
rect 15600 100869 15634 100903
rect 15668 100869 15702 100903
rect 15736 100869 15770 100903
rect 15804 100869 15838 100903
rect 15872 100869 15906 100903
rect 15940 100869 15974 100903
rect 16008 100869 16042 100903
rect 16076 100869 16110 100903
rect 16144 100869 16178 100903
rect 16212 100869 16246 100903
rect 16280 100869 16314 100903
rect 16348 100869 16382 100903
rect 16416 100869 16450 100903
rect 16484 100869 16518 100903
rect 16552 100869 16586 100903
rect 16620 100869 16654 100903
rect 16688 100869 16722 100903
rect 16756 100869 16790 100903
rect 16824 100869 16858 100903
rect 16892 100869 16926 100903
rect 16960 100869 16994 100903
rect 17028 100869 17062 100903
rect 17096 100869 17130 100903
rect 17164 100869 17198 100903
rect 17232 100869 17266 100903
rect 17300 100869 17334 100903
rect 17368 100869 17402 100903
rect 17436 100869 17470 100903
rect 17504 100869 17538 100903
rect 17572 100869 17606 100903
rect 17640 100869 17674 100903
rect 17708 100869 17742 100903
rect 17776 100869 17810 100903
rect 17844 100869 17878 100903
rect 17912 100869 17946 100903
rect 17980 100869 18014 100903
rect 18048 100869 18082 100903
rect 18116 100869 18150 100903
rect 18184 100869 18218 100903
rect 18252 100869 18286 100903
rect 18320 100869 18354 100903
rect 18388 100869 18422 100903
rect 18456 100869 18490 100903
rect 18524 100869 18558 100903
rect 18592 100869 18626 100903
rect 18660 100869 18694 100903
rect 18728 100869 18762 100903
rect 18796 100869 18830 100903
rect 18864 100869 18898 100903
rect 18932 100869 18966 100903
rect 19000 100869 19034 100903
rect 19068 100869 19102 100903
rect 19136 100869 19170 100903
rect 19204 100869 19238 100903
rect 19272 100869 19306 100903
rect 19340 100869 19374 100903
rect 19408 100869 19442 100903
rect 19476 100869 19510 100903
rect 19544 100869 19578 100903
rect 19612 100869 19646 100903
rect 19680 100869 19714 100903
rect 19748 100869 19782 100903
rect 19816 100869 19850 100903
rect 19884 100869 19918 100903
rect 19952 100869 19986 100903
rect 20020 100869 20054 100903
rect 20088 100869 20122 100903
rect 20156 100869 20190 100903
rect 20224 100869 20258 100903
rect 20292 100869 20326 100903
rect 20360 100869 20394 100903
rect 20428 100869 20462 100903
rect 20496 100869 20530 100903
rect 20564 100869 20598 100903
rect 20632 100869 20666 100903
rect 20700 100869 20734 100903
rect 20768 100869 20802 100903
rect 20836 100869 20870 100903
rect 20904 100869 20938 100903
rect 20972 100869 21006 100903
rect 21040 100869 21074 100903
rect 21108 100869 21142 100903
rect 21176 100869 21210 100903
rect 21244 100869 21278 100903
rect 21312 100869 21346 100903
rect 21380 100869 21414 100903
rect 21448 100869 21482 100903
rect 21516 100869 21550 100903
rect 21584 100869 21618 100903
rect 21652 100869 21686 100903
rect 21720 100869 21754 100903
rect 21788 100869 21822 100903
rect 21856 100869 21890 100903
rect 21924 100869 21958 100903
rect 21992 100869 22026 100903
rect 22060 100869 22094 100903
rect 22128 100869 22162 100903
rect 22196 100869 22230 100903
rect 22264 100869 22298 100903
rect 22332 100869 22366 100903
rect 22400 100869 22434 100903
rect 22468 100869 22502 100903
rect 22536 100869 22570 100903
rect 22604 100869 22638 100903
rect 22672 100869 22706 100903
rect 22740 100869 22774 100903
rect 22808 100869 22842 100903
rect 22876 100869 22910 100903
rect 22944 100869 22978 100903
rect 23012 100869 23046 100903
rect 23080 100869 23114 100903
rect 23148 100869 23182 100903
rect 23216 100869 23250 100903
rect 23284 100869 23318 100903
rect 23352 100869 23386 100903
rect 23420 100869 23454 100903
rect 23488 100869 23522 100903
rect 23556 100869 23590 100903
rect 23624 100869 23658 100903
rect 23692 100869 23726 100903
rect 23760 100869 23794 100903
rect 23828 100869 23862 100903
rect 23896 100869 23930 100903
rect 23964 100869 23998 100903
rect 24032 100869 24066 100903
rect 24100 100869 24134 100903
rect 24168 100869 24202 100903
rect 24236 100869 24270 100903
rect 24304 100869 24338 100903
rect 24372 100869 24406 100903
rect 24440 100869 24474 100903
rect 24508 100869 24542 100903
rect 24576 100869 24610 100903
rect 24644 100869 24678 100903
rect 24712 100869 24746 100903
rect 24780 100869 24814 100903
rect 24848 100869 24882 100903
rect 24916 100869 24950 100903
rect 24984 100869 25018 100903
rect 25052 100869 25086 100903
rect 25120 100869 25154 100903
rect 25188 100869 25222 100903
rect 25256 100869 25290 100903
rect 25324 100869 25358 100903
rect 25392 100869 25426 100903
rect 25460 100869 25494 100903
rect 25528 100869 25562 100903
rect 25596 100869 25630 100903
rect 25664 100869 25698 100903
rect 25732 100869 25766 100903
rect 25800 100869 25834 100903
rect 25868 100869 25902 100903
rect 25936 100869 25970 100903
rect 26004 100869 26038 100903
rect 26072 100869 26106 100903
rect 26140 100869 26174 100903
rect 26208 100869 26242 100903
rect 26276 100869 26310 100903
rect 26344 100869 26378 100903
rect 26412 100869 26446 100903
rect 26480 100869 26514 100903
rect 26548 100869 26582 100903
rect 26616 100869 26650 100903
rect 26684 100869 26718 100903
rect 26752 100869 26786 100903
rect 26820 100869 26854 100903
rect 26888 100869 26922 100903
rect 26956 100869 26990 100903
rect 27024 100869 27058 100903
rect 27092 100869 27126 100903
rect 27160 100869 27194 100903
rect 27228 100869 27262 100903
rect 27296 100869 27330 100903
rect 27364 100869 27398 100903
rect 27432 100869 27466 100903
rect 27500 100869 27534 100903
rect 27568 100869 27602 100903
rect 27636 100869 27670 100903
rect 27704 100869 27738 100903
rect 27772 100869 27806 100903
rect 27840 100869 27874 100903
rect 27908 100869 27942 100903
rect 27976 100869 28010 100903
rect 28044 100869 28078 100903
rect 28112 100869 28146 100903
rect 28180 100869 28214 100903
rect 28248 100869 28282 100903
rect 28316 100869 28350 100903
rect 28384 100869 28418 100903
rect 28452 100869 28486 100903
rect 28520 100869 28554 100903
rect 28588 100869 28622 100903
rect 28656 100869 28690 100903
rect 28724 100869 28758 100903
rect 28792 100869 28826 100903
rect 28860 100869 28894 100903
rect 28928 100869 28962 100903
rect 28996 100869 29030 100903
rect 29064 100869 29098 100903
rect 29132 100869 29166 100903
rect 29200 100869 29234 100903
rect 29268 100869 29302 100903
rect 29336 100869 29370 100903
rect 29404 100869 29438 100903
rect 29472 100869 29506 100903
rect 29540 100869 29574 100903
rect 29608 100869 29642 100903
rect 29676 100869 29710 100903
rect 29744 100869 29778 100903
rect 29812 100869 29846 100903
rect 29880 100869 29914 100903
rect 29948 100869 29982 100903
rect 30016 100869 30050 100903
rect 30084 100869 30118 100903
rect 30152 100869 30186 100903
rect 30220 100869 30254 100903
rect 30288 100869 30322 100903
rect 30356 100869 30390 100903
rect 30424 100869 30458 100903
rect 30492 100869 30526 100903
rect 30560 100869 30594 100903
rect 30628 100869 30662 100903
rect 30696 100869 30730 100903
rect 30764 100869 30798 100903
rect 30832 100869 30866 100903
rect 30900 100869 30934 100903
rect 30968 100869 31002 100903
rect 31036 100869 31070 100903
rect 31104 100869 31138 100903
rect 31172 100869 31206 100903
rect 31240 100869 31274 100903
rect 31308 100869 31342 100903
rect 31376 100869 31410 100903
rect 31444 100869 31478 100903
rect 31512 100869 31546 100903
rect 31580 100869 31614 100903
rect 31648 100869 31682 100903
rect 31716 100869 31750 100903
rect 31784 100869 31818 100903
rect 31852 100869 31886 100903
rect 31920 100869 31954 100903
rect 31988 100869 32022 100903
rect 32056 100869 32090 100903
rect 32124 100869 32158 100903
rect 32192 100869 32226 100903
rect 32260 100869 32294 100903
rect 32328 100869 32362 100903
rect 32396 100869 32430 100903
rect 32464 100869 32498 100903
rect 32532 100869 32566 100903
rect 32600 100869 32634 100903
rect 32668 100869 32702 100903
rect 32736 100869 32770 100903
rect 32804 100869 32838 100903
rect 32872 100869 32906 100903
rect 32940 100869 32974 100903
rect 33008 100869 33042 100903
rect 33076 100869 33110 100903
rect 33144 100869 33178 100903
rect 33212 100869 33246 100903
rect 33280 100869 33314 100903
rect 33348 100869 33382 100903
rect 33416 100869 33450 100903
rect 33484 100869 33518 100903
rect 33552 100869 33586 100903
rect 33620 100869 33654 100903
rect 33688 100869 33722 100903
rect 33756 100869 33790 100903
rect 33824 100869 33858 100903
rect 33892 100869 33926 100903
rect 33960 100869 33994 100903
rect 34028 100869 34062 100903
rect 34096 100869 34130 100903
rect 34164 100869 34198 100903
rect 34232 100869 34266 100903
rect 34300 100869 34334 100903
rect 34368 100869 34402 100903
rect 34436 100869 34470 100903
rect 34504 100869 34538 100903
rect 34572 100869 34606 100903
rect 34640 100869 34674 100903
rect 34708 100869 34742 100903
rect 34776 100869 34810 100903
rect 34844 100869 34878 100903
rect 34912 100869 34946 100903
rect 34980 100869 35014 100903
rect 35048 100869 35082 100903
rect 35116 100869 35150 100903
rect 35184 100869 35218 100903
rect 35252 100869 35286 100903
rect 35320 100869 35354 100903
rect 35388 100869 35422 100903
rect 35456 100869 35490 100903
rect 35524 100869 35558 100903
rect 35592 100869 35626 100903
rect 35660 100869 35694 100903
rect 35728 100869 35762 100903
rect 35796 100869 35830 100903
rect 35864 100869 35898 100903
rect 35932 100869 35966 100903
rect 36000 100869 36034 100903
rect 36068 100869 36102 100903
rect 36136 100869 36170 100903
rect 36204 100869 36238 100903
rect 36272 100869 36306 100903
rect 36340 100869 36374 100903
rect 36408 100869 36442 100903
rect 36476 100869 36510 100903
rect 36544 100869 36578 100903
rect 36612 100869 36646 100903
rect 36680 100869 36714 100903
rect 36748 100869 36782 100903
rect 36816 100869 36850 100903
rect 36884 100869 36918 100903
rect 36952 100869 36986 100903
rect 37020 100869 37054 100903
rect 37088 100869 37122 100903
rect 37156 100869 37190 100903
rect 37224 100869 37258 100903
rect 37292 100869 37326 100903
rect 37360 100869 37394 100903
rect 37428 100869 37462 100903
rect 37496 100869 37530 100903
rect 37564 100869 37598 100903
rect 37632 100869 37666 100903
rect 37700 100869 37734 100903
rect 37768 100869 37802 100903
rect 37836 100869 37870 100903
rect 37904 100869 37938 100903
rect 37972 100869 38006 100903
rect 38040 100869 38074 100903
rect 38108 100869 38142 100903
rect 38176 100869 38210 100903
rect 38244 100869 38278 100903
rect 38312 100869 38346 100903
rect 38380 100869 38414 100903
rect 38448 100869 38482 100903
rect 38516 100869 38550 100903
rect 38584 100869 38618 100903
rect 38652 100869 38686 100903
rect 38720 100869 38754 100903
rect 38788 100869 38822 100903
rect 38856 100869 38890 100903
rect 38924 100869 38958 100903
rect 38992 100869 39026 100903
rect 39060 100869 39094 100903
rect 39128 100869 39162 100903
rect 39196 100869 39230 100903
rect 39264 100869 39298 100903
rect 39332 100869 39366 100903
rect 39400 100869 39434 100903
rect 39468 100869 39502 100903
rect 39536 100869 39570 100903
rect 39604 100869 39638 100903
rect 39672 100869 39706 100903
rect 39740 100869 39774 100903
rect 39808 100869 39842 100903
rect 39876 100869 39910 100903
rect 39944 100869 39978 100903
rect 40012 100869 40046 100903
rect 40080 100869 40114 100903
rect 40148 100869 40182 100903
rect 40216 100869 40250 100903
rect 40284 100869 40318 100903
rect 40352 100869 40386 100903
rect 40420 100869 40454 100903
rect 40488 100869 40522 100903
rect 40556 100869 40590 100903
rect 40624 100869 40658 100903
rect 40692 100869 40726 100903
rect 40760 100869 40794 100903
rect 40828 100869 40862 100903
rect 40896 100869 40930 100903
rect 40964 100869 40998 100903
rect 41032 100869 41066 100903
rect 41100 100869 41134 100903
rect 41168 100869 41202 100903
rect 41236 100869 41270 100903
rect 41304 100869 41338 100903
rect 41372 100869 41406 100903
rect 41440 100869 41474 100903
rect 41508 100869 41542 100903
rect 41576 100869 41610 100903
rect 41644 100869 41678 100903
rect 41712 100869 41746 100903
rect 41780 100869 41814 100903
rect 41848 100869 41882 100903
rect 41916 100869 41950 100903
rect 41984 100869 42018 100903
rect 42052 100869 42086 100903
rect 42120 100869 42154 100903
rect 42188 100869 42222 100903
rect 42256 100869 42290 100903
rect 42324 100869 42358 100903
rect 42392 100869 42426 100903
rect 42460 100869 42494 100903
rect 42528 100869 42562 100903
rect 42596 100869 42630 100903
rect 42664 100869 42698 100903
rect 42732 100869 42766 100903
rect 42800 100869 42834 100903
rect 42868 100869 42902 100903
rect 42936 100869 42970 100903
rect 43004 100869 43038 100903
rect 43072 100869 43106 100903
rect 43140 100869 43174 100903
rect 43208 100869 43242 100903
rect 43276 100869 43310 100903
rect 43344 100869 43378 100903
rect 43412 100869 43446 100903
rect 43480 100869 43514 100903
rect 43548 100869 43582 100903
rect 43616 100869 43650 100903
rect 43684 100869 43718 100903
rect 43752 100869 43786 100903
rect 43820 100869 43854 100903
rect 43888 100869 43922 100903
rect 43956 100869 43990 100903
rect 44024 100869 44058 100903
rect 44092 100869 44126 100903
rect 44160 100869 44194 100903
rect 44228 100869 44262 100903
rect 44296 100869 44330 100903
rect 44364 100869 44398 100903
rect 44432 100869 44466 100903
rect 44500 100869 44534 100903
rect 44568 100869 44602 100903
rect 44636 100869 44670 100903
rect 44704 100869 44738 100903
rect 44772 100869 44806 100903
rect 44840 100869 44874 100903
rect 44908 100869 44942 100903
rect 44976 100869 45010 100903
rect 45044 100869 45078 100903
rect 45112 100869 45146 100903
rect 45180 100869 45214 100903
rect 45248 100869 45282 100903
rect 45316 100869 45350 100903
rect 45384 100869 45418 100903
rect 45452 100869 45486 100903
rect 45520 100869 45554 100903
rect 45588 100869 45622 100903
rect 45656 100869 45690 100903
rect 45724 100869 45758 100903
rect 45792 100869 45826 100903
rect 45860 100869 45894 100903
rect 45928 100869 45962 100903
rect 45996 100869 46030 100903
rect 46064 100869 46098 100903
rect 46132 100869 46166 100903
rect 46200 100869 46234 100903
rect 46268 100869 46302 100903
rect 46336 100869 46370 100903
rect 46404 100869 46438 100903
rect 46472 100869 46506 100903
rect 46540 100869 46574 100903
rect 46608 100869 46642 100903
rect 46676 100869 46710 100903
rect 46744 100869 46778 100903
rect 46812 100869 46846 100903
rect 46880 100869 46914 100903
rect 46948 100869 46982 100903
rect 47016 100869 47050 100903
rect 47084 100869 47118 100903
rect 47152 100869 47250 100903
rect -2416 100849 47250 100869
rect -10719 76144 -3664 76164
rect -10719 76110 -10609 76144
rect -10575 76110 -10541 76144
rect -10507 76110 -10473 76144
rect -10439 76110 -10405 76144
rect -10371 76110 -10337 76144
rect -10303 76110 -10269 76144
rect -10235 76110 -10201 76144
rect -10167 76110 -10133 76144
rect -10099 76110 -10065 76144
rect -10031 76110 -9997 76144
rect -9963 76110 -9929 76144
rect -9895 76110 -9861 76144
rect -9827 76110 -9793 76144
rect -9759 76110 -9725 76144
rect -9691 76110 -9657 76144
rect -9623 76110 -9589 76144
rect -9555 76110 -9521 76144
rect -9487 76110 -9453 76144
rect -9419 76110 -9385 76144
rect -9351 76110 -9317 76144
rect -9283 76110 -9249 76144
rect -9215 76110 -9181 76144
rect -9147 76110 -9113 76144
rect -9079 76110 -9045 76144
rect -9011 76110 -8977 76144
rect -8943 76110 -8909 76144
rect -8875 76110 -8841 76144
rect -8807 76110 -8773 76144
rect -8739 76110 -8705 76144
rect -8671 76110 -8637 76144
rect -8603 76110 -8569 76144
rect -8535 76110 -8501 76144
rect -8467 76110 -8433 76144
rect -8399 76110 -8365 76144
rect -8331 76110 -8297 76144
rect -8263 76110 -8229 76144
rect -8195 76110 -8161 76144
rect -8127 76110 -8093 76144
rect -8059 76110 -8025 76144
rect -7991 76110 -7957 76144
rect -7923 76110 -7889 76144
rect -7855 76110 -7821 76144
rect -7787 76110 -7753 76144
rect -7719 76110 -7685 76144
rect -7651 76110 -7617 76144
rect -7583 76110 -7549 76144
rect -7515 76110 -7481 76144
rect -7447 76110 -7413 76144
rect -7379 76110 -7345 76144
rect -7311 76110 -7277 76144
rect -7243 76110 -7209 76144
rect -7175 76110 -7141 76144
rect -7107 76110 -7073 76144
rect -7039 76110 -7005 76144
rect -6971 76110 -6937 76144
rect -6903 76110 -6869 76144
rect -6835 76110 -6801 76144
rect -6767 76110 -6733 76144
rect -6699 76110 -6665 76144
rect -6631 76110 -6597 76144
rect -6563 76110 -6529 76144
rect -6495 76110 -6461 76144
rect -6427 76110 -6393 76144
rect -6359 76110 -6325 76144
rect -6291 76110 -6257 76144
rect -6223 76110 -6189 76144
rect -6155 76110 -6121 76144
rect -6087 76110 -6053 76144
rect -6019 76110 -5985 76144
rect -5951 76110 -5917 76144
rect -5883 76110 -5849 76144
rect -5815 76110 -5781 76144
rect -5747 76110 -5713 76144
rect -5679 76110 -5645 76144
rect -5611 76110 -5577 76144
rect -5543 76110 -5509 76144
rect -5475 76110 -5441 76144
rect -5407 76110 -5373 76144
rect -5339 76110 -5305 76144
rect -5271 76110 -5237 76144
rect -5203 76110 -5169 76144
rect -5135 76110 -5101 76144
rect -5067 76110 -5033 76144
rect -4999 76110 -4965 76144
rect -4931 76110 -4897 76144
rect -4863 76110 -4829 76144
rect -4795 76110 -4761 76144
rect -4727 76110 -4693 76144
rect -4659 76110 -4625 76144
rect -4591 76110 -4557 76144
rect -4523 76110 -4489 76144
rect -4455 76110 -4421 76144
rect -4387 76110 -4353 76144
rect -4319 76110 -4285 76144
rect -4251 76110 -4217 76144
rect -4183 76110 -4149 76144
rect -4115 76110 -4081 76144
rect -4047 76110 -4013 76144
rect -3979 76110 -3945 76144
rect -3911 76110 -3877 76144
rect -3843 76110 -3809 76144
rect -3775 76110 -3664 76144
rect -10719 76090 -3664 76110
rect -10719 76084 -10645 76090
rect -10719 76050 -10699 76084
rect -10665 76050 -10645 76084
rect -10719 76016 -10645 76050
rect -10719 75982 -10699 76016
rect -10665 75982 -10645 76016
rect -10719 75948 -10645 75982
rect -10719 75914 -10699 75948
rect -10665 75914 -10645 75948
rect -10719 75880 -10645 75914
rect -10719 75846 -10699 75880
rect -10665 75846 -10645 75880
rect -10719 75812 -10645 75846
rect -10719 75778 -10699 75812
rect -10665 75778 -10645 75812
rect -10719 75744 -10645 75778
rect -10719 75710 -10699 75744
rect -10665 75710 -10645 75744
rect -10719 75676 -10645 75710
rect -10719 75642 -10699 75676
rect -10665 75642 -10645 75676
rect -10719 75608 -10645 75642
rect -10719 75574 -10699 75608
rect -10665 75574 -10645 75608
rect -10719 75540 -10645 75574
rect -10719 75506 -10699 75540
rect -10665 75506 -10645 75540
rect -10719 75472 -10645 75506
rect -10719 75438 -10699 75472
rect -10665 75438 -10645 75472
rect -10719 75404 -10645 75438
rect -10719 75370 -10699 75404
rect -10665 75370 -10645 75404
rect -10719 75336 -10645 75370
rect -10719 75302 -10699 75336
rect -10665 75302 -10645 75336
rect -10719 75268 -10645 75302
rect -10719 75234 -10699 75268
rect -10665 75234 -10645 75268
rect -10719 75200 -10645 75234
rect -10719 75166 -10699 75200
rect -10665 75166 -10645 75200
rect -10719 75132 -10645 75166
rect -10719 75098 -10699 75132
rect -10665 75098 -10645 75132
rect -10719 75064 -10645 75098
rect -10719 75030 -10699 75064
rect -10665 75030 -10645 75064
rect -10719 74996 -10645 75030
rect -10719 74962 -10699 74996
rect -10665 74962 -10645 74996
rect -10719 74928 -10645 74962
rect -10719 74894 -10699 74928
rect -10665 74894 -10645 74928
rect -10719 74860 -10645 74894
rect -10719 74826 -10699 74860
rect -10665 74826 -10645 74860
rect -10719 74792 -10645 74826
rect -10719 74758 -10699 74792
rect -10665 74758 -10645 74792
rect -10719 74724 -10645 74758
rect -10719 74690 -10699 74724
rect -10665 74690 -10645 74724
rect -10719 74656 -10645 74690
rect -10719 74622 -10699 74656
rect -10665 74622 -10645 74656
rect -10719 74588 -10645 74622
rect -10719 74554 -10699 74588
rect -10665 74554 -10645 74588
rect -10719 74520 -10645 74554
rect -10719 74486 -10699 74520
rect -10665 74486 -10645 74520
rect -10719 74452 -10645 74486
rect -10719 74418 -10699 74452
rect -10665 74418 -10645 74452
rect -10719 74384 -10645 74418
rect -10719 74350 -10699 74384
rect -10665 74350 -10645 74384
rect -10719 74316 -10645 74350
rect -10719 74282 -10699 74316
rect -10665 74282 -10645 74316
rect -10719 74248 -10645 74282
rect -10719 74214 -10699 74248
rect -10665 74214 -10645 74248
rect -10719 74180 -10645 74214
rect -10719 74146 -10699 74180
rect -10665 74146 -10645 74180
rect -10719 74112 -10645 74146
rect -10719 74078 -10699 74112
rect -10665 74078 -10645 74112
rect -10719 74044 -10645 74078
rect -10719 74010 -10699 74044
rect -10665 74010 -10645 74044
rect -10719 73976 -10645 74010
rect -10719 73942 -10699 73976
rect -10665 73942 -10645 73976
rect -10719 73908 -10645 73942
rect -10719 73874 -10699 73908
rect -10665 73874 -10645 73908
rect -10719 73840 -10645 73874
rect -10719 73806 -10699 73840
rect -10665 73806 -10645 73840
rect -10719 73772 -10645 73806
rect -10719 73738 -10699 73772
rect -10665 73738 -10645 73772
rect -10719 73704 -10645 73738
rect -10719 73670 -10699 73704
rect -10665 73670 -10645 73704
rect -10719 73636 -10645 73670
rect -10719 73602 -10699 73636
rect -10665 73602 -10645 73636
rect -10719 73568 -10645 73602
rect -10719 73534 -10699 73568
rect -10665 73534 -10645 73568
rect -10719 73500 -10645 73534
rect -10719 73466 -10699 73500
rect -10665 73466 -10645 73500
rect -10719 73432 -10645 73466
rect -10719 73398 -10699 73432
rect -10665 73398 -10645 73432
rect -10719 73364 -10645 73398
rect -10719 73330 -10699 73364
rect -10665 73330 -10645 73364
rect -10719 73296 -10645 73330
rect -10719 73262 -10699 73296
rect -10665 73262 -10645 73296
rect -10719 73228 -10645 73262
rect -10719 73194 -10699 73228
rect -10665 73194 -10645 73228
rect -10719 73160 -10645 73194
rect -10719 73126 -10699 73160
rect -10665 73126 -10645 73160
rect -10719 73092 -10645 73126
rect -10719 73058 -10699 73092
rect -10665 73058 -10645 73092
rect -10719 73024 -10645 73058
rect -10719 72990 -10699 73024
rect -10665 72990 -10645 73024
rect -10719 72956 -10645 72990
rect -10719 72922 -10699 72956
rect -10665 72922 -10645 72956
rect -10719 72888 -10645 72922
rect -10719 72854 -10699 72888
rect -10665 72854 -10645 72888
rect -10719 72820 -10645 72854
rect -10719 72786 -10699 72820
rect -10665 72786 -10645 72820
rect -10719 72752 -10645 72786
rect -10719 72718 -10699 72752
rect -10665 72718 -10645 72752
rect -10719 72684 -10645 72718
rect -10719 72650 -10699 72684
rect -10665 72650 -10645 72684
rect -10719 72616 -10645 72650
rect -10719 72582 -10699 72616
rect -10665 72582 -10645 72616
rect -10719 72548 -10645 72582
rect -10719 72514 -10699 72548
rect -10665 72514 -10645 72548
rect -10719 72480 -10645 72514
rect -10719 72446 -10699 72480
rect -10665 72446 -10645 72480
rect -10719 72412 -10645 72446
rect -10719 72378 -10699 72412
rect -10665 72378 -10645 72412
rect -10719 72344 -10645 72378
rect -10719 72310 -10699 72344
rect -10665 72310 -10645 72344
rect -10719 72276 -10645 72310
rect -10719 72242 -10699 72276
rect -10665 72242 -10645 72276
rect -10719 72208 -10645 72242
rect -10719 72174 -10699 72208
rect -10665 72174 -10645 72208
rect -10719 72140 -10645 72174
rect -10719 72106 -10699 72140
rect -10665 72106 -10645 72140
rect -10719 72072 -10645 72106
rect -10719 72038 -10699 72072
rect -10665 72038 -10645 72072
rect -10719 72004 -10645 72038
rect -10719 71970 -10699 72004
rect -10665 71970 -10645 72004
rect -10719 71936 -10645 71970
rect -10719 71902 -10699 71936
rect -10665 71902 -10645 71936
rect -10719 71868 -10645 71902
rect -10719 71834 -10699 71868
rect -10665 71834 -10645 71868
rect -10719 71800 -10645 71834
rect -10719 71766 -10699 71800
rect -10665 71766 -10645 71800
rect -10719 71732 -10645 71766
rect -10719 71698 -10699 71732
rect -10665 71698 -10645 71732
rect -10719 71664 -10645 71698
rect -10719 71630 -10699 71664
rect -10665 71630 -10645 71664
rect -10719 71596 -10645 71630
rect -10719 71562 -10699 71596
rect -10665 71562 -10645 71596
rect -10719 71528 -10645 71562
rect -10719 71494 -10699 71528
rect -10665 71494 -10645 71528
rect -10719 71460 -10645 71494
rect -10719 71426 -10699 71460
rect -10665 71426 -10645 71460
rect -10719 71392 -10645 71426
rect -10719 71358 -10699 71392
rect -10665 71358 -10645 71392
rect -10719 71324 -10645 71358
rect -10719 71290 -10699 71324
rect -10665 71290 -10645 71324
rect -10719 71256 -10645 71290
rect -10719 71222 -10699 71256
rect -10665 71222 -10645 71256
rect -10719 71188 -10645 71222
rect -10719 71154 -10699 71188
rect -10665 71154 -10645 71188
rect -10719 71120 -10645 71154
rect -10719 71086 -10699 71120
rect -10665 71086 -10645 71120
rect -10719 71052 -10645 71086
rect -10719 71018 -10699 71052
rect -10665 71018 -10645 71052
rect -10719 70984 -10645 71018
rect -10719 70950 -10699 70984
rect -10665 70950 -10645 70984
rect -10719 70916 -10645 70950
rect -10719 70882 -10699 70916
rect -10665 70882 -10645 70916
rect -10719 70848 -10645 70882
rect -10719 70814 -10699 70848
rect -10665 70814 -10645 70848
rect -10719 70780 -10645 70814
rect -10719 70746 -10699 70780
rect -10665 70746 -10645 70780
rect -10719 70712 -10645 70746
rect -10719 70678 -10699 70712
rect -10665 70678 -10645 70712
rect -10719 70644 -10645 70678
rect -10719 70610 -10699 70644
rect -10665 70610 -10645 70644
rect -10719 70576 -10645 70610
rect -10719 70542 -10699 70576
rect -10665 70542 -10645 70576
rect -10719 70508 -10645 70542
rect -10719 70474 -10699 70508
rect -10665 70474 -10645 70508
rect -10719 70440 -10645 70474
rect -10719 70406 -10699 70440
rect -10665 70406 -10645 70440
rect -10719 70372 -10645 70406
rect -10719 70338 -10699 70372
rect -10665 70338 -10645 70372
rect -10719 70304 -10645 70338
rect -10719 70270 -10699 70304
rect -10665 70270 -10645 70304
rect -10719 70236 -10645 70270
rect -10719 70202 -10699 70236
rect -10665 70202 -10645 70236
rect -10719 70168 -10645 70202
rect -10719 70134 -10699 70168
rect -10665 70134 -10645 70168
rect -10719 70100 -10645 70134
rect -10719 70066 -10699 70100
rect -10665 70066 -10645 70100
rect -10719 70032 -10645 70066
rect -10719 69998 -10699 70032
rect -10665 69998 -10645 70032
rect -10719 69964 -10645 69998
rect -10719 69930 -10699 69964
rect -10665 69930 -10645 69964
rect -10719 69896 -10645 69930
rect -10719 69862 -10699 69896
rect -10665 69862 -10645 69896
rect -10719 69828 -10645 69862
rect -10719 69794 -10699 69828
rect -10665 69794 -10645 69828
rect -10719 69760 -10645 69794
rect -10719 69726 -10699 69760
rect -10665 69726 -10645 69760
rect -10719 69692 -10645 69726
rect -10719 69658 -10699 69692
rect -10665 69658 -10645 69692
rect -10719 69624 -10645 69658
rect -10719 69590 -10699 69624
rect -10665 69590 -10645 69624
rect -10719 69556 -10645 69590
rect -10719 69522 -10699 69556
rect -10665 69522 -10645 69556
rect -10719 69488 -10645 69522
rect -10719 69454 -10699 69488
rect -10665 69454 -10645 69488
rect -10719 69420 -10645 69454
rect -10719 69386 -10699 69420
rect -10665 69386 -10645 69420
rect -10719 69352 -10645 69386
rect -10719 69318 -10699 69352
rect -10665 69318 -10645 69352
rect -10719 69284 -10645 69318
rect -10719 69250 -10699 69284
rect -10665 69250 -10645 69284
rect -10719 69216 -10645 69250
rect -10719 69182 -10699 69216
rect -10665 69182 -10645 69216
rect -10719 69148 -10645 69182
rect -10719 69114 -10699 69148
rect -10665 69114 -10645 69148
rect -10719 69080 -10645 69114
rect -10719 69046 -10699 69080
rect -10665 69046 -10645 69080
rect -10719 69012 -10645 69046
rect -10719 68978 -10699 69012
rect -10665 68978 -10645 69012
rect -10719 68944 -10645 68978
rect -10719 68910 -10699 68944
rect -10665 68910 -10645 68944
rect -10719 68876 -10645 68910
rect -10719 68842 -10699 68876
rect -10665 68842 -10645 68876
rect -10719 68808 -10645 68842
rect -10719 68774 -10699 68808
rect -10665 68774 -10645 68808
rect -10719 68740 -10645 68774
rect -10719 68706 -10699 68740
rect -10665 68706 -10645 68740
rect -10719 68672 -10645 68706
rect -10719 68638 -10699 68672
rect -10665 68638 -10645 68672
rect -10719 68604 -10645 68638
rect -10719 68570 -10699 68604
rect -10665 68570 -10645 68604
rect -10719 68536 -10645 68570
rect -10719 68502 -10699 68536
rect -10665 68502 -10645 68536
rect -10719 68468 -10645 68502
rect -10719 68434 -10699 68468
rect -10665 68434 -10645 68468
rect -10719 68400 -10645 68434
rect -10719 68366 -10699 68400
rect -10665 68366 -10645 68400
rect -10719 68332 -10645 68366
rect -10719 68298 -10699 68332
rect -10665 68298 -10645 68332
rect -10719 68264 -10645 68298
rect -10719 68230 -10699 68264
rect -10665 68230 -10645 68264
rect -10719 68196 -10645 68230
rect -10719 68162 -10699 68196
rect -10665 68162 -10645 68196
rect -10719 68128 -10645 68162
rect -10719 68094 -10699 68128
rect -10665 68094 -10645 68128
rect -10719 68060 -10645 68094
rect -10719 68026 -10699 68060
rect -10665 68026 -10645 68060
rect -10719 67992 -10645 68026
rect -10719 67958 -10699 67992
rect -10665 67958 -10645 67992
rect -10719 67924 -10645 67958
rect -10719 67890 -10699 67924
rect -10665 67890 -10645 67924
rect -10719 67856 -10645 67890
rect -10719 67822 -10699 67856
rect -10665 67822 -10645 67856
rect -10719 67788 -10645 67822
rect -10719 67754 -10699 67788
rect -10665 67754 -10645 67788
rect -10719 67720 -10645 67754
rect -10719 67686 -10699 67720
rect -10665 67686 -10645 67720
rect -10719 67652 -10645 67686
rect -10719 67618 -10699 67652
rect -10665 67618 -10645 67652
rect -10719 67584 -10645 67618
rect -10719 67550 -10699 67584
rect -10665 67550 -10645 67584
rect -10719 67516 -10645 67550
rect -10719 67482 -10699 67516
rect -10665 67482 -10645 67516
rect -10719 67448 -10645 67482
rect -10719 67414 -10699 67448
rect -10665 67414 -10645 67448
rect -10719 67380 -10645 67414
rect -10719 67346 -10699 67380
rect -10665 67346 -10645 67380
rect -10719 67312 -10645 67346
rect -10719 67278 -10699 67312
rect -10665 67278 -10645 67312
rect -10719 67244 -10645 67278
rect -10719 67210 -10699 67244
rect -10665 67210 -10645 67244
rect -10719 67176 -10645 67210
rect -10719 67142 -10699 67176
rect -10665 67142 -10645 67176
rect -10719 67108 -10645 67142
rect -10719 67074 -10699 67108
rect -10665 67074 -10645 67108
rect -10719 67040 -10645 67074
rect -10719 67006 -10699 67040
rect -10665 67006 -10645 67040
rect -10719 66972 -10645 67006
rect -10719 66938 -10699 66972
rect -10665 66938 -10645 66972
rect -10719 66904 -10645 66938
rect -10719 66870 -10699 66904
rect -10665 66870 -10645 66904
rect -10719 66836 -10645 66870
rect -10719 66802 -10699 66836
rect -10665 66802 -10645 66836
rect -10719 66768 -10645 66802
rect -10719 66734 -10699 66768
rect -10665 66734 -10645 66768
rect -10719 66700 -10645 66734
rect -10719 66666 -10699 66700
rect -10665 66666 -10645 66700
rect -10719 66632 -10645 66666
rect -10719 66598 -10699 66632
rect -10665 66598 -10645 66632
rect -10719 66564 -10645 66598
rect -10719 66530 -10699 66564
rect -10665 66530 -10645 66564
rect -10719 66496 -10645 66530
rect -10719 66462 -10699 66496
rect -10665 66462 -10645 66496
rect -10719 66428 -10645 66462
rect -10719 66394 -10699 66428
rect -10665 66394 -10645 66428
rect -10719 66360 -10645 66394
rect -10719 66326 -10699 66360
rect -10665 66326 -10645 66360
rect -10719 66292 -10645 66326
rect -10719 66258 -10699 66292
rect -10665 66258 -10645 66292
rect -10719 66224 -10645 66258
rect -10719 66190 -10699 66224
rect -10665 66190 -10645 66224
rect -10719 66156 -10645 66190
rect -10719 66122 -10699 66156
rect -10665 66122 -10645 66156
rect -10719 66088 -10645 66122
rect -10719 66054 -10699 66088
rect -10665 66054 -10645 66088
rect -10719 66020 -10645 66054
rect -10719 65986 -10699 66020
rect -10665 65986 -10645 66020
rect -10719 65952 -10645 65986
rect -10719 65918 -10699 65952
rect -10665 65918 -10645 65952
rect -10719 65884 -10645 65918
rect -10719 65850 -10699 65884
rect -10665 65850 -10645 65884
rect -10719 65816 -10645 65850
rect -10719 65782 -10699 65816
rect -10665 65782 -10645 65816
rect -10719 65748 -10645 65782
rect -10719 65714 -10699 65748
rect -10665 65714 -10645 65748
rect -10719 65680 -10645 65714
rect -10719 65646 -10699 65680
rect -10665 65646 -10645 65680
rect -10719 65612 -10645 65646
rect -10719 65578 -10699 65612
rect -10665 65578 -10645 65612
rect -10719 65544 -10645 65578
rect -10719 65510 -10699 65544
rect -10665 65510 -10645 65544
rect -10719 65476 -10645 65510
rect -10719 65442 -10699 65476
rect -10665 65442 -10645 65476
rect -10719 65408 -10645 65442
rect -10719 65374 -10699 65408
rect -10665 65374 -10645 65408
rect -10719 65340 -10645 65374
rect -10719 65306 -10699 65340
rect -10665 65306 -10645 65340
rect -10719 65272 -10645 65306
rect -10719 65238 -10699 65272
rect -10665 65238 -10645 65272
rect -10719 65204 -10645 65238
rect -10719 65170 -10699 65204
rect -10665 65170 -10645 65204
rect -10719 65136 -10645 65170
rect -10719 65102 -10699 65136
rect -10665 65102 -10645 65136
rect -10719 65068 -10645 65102
rect -10719 65034 -10699 65068
rect -10665 65034 -10645 65068
rect -10719 65000 -10645 65034
rect -10719 64966 -10699 65000
rect -10665 64966 -10645 65000
rect -10719 64932 -10645 64966
rect -10719 64898 -10699 64932
rect -10665 64898 -10645 64932
rect -10719 64864 -10645 64898
rect -10719 64830 -10699 64864
rect -10665 64830 -10645 64864
rect -10719 64796 -10645 64830
rect -10719 64762 -10699 64796
rect -10665 64762 -10645 64796
rect -10719 64728 -10645 64762
rect -10719 64694 -10699 64728
rect -10665 64694 -10645 64728
rect -10719 64660 -10645 64694
rect -10719 64626 -10699 64660
rect -10665 64626 -10645 64660
rect -10719 64592 -10645 64626
rect -10719 64558 -10699 64592
rect -10665 64558 -10645 64592
rect -10719 64524 -10645 64558
rect -10719 64490 -10699 64524
rect -10665 64490 -10645 64524
rect -10719 64456 -10645 64490
rect -10719 64422 -10699 64456
rect -10665 64422 -10645 64456
rect -10719 64388 -10645 64422
rect -10719 64354 -10699 64388
rect -10665 64354 -10645 64388
rect -10719 64320 -10645 64354
rect -10719 64286 -10699 64320
rect -10665 64286 -10645 64320
rect -10719 64252 -10645 64286
rect -10719 64218 -10699 64252
rect -10665 64218 -10645 64252
rect -10719 64184 -10645 64218
rect -10719 64150 -10699 64184
rect -10665 64150 -10645 64184
rect -10719 64140 -10645 64150
rect -3738 76056 -3664 76090
rect -3738 76022 -3718 76056
rect -3684 76022 -3664 76056
rect -3738 75988 -3664 76022
rect -3738 75954 -3718 75988
rect -3684 75954 -3664 75988
rect -3738 75920 -3664 75954
rect -3738 75886 -3718 75920
rect -3684 75886 -3664 75920
rect -3738 75852 -3664 75886
rect -3738 75818 -3718 75852
rect -3684 75818 -3664 75852
rect -3738 75784 -3664 75818
rect -3738 75750 -3718 75784
rect -3684 75750 -3664 75784
rect -3738 75716 -3664 75750
rect -3738 75682 -3718 75716
rect -3684 75682 -3664 75716
rect -3738 75648 -3664 75682
rect -3738 75614 -3718 75648
rect -3684 75614 -3664 75648
rect -3738 75580 -3664 75614
rect -3738 75546 -3718 75580
rect -3684 75546 -3664 75580
rect -3738 75512 -3664 75546
rect -3738 75478 -3718 75512
rect -3684 75478 -3664 75512
rect -3738 75444 -3664 75478
rect -3738 75410 -3718 75444
rect -3684 75410 -3664 75444
rect -3738 75376 -3664 75410
rect -3738 75342 -3718 75376
rect -3684 75342 -3664 75376
rect -3738 75308 -3664 75342
rect -3738 75274 -3718 75308
rect -3684 75274 -3664 75308
rect -3738 75240 -3664 75274
rect -3738 75206 -3718 75240
rect -3684 75206 -3664 75240
rect -3738 75172 -3664 75206
rect -3738 75138 -3718 75172
rect -3684 75138 -3664 75172
rect -3738 75104 -3664 75138
rect -3738 75070 -3718 75104
rect -3684 75070 -3664 75104
rect -3738 75036 -3664 75070
rect -3738 75002 -3718 75036
rect -3684 75002 -3664 75036
rect -3738 74968 -3664 75002
rect -3738 74934 -3718 74968
rect -3684 74934 -3664 74968
rect -3738 74900 -3664 74934
rect -3738 74866 -3718 74900
rect -3684 74866 -3664 74900
rect -3738 74832 -3664 74866
rect -3738 74798 -3718 74832
rect -3684 74798 -3664 74832
rect -3738 74764 -3664 74798
rect -3738 74730 -3718 74764
rect -3684 74730 -3664 74764
rect -3738 74696 -3664 74730
rect -3738 74662 -3718 74696
rect -3684 74662 -3664 74696
rect -3738 74628 -3664 74662
rect -3738 74594 -3718 74628
rect -3684 74594 -3664 74628
rect -3738 74560 -3664 74594
rect -3738 74526 -3718 74560
rect -3684 74526 -3664 74560
rect -3738 74492 -3664 74526
rect -3738 74458 -3718 74492
rect -3684 74458 -3664 74492
rect -3738 74424 -3664 74458
rect -3738 74390 -3718 74424
rect -3684 74390 -3664 74424
rect -3738 74356 -3664 74390
rect -3738 74322 -3718 74356
rect -3684 74322 -3664 74356
rect -3738 74288 -3664 74322
rect -3738 74254 -3718 74288
rect -3684 74254 -3664 74288
rect -3738 74220 -3664 74254
rect -3738 74186 -3718 74220
rect -3684 74186 -3664 74220
rect -3738 74152 -3664 74186
rect -3738 74118 -3718 74152
rect -3684 74118 -3664 74152
rect -3738 74084 -3664 74118
rect -3738 74050 -3718 74084
rect -3684 74050 -3664 74084
rect -3738 74016 -3664 74050
rect -3738 73982 -3718 74016
rect -3684 73982 -3664 74016
rect -3738 73948 -3664 73982
rect -3738 73914 -3718 73948
rect -3684 73914 -3664 73948
rect -3738 73880 -3664 73914
rect -3738 73846 -3718 73880
rect -3684 73846 -3664 73880
rect -3738 73812 -3664 73846
rect -3738 73778 -3718 73812
rect -3684 73778 -3664 73812
rect -3738 73744 -3664 73778
rect -3738 73710 -3718 73744
rect -3684 73710 -3664 73744
rect -3738 73676 -3664 73710
rect -3738 73642 -3718 73676
rect -3684 73642 -3664 73676
rect -3738 73608 -3664 73642
rect -3738 73574 -3718 73608
rect -3684 73574 -3664 73608
rect -3738 73540 -3664 73574
rect -3738 73506 -3718 73540
rect -3684 73506 -3664 73540
rect -3738 73472 -3664 73506
rect -3738 73438 -3718 73472
rect -3684 73438 -3664 73472
rect -3738 73404 -3664 73438
rect -3738 73370 -3718 73404
rect -3684 73370 -3664 73404
rect -3738 73336 -3664 73370
rect -3738 73302 -3718 73336
rect -3684 73302 -3664 73336
rect -3738 73268 -3664 73302
rect -3738 73234 -3718 73268
rect -3684 73234 -3664 73268
rect -3738 73200 -3664 73234
rect -3738 73166 -3718 73200
rect -3684 73166 -3664 73200
rect -3738 73132 -3664 73166
rect -3738 73098 -3718 73132
rect -3684 73098 -3664 73132
rect -3738 73064 -3664 73098
rect -3738 73030 -3718 73064
rect -3684 73030 -3664 73064
rect -3738 72996 -3664 73030
rect -3738 72962 -3718 72996
rect -3684 72962 -3664 72996
rect -3738 72928 -3664 72962
rect -3738 72894 -3718 72928
rect -3684 72894 -3664 72928
rect -3738 72860 -3664 72894
rect -3738 72826 -3718 72860
rect -3684 72826 -3664 72860
rect -3738 72792 -3664 72826
rect -3738 72758 -3718 72792
rect -3684 72758 -3664 72792
rect -3738 72724 -3664 72758
rect -3738 72690 -3718 72724
rect -3684 72690 -3664 72724
rect -3738 72656 -3664 72690
rect -3738 72622 -3718 72656
rect -3684 72622 -3664 72656
rect -3738 72588 -3664 72622
rect -3738 72554 -3718 72588
rect -3684 72554 -3664 72588
rect -3738 72520 -3664 72554
rect -3738 72486 -3718 72520
rect -3684 72486 -3664 72520
rect -3738 72452 -3664 72486
rect -3738 72418 -3718 72452
rect -3684 72418 -3664 72452
rect -3738 72384 -3664 72418
rect -3738 72350 -3718 72384
rect -3684 72350 -3664 72384
rect -3738 72316 -3664 72350
rect -3738 72282 -3718 72316
rect -3684 72282 -3664 72316
rect -3738 72248 -3664 72282
rect -3738 72214 -3718 72248
rect -3684 72214 -3664 72248
rect -3738 72180 -3664 72214
rect -3738 72146 -3718 72180
rect -3684 72146 -3664 72180
rect -3738 72112 -3664 72146
rect -3738 72078 -3718 72112
rect -3684 72078 -3664 72112
rect -3738 72044 -3664 72078
rect -3738 72010 -3718 72044
rect -3684 72010 -3664 72044
rect -3738 71976 -3664 72010
rect -3738 71942 -3718 71976
rect -3684 71942 -3664 71976
rect -3738 71908 -3664 71942
rect -3738 71874 -3718 71908
rect -3684 71874 -3664 71908
rect -3738 71840 -3664 71874
rect -3738 71806 -3718 71840
rect -3684 71806 -3664 71840
rect -3738 71772 -3664 71806
rect -3738 71738 -3718 71772
rect -3684 71738 -3664 71772
rect -3738 71704 -3664 71738
rect -3738 71670 -3718 71704
rect -3684 71670 -3664 71704
rect -3738 71636 -3664 71670
rect -3738 71602 -3718 71636
rect -3684 71602 -3664 71636
rect -3738 71568 -3664 71602
rect -3738 71534 -3718 71568
rect -3684 71534 -3664 71568
rect -3738 71500 -3664 71534
rect -3738 71466 -3718 71500
rect -3684 71466 -3664 71500
rect -3738 71432 -3664 71466
rect -3738 71398 -3718 71432
rect -3684 71398 -3664 71432
rect -3738 71364 -3664 71398
rect -3738 71330 -3718 71364
rect -3684 71330 -3664 71364
rect -3738 71296 -3664 71330
rect -3738 71262 -3718 71296
rect -3684 71262 -3664 71296
rect -3738 71228 -3664 71262
rect -3738 71194 -3718 71228
rect -3684 71194 -3664 71228
rect -3738 71160 -3664 71194
rect -3738 71126 -3718 71160
rect -3684 71126 -3664 71160
rect -3738 71092 -3664 71126
rect -3738 71058 -3718 71092
rect -3684 71058 -3664 71092
rect -3738 71024 -3664 71058
rect -3738 70990 -3718 71024
rect -3684 70990 -3664 71024
rect -3738 70956 -3664 70990
rect -3738 70922 -3718 70956
rect -3684 70922 -3664 70956
rect -3738 70888 -3664 70922
rect -3738 70854 -3718 70888
rect -3684 70854 -3664 70888
rect -3738 70820 -3664 70854
rect -3738 70786 -3718 70820
rect -3684 70786 -3664 70820
rect -3738 70752 -3664 70786
rect -3738 70718 -3718 70752
rect -3684 70718 -3664 70752
rect -3738 70684 -3664 70718
rect -3738 70650 -3718 70684
rect -3684 70650 -3664 70684
rect -3738 70616 -3664 70650
rect -3738 70582 -3718 70616
rect -3684 70582 -3664 70616
rect -3738 70548 -3664 70582
rect -3738 70514 -3718 70548
rect -3684 70514 -3664 70548
rect -3738 70480 -3664 70514
rect -3738 70446 -3718 70480
rect -3684 70446 -3664 70480
rect -3738 70412 -3664 70446
rect -3738 70378 -3718 70412
rect -3684 70378 -3664 70412
rect -3738 70344 -3664 70378
rect -3738 70310 -3718 70344
rect -3684 70310 -3664 70344
rect -3738 70276 -3664 70310
rect -3738 70242 -3718 70276
rect -3684 70242 -3664 70276
rect -3738 70208 -3664 70242
rect -3738 70174 -3718 70208
rect -3684 70174 -3664 70208
rect -3738 70140 -3664 70174
rect -3738 70106 -3718 70140
rect -3684 70106 -3664 70140
rect -3738 70072 -3664 70106
rect -3738 70038 -3718 70072
rect -3684 70038 -3664 70072
rect -3738 70004 -3664 70038
rect -3738 69970 -3718 70004
rect -3684 69970 -3664 70004
rect -3738 69936 -3664 69970
rect -3738 69902 -3718 69936
rect -3684 69902 -3664 69936
rect -3738 69868 -3664 69902
rect -3738 69834 -3718 69868
rect -3684 69834 -3664 69868
rect -3738 69800 -3664 69834
rect -3738 69766 -3718 69800
rect -3684 69766 -3664 69800
rect -3738 69732 -3664 69766
rect -3738 69698 -3718 69732
rect -3684 69698 -3664 69732
rect -3738 69664 -3664 69698
rect -3738 69630 -3718 69664
rect -3684 69630 -3664 69664
rect -3738 69596 -3664 69630
rect -3738 69562 -3718 69596
rect -3684 69562 -3664 69596
rect -3738 69528 -3664 69562
rect -3738 69494 -3718 69528
rect -3684 69494 -3664 69528
rect -3738 69460 -3664 69494
rect -3738 69426 -3718 69460
rect -3684 69426 -3664 69460
rect -3738 69392 -3664 69426
rect -3738 69358 -3718 69392
rect -3684 69358 -3664 69392
rect -3738 69324 -3664 69358
rect -3738 69290 -3718 69324
rect -3684 69290 -3664 69324
rect -3738 69256 -3664 69290
rect -3738 69222 -3718 69256
rect -3684 69222 -3664 69256
rect -3738 69188 -3664 69222
rect -3738 69154 -3718 69188
rect -3684 69154 -3664 69188
rect -3738 69120 -3664 69154
rect -3738 69086 -3718 69120
rect -3684 69086 -3664 69120
rect -3738 69052 -3664 69086
rect -3738 69018 -3718 69052
rect -3684 69018 -3664 69052
rect -3738 68984 -3664 69018
rect -3738 68950 -3718 68984
rect -3684 68950 -3664 68984
rect -3738 68916 -3664 68950
rect -3738 68882 -3718 68916
rect -3684 68882 -3664 68916
rect -3738 68848 -3664 68882
rect -3738 68814 -3718 68848
rect -3684 68814 -3664 68848
rect -3738 68780 -3664 68814
rect -3738 68746 -3718 68780
rect -3684 68746 -3664 68780
rect -3738 68712 -3664 68746
rect -3738 68678 -3718 68712
rect -3684 68678 -3664 68712
rect -3738 68644 -3664 68678
rect -3738 68610 -3718 68644
rect -3684 68610 -3664 68644
rect -3738 68576 -3664 68610
rect -3738 68542 -3718 68576
rect -3684 68542 -3664 68576
rect -3738 68508 -3664 68542
rect -3738 68474 -3718 68508
rect -3684 68474 -3664 68508
rect -3738 68440 -3664 68474
rect -3738 68406 -3718 68440
rect -3684 68406 -3664 68440
rect -3738 68372 -3664 68406
rect -3738 68338 -3718 68372
rect -3684 68338 -3664 68372
rect -3738 68304 -3664 68338
rect -3738 68270 -3718 68304
rect -3684 68270 -3664 68304
rect -3738 68236 -3664 68270
rect -3738 68202 -3718 68236
rect -3684 68202 -3664 68236
rect -3738 68168 -3664 68202
rect -3738 68134 -3718 68168
rect -3684 68134 -3664 68168
rect -3738 68100 -3664 68134
rect -3738 68066 -3718 68100
rect -3684 68066 -3664 68100
rect -3738 68032 -3664 68066
rect -3738 67998 -3718 68032
rect -3684 67998 -3664 68032
rect -3738 67964 -3664 67998
rect -3738 67930 -3718 67964
rect -3684 67930 -3664 67964
rect -3738 67896 -3664 67930
rect -3738 67862 -3718 67896
rect -3684 67862 -3664 67896
rect -3738 67828 -3664 67862
rect -3738 67794 -3718 67828
rect -3684 67794 -3664 67828
rect -3738 67760 -3664 67794
rect -3738 67726 -3718 67760
rect -3684 67726 -3664 67760
rect -3738 67692 -3664 67726
rect -3738 67658 -3718 67692
rect -3684 67658 -3664 67692
rect -3738 67624 -3664 67658
rect -3738 67590 -3718 67624
rect -3684 67590 -3664 67624
rect -3738 67556 -3664 67590
rect -3738 67522 -3718 67556
rect -3684 67522 -3664 67556
rect -3738 67488 -3664 67522
rect -3738 67454 -3718 67488
rect -3684 67454 -3664 67488
rect -3738 67420 -3664 67454
rect -3738 67386 -3718 67420
rect -3684 67386 -3664 67420
rect -3738 67352 -3664 67386
rect -3738 67318 -3718 67352
rect -3684 67318 -3664 67352
rect -3738 67284 -3664 67318
rect -3738 67250 -3718 67284
rect -3684 67250 -3664 67284
rect -3738 67216 -3664 67250
rect -3738 67182 -3718 67216
rect -3684 67182 -3664 67216
rect -3738 67148 -3664 67182
rect -3738 67114 -3718 67148
rect -3684 67114 -3664 67148
rect -3738 67080 -3664 67114
rect -3738 67046 -3718 67080
rect -3684 67046 -3664 67080
rect -3738 67012 -3664 67046
rect -3738 66978 -3718 67012
rect -3684 66978 -3664 67012
rect -3738 66944 -3664 66978
rect -3738 66910 -3718 66944
rect -3684 66910 -3664 66944
rect -3738 66876 -3664 66910
rect -3738 66842 -3718 66876
rect -3684 66842 -3664 66876
rect -3738 66808 -3664 66842
rect -3738 66774 -3718 66808
rect -3684 66774 -3664 66808
rect -3738 66740 -3664 66774
rect -3738 66706 -3718 66740
rect -3684 66706 -3664 66740
rect -3738 66672 -3664 66706
rect -3738 66638 -3718 66672
rect -3684 66638 -3664 66672
rect -3738 66604 -3664 66638
rect -3738 66570 -3718 66604
rect -3684 66570 -3664 66604
rect -3738 66536 -3664 66570
rect -3738 66502 -3718 66536
rect -3684 66502 -3664 66536
rect -3738 66468 -3664 66502
rect -3738 66434 -3718 66468
rect -3684 66434 -3664 66468
rect -3738 66400 -3664 66434
rect -3738 66366 -3718 66400
rect -3684 66366 -3664 66400
rect -3738 66332 -3664 66366
rect -3738 66298 -3718 66332
rect -3684 66298 -3664 66332
rect -3738 66264 -3664 66298
rect -3738 66230 -3718 66264
rect -3684 66230 -3664 66264
rect -3738 66196 -3664 66230
rect -3738 66162 -3718 66196
rect -3684 66162 -3664 66196
rect -3738 66128 -3664 66162
rect -3738 66094 -3718 66128
rect -3684 66094 -3664 66128
rect -3738 66060 -3664 66094
rect -3738 66026 -3718 66060
rect -3684 66026 -3664 66060
rect -3738 65992 -3664 66026
rect -3738 65958 -3718 65992
rect -3684 65958 -3664 65992
rect -3738 65924 -3664 65958
rect -3738 65890 -3718 65924
rect -3684 65890 -3664 65924
rect -3738 65856 -3664 65890
rect -3738 65822 -3718 65856
rect -3684 65822 -3664 65856
rect -3738 65788 -3664 65822
rect -3738 65754 -3718 65788
rect -3684 65754 -3664 65788
rect -3738 65720 -3664 65754
rect -3738 65686 -3718 65720
rect -3684 65686 -3664 65720
rect -3738 65652 -3664 65686
rect -3738 65618 -3718 65652
rect -3684 65618 -3664 65652
rect -3738 65584 -3664 65618
rect -3738 65550 -3718 65584
rect -3684 65550 -3664 65584
rect -3738 65516 -3664 65550
rect -3738 65482 -3718 65516
rect -3684 65482 -3664 65516
rect -3738 65448 -3664 65482
rect -3738 65414 -3718 65448
rect -3684 65414 -3664 65448
rect -3738 65380 -3664 65414
rect -3738 65346 -3718 65380
rect -3684 65346 -3664 65380
rect -3738 65312 -3664 65346
rect -3738 65278 -3718 65312
rect -3684 65278 -3664 65312
rect -3738 65244 -3664 65278
rect -3738 65210 -3718 65244
rect -3684 65210 -3664 65244
rect -3738 65176 -3664 65210
rect -3738 65142 -3718 65176
rect -3684 65142 -3664 65176
rect -3738 65108 -3664 65142
rect -3738 65074 -3718 65108
rect -3684 65074 -3664 65108
rect -3738 65040 -3664 65074
rect -3738 65006 -3718 65040
rect -3684 65006 -3664 65040
rect -3738 64972 -3664 65006
rect -3738 64938 -3718 64972
rect -3684 64938 -3664 64972
rect -3738 64904 -3664 64938
rect -3738 64870 -3718 64904
rect -3684 64870 -3664 64904
rect -3738 64836 -3664 64870
rect -3738 64802 -3718 64836
rect -3684 64802 -3664 64836
rect -3738 64768 -3664 64802
rect -3738 64734 -3718 64768
rect -3684 64734 -3664 64768
rect -3738 64700 -3664 64734
rect -3738 64666 -3718 64700
rect -3684 64666 -3664 64700
rect -3738 64632 -3664 64666
rect -3738 64598 -3718 64632
rect -3684 64598 -3664 64632
rect -3738 64564 -3664 64598
rect -3738 64530 -3718 64564
rect -3684 64530 -3664 64564
rect -3738 64496 -3664 64530
rect -3738 64462 -3718 64496
rect -3684 64462 -3664 64496
rect -3738 64428 -3664 64462
rect -3738 64394 -3718 64428
rect -3684 64394 -3664 64428
rect -3738 64360 -3664 64394
rect -3738 64326 -3718 64360
rect -3684 64326 -3664 64360
rect -3738 64292 -3664 64326
rect -3738 64258 -3718 64292
rect -3684 64258 -3664 64292
rect -3738 64224 -3664 64258
rect -3738 64190 -3718 64224
rect -3684 64190 -3664 64224
rect -3738 64156 -3664 64190
rect -10719 64120 -7153 64140
rect -10719 64086 -10624 64120
rect -10590 64086 -10556 64120
rect -10522 64086 -10488 64120
rect -10454 64086 -10420 64120
rect -10386 64086 -10352 64120
rect -10318 64086 -10284 64120
rect -10250 64086 -10216 64120
rect -10182 64086 -10148 64120
rect -10114 64086 -10080 64120
rect -10046 64086 -10012 64120
rect -9978 64086 -9944 64120
rect -9910 64086 -9876 64120
rect -9842 64086 -9808 64120
rect -9774 64086 -9740 64120
rect -9706 64086 -9672 64120
rect -9638 64086 -9604 64120
rect -9570 64086 -9536 64120
rect -9502 64086 -9468 64120
rect -9434 64086 -9400 64120
rect -9366 64086 -9332 64120
rect -9298 64086 -9264 64120
rect -9230 64086 -9196 64120
rect -9162 64086 -9128 64120
rect -9094 64086 -9060 64120
rect -9026 64086 -8992 64120
rect -8958 64086 -8924 64120
rect -8890 64086 -8856 64120
rect -8822 64086 -8788 64120
rect -8754 64086 -8720 64120
rect -8686 64086 -8652 64120
rect -8618 64086 -8584 64120
rect -8550 64086 -8516 64120
rect -8482 64086 -8448 64120
rect -8414 64086 -8380 64120
rect -8346 64086 -8312 64120
rect -8278 64086 -8244 64120
rect -8210 64086 -8176 64120
rect -8142 64086 -8108 64120
rect -8074 64086 -8040 64120
rect -8006 64086 -7972 64120
rect -7938 64086 -7904 64120
rect -7870 64086 -7836 64120
rect -7802 64086 -7768 64120
rect -7734 64086 -7700 64120
rect -7666 64086 -7632 64120
rect -7598 64086 -7564 64120
rect -7530 64086 -7496 64120
rect -7462 64086 -7428 64120
rect -7394 64086 -7360 64120
rect -7326 64086 -7292 64120
rect -7258 64086 -7153 64120
rect -10719 64066 -7153 64086
rect -7227 64059 -7153 64066
rect -7227 64025 -7207 64059
rect -7173 64025 -7153 64059
rect -7227 63991 -7153 64025
rect -7227 63957 -7207 63991
rect -7173 63957 -7153 63991
rect -7227 63923 -7153 63957
rect -7227 63889 -7207 63923
rect -7173 63889 -7153 63923
rect -7227 63855 -7153 63889
rect -7227 63821 -7207 63855
rect -7173 63821 -7153 63855
rect -7227 63787 -7153 63821
rect -7227 63753 -7207 63787
rect -7173 63753 -7153 63787
rect -7227 63719 -7153 63753
rect -7227 63685 -7207 63719
rect -7173 63685 -7153 63719
rect -7227 63651 -7153 63685
rect -7227 63617 -7207 63651
rect -7173 63617 -7153 63651
rect -7227 63583 -7153 63617
rect -7227 63549 -7207 63583
rect -7173 63549 -7153 63583
rect -7227 63515 -7153 63549
rect -7227 63481 -7207 63515
rect -7173 63481 -7153 63515
rect -7227 63447 -7153 63481
rect -7227 63413 -7207 63447
rect -7173 63413 -7153 63447
rect -7227 63379 -7153 63413
rect -7227 63345 -7207 63379
rect -7173 63345 -7153 63379
rect -7227 63311 -7153 63345
rect -7227 63277 -7207 63311
rect -7173 63277 -7153 63311
rect -7227 63243 -7153 63277
rect -7227 63209 -7207 63243
rect -7173 63209 -7153 63243
rect -7227 63175 -7153 63209
rect -7227 63141 -7207 63175
rect -7173 63141 -7153 63175
rect -7227 63107 -7153 63141
rect -7227 63073 -7207 63107
rect -7173 63073 -7153 63107
rect -7227 63039 -7153 63073
rect -7227 63005 -7207 63039
rect -7173 63005 -7153 63039
rect -7227 62971 -7153 63005
rect -7227 62937 -7207 62971
rect -7173 62937 -7153 62971
rect -7227 62903 -7153 62937
rect -7227 62869 -7207 62903
rect -7173 62869 -7153 62903
rect -7227 62835 -7153 62869
rect -7227 62801 -7207 62835
rect -7173 62801 -7153 62835
rect -7227 62767 -7153 62801
rect -7227 62733 -7207 62767
rect -7173 62733 -7153 62767
rect -7227 62699 -7153 62733
rect -7227 62665 -7207 62699
rect -7173 62665 -7153 62699
rect -7227 62631 -7153 62665
rect -7227 62597 -7207 62631
rect -7173 62597 -7153 62631
rect -7227 62563 -7153 62597
rect -7227 62529 -7207 62563
rect -7173 62529 -7153 62563
rect -7227 62495 -7153 62529
rect -7227 62461 -7207 62495
rect -7173 62461 -7153 62495
rect -7227 62427 -7153 62461
rect -7227 62393 -7207 62427
rect -7173 62393 -7153 62427
rect -7227 62359 -7153 62393
rect -7227 62325 -7207 62359
rect -7173 62325 -7153 62359
rect -7227 62291 -7153 62325
rect -7227 62257 -7207 62291
rect -7173 62257 -7153 62291
rect -7227 62223 -7153 62257
rect -7227 62189 -7207 62223
rect -7173 62189 -7153 62223
rect -7227 62155 -7153 62189
rect -7227 62121 -7207 62155
rect -7173 62121 -7153 62155
rect -7227 62087 -7153 62121
rect -7227 62053 -7207 62087
rect -7173 62053 -7153 62087
rect -7227 62019 -7153 62053
rect -7227 61985 -7207 62019
rect -7173 61985 -7153 62019
rect -7227 61951 -7153 61985
rect -7227 61917 -7207 61951
rect -7173 61917 -7153 61951
rect -7227 61883 -7153 61917
rect -7227 61849 -7207 61883
rect -7173 61849 -7153 61883
rect -7227 61815 -7153 61849
rect -7227 61781 -7207 61815
rect -7173 61781 -7153 61815
rect -7227 61747 -7153 61781
rect -7227 61713 -7207 61747
rect -7173 61713 -7153 61747
rect -7227 61679 -7153 61713
rect -7227 61645 -7207 61679
rect -7173 61645 -7153 61679
rect -7227 61611 -7153 61645
rect -7227 61577 -7207 61611
rect -7173 61577 -7153 61611
rect -7227 61543 -7153 61577
rect -7227 61509 -7207 61543
rect -7173 61509 -7153 61543
rect -7227 61475 -7153 61509
rect -7227 61441 -7207 61475
rect -7173 61441 -7153 61475
rect -7227 61407 -7153 61441
rect -7227 61373 -7207 61407
rect -7173 61373 -7153 61407
rect -7227 61339 -7153 61373
rect -7227 61305 -7207 61339
rect -7173 61305 -7153 61339
rect -7227 61271 -7153 61305
rect -7227 61237 -7207 61271
rect -7173 61237 -7153 61271
rect -7227 61203 -7153 61237
rect -7227 61169 -7207 61203
rect -7173 61169 -7153 61203
rect -7227 61135 -7153 61169
rect -7227 61101 -7207 61135
rect -7173 61101 -7153 61135
rect -7227 61067 -7153 61101
rect -7227 61033 -7207 61067
rect -7173 61033 -7153 61067
rect -7227 60999 -7153 61033
rect -7227 60965 -7207 60999
rect -7173 60965 -7153 60999
rect -7227 60931 -7153 60965
rect -7227 60897 -7207 60931
rect -7173 60897 -7153 60931
rect -7227 60863 -7153 60897
rect -7227 60829 -7207 60863
rect -7173 60829 -7153 60863
rect -7227 60795 -7153 60829
rect -7227 60761 -7207 60795
rect -7173 60761 -7153 60795
rect -7227 60727 -7153 60761
rect -7227 60693 -7207 60727
rect -7173 60693 -7153 60727
rect -7227 60659 -7153 60693
rect -7227 60625 -7207 60659
rect -7173 60625 -7153 60659
rect -7227 60591 -7153 60625
rect -7227 60557 -7207 60591
rect -7173 60557 -7153 60591
rect -7227 60523 -7153 60557
rect -7227 60489 -7207 60523
rect -7173 60489 -7153 60523
rect -7227 60455 -7153 60489
rect -7227 60421 -7207 60455
rect -7173 60421 -7153 60455
rect -7227 60387 -7153 60421
rect -7227 60353 -7207 60387
rect -7173 60353 -7153 60387
rect -7227 60319 -7153 60353
rect -7227 60285 -7207 60319
rect -7173 60285 -7153 60319
rect -7227 60251 -7153 60285
rect -7227 60217 -7207 60251
rect -7173 60217 -7153 60251
rect -7227 60183 -7153 60217
rect -7227 60149 -7207 60183
rect -7173 60149 -7153 60183
rect -7227 60115 -7153 60149
rect -7227 60081 -7207 60115
rect -7173 60081 -7153 60115
rect -7227 60047 -7153 60081
rect -7227 60013 -7207 60047
rect -7173 60013 -7153 60047
rect -7227 59979 -7153 60013
rect -7227 59945 -7207 59979
rect -7173 59945 -7153 59979
rect -7227 59911 -7153 59945
rect -7227 59877 -7207 59911
rect -7173 59877 -7153 59911
rect -7227 59843 -7153 59877
rect -7227 59809 -7207 59843
rect -7173 59809 -7153 59843
rect -7227 59775 -7153 59809
rect -7227 59741 -7207 59775
rect -7173 59741 -7153 59775
rect -7227 59707 -7153 59741
rect -7227 59673 -7207 59707
rect -7173 59673 -7153 59707
rect -7227 59639 -7153 59673
rect -7227 59605 -7207 59639
rect -7173 59605 -7153 59639
rect -7227 59571 -7153 59605
rect -7227 59537 -7207 59571
rect -7173 59537 -7153 59571
rect -7227 59503 -7153 59537
rect -7227 59469 -7207 59503
rect -7173 59469 -7153 59503
rect -7227 59435 -7153 59469
rect -7227 59401 -7207 59435
rect -7173 59401 -7153 59435
rect -7227 59367 -7153 59401
rect -7227 59333 -7207 59367
rect -7173 59333 -7153 59367
rect -7227 59299 -7153 59333
rect -7227 59265 -7207 59299
rect -7173 59265 -7153 59299
rect -7227 59231 -7153 59265
rect -7227 59197 -7207 59231
rect -7173 59197 -7153 59231
rect -7227 59163 -7153 59197
rect -7227 59129 -7207 59163
rect -7173 59129 -7153 59163
rect -7227 59095 -7153 59129
rect -7227 59061 -7207 59095
rect -7173 59061 -7153 59095
rect -7227 59027 -7153 59061
rect -7227 58993 -7207 59027
rect -7173 58993 -7153 59027
rect -7227 58959 -7153 58993
rect -7227 58925 -7207 58959
rect -7173 58925 -7153 58959
rect -7227 58891 -7153 58925
rect -7227 58857 -7207 58891
rect -7173 58857 -7153 58891
rect -7227 58823 -7153 58857
rect -7227 58789 -7207 58823
rect -7173 58789 -7153 58823
rect -7227 58755 -7153 58789
rect -7227 58721 -7207 58755
rect -7173 58721 -7153 58755
rect -7227 58687 -7153 58721
rect -7227 58653 -7207 58687
rect -7173 58653 -7153 58687
rect -7227 58619 -7153 58653
rect -7227 58585 -7207 58619
rect -7173 58585 -7153 58619
rect -7227 58551 -7153 58585
rect -7227 58517 -7207 58551
rect -7173 58517 -7153 58551
rect -7227 58483 -7153 58517
rect -7227 58449 -7207 58483
rect -7173 58449 -7153 58483
rect -7227 58415 -7153 58449
rect -7227 58381 -7207 58415
rect -7173 58381 -7153 58415
rect -7227 58347 -7153 58381
rect -7227 58313 -7207 58347
rect -7173 58313 -7153 58347
rect -7227 58279 -7153 58313
rect -7227 58245 -7207 58279
rect -7173 58245 -7153 58279
rect -7227 58211 -7153 58245
rect -7227 58177 -7207 58211
rect -7173 58177 -7153 58211
rect -7227 58143 -7153 58177
rect -7227 58109 -7207 58143
rect -7173 58109 -7153 58143
rect -7227 58075 -7153 58109
rect -7227 58041 -7207 58075
rect -7173 58041 -7153 58075
rect -7227 58007 -7153 58041
rect -7227 57973 -7207 58007
rect -7173 57973 -7153 58007
rect -7227 57939 -7153 57973
rect -7227 57905 -7207 57939
rect -7173 57905 -7153 57939
rect -7227 57871 -7153 57905
rect -7227 57837 -7207 57871
rect -7173 57837 -7153 57871
rect -7227 57803 -7153 57837
rect -7227 57769 -7207 57803
rect -7173 57769 -7153 57803
rect -7227 57735 -7153 57769
rect -7227 57701 -7207 57735
rect -7173 57701 -7153 57735
rect -7227 57667 -7153 57701
rect -7227 57633 -7207 57667
rect -7173 57633 -7153 57667
rect -7227 57599 -7153 57633
rect -7227 57565 -7207 57599
rect -7173 57565 -7153 57599
rect -7227 57531 -7153 57565
rect -7227 57497 -7207 57531
rect -7173 57497 -7153 57531
rect -7227 57463 -7153 57497
rect -7227 57429 -7207 57463
rect -7173 57429 -7153 57463
rect -7227 57395 -7153 57429
rect -7227 57361 -7207 57395
rect -7173 57361 -7153 57395
rect -7227 57327 -7153 57361
rect -7227 57293 -7207 57327
rect -7173 57293 -7153 57327
rect -7227 57259 -7153 57293
rect -7227 57225 -7207 57259
rect -7173 57225 -7153 57259
rect -7227 57191 -7153 57225
rect -7227 57157 -7207 57191
rect -7173 57157 -7153 57191
rect -7227 57123 -7153 57157
rect -7227 57089 -7207 57123
rect -7173 57089 -7153 57123
rect -7227 57055 -7153 57089
rect -7227 57021 -7207 57055
rect -7173 57021 -7153 57055
rect -7227 56987 -7153 57021
rect -7227 56953 -7207 56987
rect -7173 56953 -7153 56987
rect -7227 56919 -7153 56953
rect -7227 56885 -7207 56919
rect -7173 56885 -7153 56919
rect -7227 56851 -7153 56885
rect -7227 56817 -7207 56851
rect -7173 56817 -7153 56851
rect -7227 56783 -7153 56817
rect -7227 56749 -7207 56783
rect -7173 56749 -7153 56783
rect -7227 56715 -7153 56749
rect -7227 56681 -7207 56715
rect -7173 56681 -7153 56715
rect -7227 56647 -7153 56681
rect -7227 56613 -7207 56647
rect -7173 56613 -7153 56647
rect -7227 56579 -7153 56613
rect -7227 56545 -7207 56579
rect -7173 56545 -7153 56579
rect -7227 56511 -7153 56545
rect -7227 56477 -7207 56511
rect -7173 56477 -7153 56511
rect -7227 56443 -7153 56477
rect -7227 56409 -7207 56443
rect -7173 56409 -7153 56443
rect -7227 56375 -7153 56409
rect -7227 56341 -7207 56375
rect -7173 56341 -7153 56375
rect -7227 56324 -7153 56341
rect -10719 56304 -7153 56324
rect -10719 56270 -10614 56304
rect -10580 56270 -10546 56304
rect -10512 56270 -10478 56304
rect -10444 56270 -10410 56304
rect -10376 56270 -10342 56304
rect -10308 56270 -10274 56304
rect -10240 56270 -10206 56304
rect -10172 56270 -10138 56304
rect -10104 56270 -10070 56304
rect -10036 56270 -10002 56304
rect -9968 56270 -9934 56304
rect -9900 56270 -9866 56304
rect -9832 56270 -9798 56304
rect -9764 56270 -9730 56304
rect -9696 56270 -9662 56304
rect -9628 56270 -9594 56304
rect -9560 56270 -9526 56304
rect -9492 56270 -9458 56304
rect -9424 56270 -9390 56304
rect -9356 56270 -9322 56304
rect -9288 56270 -9254 56304
rect -9220 56270 -9186 56304
rect -9152 56270 -9118 56304
rect -9084 56270 -9050 56304
rect -9016 56270 -8982 56304
rect -8948 56270 -8914 56304
rect -8880 56270 -8846 56304
rect -8812 56270 -8778 56304
rect -8744 56270 -8710 56304
rect -8676 56270 -8642 56304
rect -8608 56270 -8574 56304
rect -8540 56270 -8506 56304
rect -8472 56270 -8438 56304
rect -8404 56270 -8370 56304
rect -8336 56270 -8302 56304
rect -8268 56270 -8234 56304
rect -8200 56270 -8166 56304
rect -8132 56270 -8098 56304
rect -8064 56270 -8030 56304
rect -7996 56270 -7962 56304
rect -7928 56270 -7894 56304
rect -7860 56270 -7826 56304
rect -7792 56270 -7758 56304
rect -7724 56270 -7690 56304
rect -7656 56270 -7622 56304
rect -7588 56270 -7554 56304
rect -7520 56270 -7486 56304
rect -7452 56270 -7418 56304
rect -7384 56270 -7350 56304
rect -7316 56270 -7282 56304
rect -7248 56270 -7153 56304
rect -10719 56250 -7153 56270
rect -3738 64122 -3718 64156
rect -3684 64122 -3664 64156
rect -3738 64088 -3664 64122
rect -3738 64054 -3718 64088
rect -3684 64054 -3664 64088
rect -3738 64020 -3664 64054
rect -3738 63986 -3718 64020
rect -3684 63986 -3664 64020
rect -3738 63952 -3664 63986
rect -3738 63918 -3718 63952
rect -3684 63918 -3664 63952
rect -3738 63884 -3664 63918
rect -3738 63850 -3718 63884
rect -3684 63850 -3664 63884
rect -3738 63816 -3664 63850
rect -3738 63782 -3718 63816
rect -3684 63782 -3664 63816
rect -3738 63748 -3664 63782
rect -3738 63714 -3718 63748
rect -3684 63714 -3664 63748
rect -3738 63680 -3664 63714
rect -3738 63646 -3718 63680
rect -3684 63646 -3664 63680
rect -3738 63612 -3664 63646
rect -3738 63578 -3718 63612
rect -3684 63578 -3664 63612
rect -3738 63544 -3664 63578
rect -3738 63510 -3718 63544
rect -3684 63510 -3664 63544
rect -3738 63476 -3664 63510
rect -3738 63442 -3718 63476
rect -3684 63442 -3664 63476
rect -3738 63408 -3664 63442
rect -3738 63374 -3718 63408
rect -3684 63374 -3664 63408
rect -3738 63340 -3664 63374
rect -3738 63306 -3718 63340
rect -3684 63306 -3664 63340
rect -3738 63272 -3664 63306
rect -3738 63238 -3718 63272
rect -3684 63238 -3664 63272
rect -3738 63204 -3664 63238
rect -3738 63170 -3718 63204
rect -3684 63170 -3664 63204
rect -3738 63136 -3664 63170
rect -3738 63102 -3718 63136
rect -3684 63102 -3664 63136
rect -3738 63068 -3664 63102
rect -3738 63034 -3718 63068
rect -3684 63034 -3664 63068
rect -3738 63000 -3664 63034
rect -3738 62966 -3718 63000
rect -3684 62966 -3664 63000
rect -3738 62932 -3664 62966
rect -3738 62898 -3718 62932
rect -3684 62898 -3664 62932
rect -3738 62864 -3664 62898
rect -3738 62830 -3718 62864
rect -3684 62830 -3664 62864
rect -3738 62796 -3664 62830
rect -3738 62762 -3718 62796
rect -3684 62762 -3664 62796
rect -3738 62728 -3664 62762
rect -3738 62694 -3718 62728
rect -3684 62694 -3664 62728
rect -3738 62660 -3664 62694
rect -3738 62626 -3718 62660
rect -3684 62626 -3664 62660
rect -3738 62592 -3664 62626
rect -3738 62558 -3718 62592
rect -3684 62558 -3664 62592
rect -3738 62524 -3664 62558
rect -3738 62490 -3718 62524
rect -3684 62490 -3664 62524
rect -3738 62456 -3664 62490
rect -3738 62422 -3718 62456
rect -3684 62422 -3664 62456
rect -3738 62388 -3664 62422
rect -3738 62354 -3718 62388
rect -3684 62354 -3664 62388
rect -3738 62320 -3664 62354
rect -3738 62286 -3718 62320
rect -3684 62286 -3664 62320
rect -3738 62252 -3664 62286
rect -3738 62218 -3718 62252
rect -3684 62218 -3664 62252
rect -3738 62184 -3664 62218
rect -3738 62150 -3718 62184
rect -3684 62150 -3664 62184
rect -3738 62116 -3664 62150
rect -3738 62082 -3718 62116
rect -3684 62082 -3664 62116
rect -3738 62048 -3664 62082
rect 59084 74806 70892 74826
rect 59084 74772 59191 74806
rect 59225 74772 59259 74806
rect 59293 74772 59327 74806
rect 59361 74772 59395 74806
rect 59429 74772 59463 74806
rect 59497 74772 59531 74806
rect 59565 74772 59599 74806
rect 59633 74772 59667 74806
rect 59701 74772 59735 74806
rect 59769 74772 59803 74806
rect 59837 74772 59871 74806
rect 59905 74772 59939 74806
rect 59973 74772 60007 74806
rect 60041 74772 60075 74806
rect 60109 74772 60143 74806
rect 60177 74772 60211 74806
rect 60245 74772 60279 74806
rect 60313 74772 60347 74806
rect 60381 74772 60415 74806
rect 60449 74772 60483 74806
rect 60517 74772 60551 74806
rect 60585 74772 60619 74806
rect 60653 74772 60687 74806
rect 60721 74772 60755 74806
rect 60789 74772 60823 74806
rect 60857 74772 60891 74806
rect 60925 74772 60959 74806
rect 60993 74772 61027 74806
rect 61061 74772 61095 74806
rect 61129 74772 61163 74806
rect 61197 74772 61231 74806
rect 61265 74772 61299 74806
rect 61333 74772 61367 74806
rect 61401 74772 61435 74806
rect 61469 74772 61503 74806
rect 61537 74772 61571 74806
rect 61605 74772 61639 74806
rect 61673 74772 61707 74806
rect 61741 74772 61775 74806
rect 61809 74772 61843 74806
rect 61877 74772 61911 74806
rect 61945 74772 61979 74806
rect 62013 74772 62047 74806
rect 62081 74772 62115 74806
rect 62149 74772 62183 74806
rect 62217 74772 62251 74806
rect 62285 74772 62319 74806
rect 62353 74772 62387 74806
rect 62421 74772 62455 74806
rect 62489 74772 62523 74806
rect 62557 74772 62591 74806
rect 62625 74772 62659 74806
rect 62693 74772 62727 74806
rect 62761 74772 62795 74806
rect 62829 74772 62863 74806
rect 62897 74772 62931 74806
rect 62965 74772 62999 74806
rect 63033 74772 63067 74806
rect 63101 74772 63135 74806
rect 63169 74772 63203 74806
rect 63237 74772 63271 74806
rect 63305 74772 63339 74806
rect 63373 74772 63407 74806
rect 63441 74772 63475 74806
rect 63509 74772 63543 74806
rect 63577 74772 63611 74806
rect 63645 74772 63679 74806
rect 63713 74772 63747 74806
rect 63781 74772 63815 74806
rect 63849 74772 63883 74806
rect 63917 74772 63951 74806
rect 63985 74772 64019 74806
rect 64053 74772 64087 74806
rect 64121 74772 64155 74806
rect 64189 74772 64223 74806
rect 64257 74772 64291 74806
rect 64325 74772 64359 74806
rect 64393 74772 64427 74806
rect 64461 74772 64495 74806
rect 64529 74772 64563 74806
rect 64597 74772 64631 74806
rect 64665 74772 64699 74806
rect 64733 74772 64767 74806
rect 64801 74772 64835 74806
rect 64869 74772 64903 74806
rect 64937 74772 64971 74806
rect 65005 74772 65039 74806
rect 65073 74772 65107 74806
rect 65141 74772 65175 74806
rect 65209 74772 65243 74806
rect 65277 74772 65311 74806
rect 65345 74772 65379 74806
rect 65413 74772 65447 74806
rect 65481 74772 65515 74806
rect 65549 74772 65583 74806
rect 65617 74772 65651 74806
rect 65685 74772 65719 74806
rect 65753 74772 65787 74806
rect 65821 74772 65855 74806
rect 65889 74772 65923 74806
rect 65957 74772 65991 74806
rect 66025 74772 66059 74806
rect 66093 74772 66127 74806
rect 66161 74772 66195 74806
rect 66229 74772 66263 74806
rect 66297 74772 66331 74806
rect 66365 74772 66399 74806
rect 66433 74772 66467 74806
rect 66501 74772 66535 74806
rect 66569 74772 66603 74806
rect 66637 74772 66671 74806
rect 66705 74772 66739 74806
rect 66773 74772 66807 74806
rect 66841 74772 66875 74806
rect 66909 74772 66943 74806
rect 66977 74772 67011 74806
rect 67045 74772 67079 74806
rect 67113 74772 67147 74806
rect 67181 74772 67215 74806
rect 67249 74772 67283 74806
rect 67317 74772 67351 74806
rect 67385 74772 67419 74806
rect 67453 74772 67487 74806
rect 67521 74772 67555 74806
rect 67589 74772 67623 74806
rect 67657 74772 67691 74806
rect 67725 74772 67759 74806
rect 67793 74772 67827 74806
rect 67861 74772 67895 74806
rect 67929 74772 67963 74806
rect 67997 74772 68031 74806
rect 68065 74772 68099 74806
rect 68133 74772 68167 74806
rect 68201 74772 68235 74806
rect 68269 74772 68303 74806
rect 68337 74772 68371 74806
rect 68405 74772 68439 74806
rect 68473 74772 68507 74806
rect 68541 74772 68575 74806
rect 68609 74772 68643 74806
rect 68677 74772 68711 74806
rect 68745 74772 68779 74806
rect 68813 74772 68847 74806
rect 68881 74772 68915 74806
rect 68949 74772 68983 74806
rect 69017 74772 69051 74806
rect 69085 74772 69119 74806
rect 69153 74772 69187 74806
rect 69221 74772 69255 74806
rect 69289 74772 69323 74806
rect 69357 74772 69391 74806
rect 69425 74772 69459 74806
rect 69493 74772 69527 74806
rect 69561 74772 69595 74806
rect 69629 74772 69663 74806
rect 69697 74772 69731 74806
rect 69765 74772 69799 74806
rect 69833 74772 69867 74806
rect 69901 74772 69935 74806
rect 69969 74772 70003 74806
rect 70037 74772 70071 74806
rect 70105 74772 70139 74806
rect 70173 74772 70207 74806
rect 70241 74772 70275 74806
rect 70309 74772 70343 74806
rect 70377 74772 70411 74806
rect 70445 74772 70479 74806
rect 70513 74772 70547 74806
rect 70581 74772 70615 74806
rect 70649 74772 70683 74806
rect 70717 74772 70751 74806
rect 70785 74772 70892 74806
rect 59084 74752 70892 74772
rect 59084 74745 59158 74752
rect 59084 74711 59104 74745
rect 59138 74711 59158 74745
rect 59084 74677 59158 74711
rect 59084 74643 59104 74677
rect 59138 74643 59158 74677
rect 59084 74609 59158 74643
rect 59084 74575 59104 74609
rect 59138 74575 59158 74609
rect 59084 74541 59158 74575
rect 59084 74507 59104 74541
rect 59138 74507 59158 74541
rect 59084 74473 59158 74507
rect 59084 74439 59104 74473
rect 59138 74439 59158 74473
rect 59084 74405 59158 74439
rect 59084 74371 59104 74405
rect 59138 74371 59158 74405
rect 59084 74337 59158 74371
rect 59084 74303 59104 74337
rect 59138 74303 59158 74337
rect 59084 74269 59158 74303
rect 59084 74235 59104 74269
rect 59138 74235 59158 74269
rect 59084 74201 59158 74235
rect 59084 74167 59104 74201
rect 59138 74167 59158 74201
rect 59084 74133 59158 74167
rect 59084 74099 59104 74133
rect 59138 74099 59158 74133
rect 59084 74065 59158 74099
rect 59084 74031 59104 74065
rect 59138 74031 59158 74065
rect 59084 73997 59158 74031
rect 59084 73963 59104 73997
rect 59138 73963 59158 73997
rect 59084 73929 59158 73963
rect 59084 73895 59104 73929
rect 59138 73895 59158 73929
rect 59084 73861 59158 73895
rect 59084 73827 59104 73861
rect 59138 73827 59158 73861
rect 59084 73793 59158 73827
rect 59084 73759 59104 73793
rect 59138 73759 59158 73793
rect 59084 73725 59158 73759
rect 59084 73691 59104 73725
rect 59138 73691 59158 73725
rect 59084 73657 59158 73691
rect 59084 73623 59104 73657
rect 59138 73623 59158 73657
rect 59084 73589 59158 73623
rect 59084 73555 59104 73589
rect 59138 73555 59158 73589
rect 59084 73521 59158 73555
rect 59084 73487 59104 73521
rect 59138 73487 59158 73521
rect 59084 73453 59158 73487
rect 59084 73419 59104 73453
rect 59138 73419 59158 73453
rect 59084 73385 59158 73419
rect 59084 73351 59104 73385
rect 59138 73351 59158 73385
rect 59084 73317 59158 73351
rect 59084 73283 59104 73317
rect 59138 73283 59158 73317
rect 59084 73249 59158 73283
rect 59084 73215 59104 73249
rect 59138 73215 59158 73249
rect 59084 73181 59158 73215
rect 59084 73147 59104 73181
rect 59138 73147 59158 73181
rect 59084 73113 59158 73147
rect 59084 73079 59104 73113
rect 59138 73079 59158 73113
rect 59084 73045 59158 73079
rect 59084 73011 59104 73045
rect 59138 73011 59158 73045
rect 59084 72977 59158 73011
rect 59084 72943 59104 72977
rect 59138 72943 59158 72977
rect 59084 72909 59158 72943
rect 59084 72875 59104 72909
rect 59138 72875 59158 72909
rect 59084 72841 59158 72875
rect 59084 72807 59104 72841
rect 59138 72807 59158 72841
rect 59084 72773 59158 72807
rect 59084 72739 59104 72773
rect 59138 72739 59158 72773
rect 59084 72705 59158 72739
rect 59084 72671 59104 72705
rect 59138 72671 59158 72705
rect 59084 72637 59158 72671
rect 59084 72603 59104 72637
rect 59138 72603 59158 72637
rect 59084 72569 59158 72603
rect 59084 72535 59104 72569
rect 59138 72535 59158 72569
rect 59084 72501 59158 72535
rect 59084 72467 59104 72501
rect 59138 72467 59158 72501
rect 59084 72433 59158 72467
rect 59084 72399 59104 72433
rect 59138 72399 59158 72433
rect 59084 72365 59158 72399
rect 59084 72331 59104 72365
rect 59138 72331 59158 72365
rect 59084 72297 59158 72331
rect 59084 72263 59104 72297
rect 59138 72263 59158 72297
rect 59084 72229 59158 72263
rect 59084 72195 59104 72229
rect 59138 72195 59158 72229
rect 59084 72161 59158 72195
rect 59084 72127 59104 72161
rect 59138 72127 59158 72161
rect 59084 72093 59158 72127
rect 59084 72059 59104 72093
rect 59138 72059 59158 72093
rect 59084 72025 59158 72059
rect 59084 71991 59104 72025
rect 59138 71991 59158 72025
rect 59084 71957 59158 71991
rect 59084 71923 59104 71957
rect 59138 71923 59158 71957
rect 59084 71889 59158 71923
rect 59084 71855 59104 71889
rect 59138 71855 59158 71889
rect 59084 71821 59158 71855
rect 59084 71787 59104 71821
rect 59138 71787 59158 71821
rect 59084 71753 59158 71787
rect 59084 71719 59104 71753
rect 59138 71719 59158 71753
rect 59084 71685 59158 71719
rect 59084 71651 59104 71685
rect 59138 71651 59158 71685
rect 59084 71617 59158 71651
rect 59084 71583 59104 71617
rect 59138 71583 59158 71617
rect 59084 71549 59158 71583
rect 59084 71515 59104 71549
rect 59138 71515 59158 71549
rect 59084 71481 59158 71515
rect 59084 71447 59104 71481
rect 59138 71447 59158 71481
rect 59084 71413 59158 71447
rect 59084 71379 59104 71413
rect 59138 71379 59158 71413
rect 59084 71345 59158 71379
rect 59084 71311 59104 71345
rect 59138 71311 59158 71345
rect 59084 71277 59158 71311
rect 59084 71243 59104 71277
rect 59138 71243 59158 71277
rect 59084 71209 59158 71243
rect 59084 71175 59104 71209
rect 59138 71175 59158 71209
rect 59084 71141 59158 71175
rect 59084 71107 59104 71141
rect 59138 71107 59158 71141
rect 59084 71073 59158 71107
rect 59084 71039 59104 71073
rect 59138 71039 59158 71073
rect 59084 71005 59158 71039
rect 59084 70971 59104 71005
rect 59138 70971 59158 71005
rect 59084 70937 59158 70971
rect 59084 70903 59104 70937
rect 59138 70903 59158 70937
rect 59084 70869 59158 70903
rect 59084 70835 59104 70869
rect 59138 70835 59158 70869
rect 59084 70801 59158 70835
rect 59084 70767 59104 70801
rect 59138 70767 59158 70801
rect 59084 70733 59158 70767
rect 59084 70699 59104 70733
rect 59138 70699 59158 70733
rect 59084 70665 59158 70699
rect 59084 70631 59104 70665
rect 59138 70631 59158 70665
rect 59084 70597 59158 70631
rect 59084 70563 59104 70597
rect 59138 70563 59158 70597
rect 59084 70529 59158 70563
rect 59084 70495 59104 70529
rect 59138 70495 59158 70529
rect 59084 70461 59158 70495
rect 59084 70427 59104 70461
rect 59138 70427 59158 70461
rect 59084 70393 59158 70427
rect 59084 70359 59104 70393
rect 59138 70359 59158 70393
rect 59084 70325 59158 70359
rect 59084 70291 59104 70325
rect 59138 70291 59158 70325
rect 59084 70257 59158 70291
rect 59084 70223 59104 70257
rect 59138 70223 59158 70257
rect 59084 70189 59158 70223
rect 59084 70155 59104 70189
rect 59138 70155 59158 70189
rect 59084 70121 59158 70155
rect 59084 70087 59104 70121
rect 59138 70087 59158 70121
rect 59084 70053 59158 70087
rect 59084 70019 59104 70053
rect 59138 70019 59158 70053
rect 59084 69985 59158 70019
rect 59084 69951 59104 69985
rect 59138 69951 59158 69985
rect 59084 69917 59158 69951
rect 59084 69883 59104 69917
rect 59138 69883 59158 69917
rect 59084 69849 59158 69883
rect 59084 69815 59104 69849
rect 59138 69815 59158 69849
rect 59084 69781 59158 69815
rect 59084 69747 59104 69781
rect 59138 69747 59158 69781
rect 59084 69713 59158 69747
rect 59084 69679 59104 69713
rect 59138 69679 59158 69713
rect 59084 69645 59158 69679
rect 59084 69611 59104 69645
rect 59138 69611 59158 69645
rect 59084 69577 59158 69611
rect 59084 69543 59104 69577
rect 59138 69543 59158 69577
rect 59084 69509 59158 69543
rect 59084 69475 59104 69509
rect 59138 69475 59158 69509
rect 59084 69441 59158 69475
rect 59084 69407 59104 69441
rect 59138 69407 59158 69441
rect 59084 69373 59158 69407
rect 59084 69339 59104 69373
rect 59138 69339 59158 69373
rect 59084 69305 59158 69339
rect 59084 69271 59104 69305
rect 59138 69271 59158 69305
rect 59084 69237 59158 69271
rect 59084 69203 59104 69237
rect 59138 69203 59158 69237
rect 59084 69169 59158 69203
rect 59084 69135 59104 69169
rect 59138 69135 59158 69169
rect 59084 69101 59158 69135
rect 59084 69067 59104 69101
rect 59138 69067 59158 69101
rect 59084 69033 59158 69067
rect 59084 68999 59104 69033
rect 59138 68999 59158 69033
rect 59084 68965 59158 68999
rect 59084 68931 59104 68965
rect 59138 68931 59158 68965
rect 59084 68897 59158 68931
rect 59084 68863 59104 68897
rect 59138 68863 59158 68897
rect 59084 68829 59158 68863
rect 59084 68795 59104 68829
rect 59138 68795 59158 68829
rect 59084 68761 59158 68795
rect 59084 68727 59104 68761
rect 59138 68727 59158 68761
rect 59084 68693 59158 68727
rect 59084 68659 59104 68693
rect 59138 68659 59158 68693
rect 59084 68625 59158 68659
rect 59084 68591 59104 68625
rect 59138 68591 59158 68625
rect 59084 68557 59158 68591
rect 59084 68523 59104 68557
rect 59138 68523 59158 68557
rect 59084 68489 59158 68523
rect 59084 68455 59104 68489
rect 59138 68455 59158 68489
rect 59084 68421 59158 68455
rect 59084 68387 59104 68421
rect 59138 68387 59158 68421
rect 59084 68353 59158 68387
rect 59084 68319 59104 68353
rect 59138 68319 59158 68353
rect 59084 68285 59158 68319
rect 59084 68251 59104 68285
rect 59138 68251 59158 68285
rect 59084 68217 59158 68251
rect 59084 68183 59104 68217
rect 59138 68183 59158 68217
rect 59084 68149 59158 68183
rect 59084 68115 59104 68149
rect 59138 68115 59158 68149
rect 59084 68081 59158 68115
rect 59084 68047 59104 68081
rect 59138 68047 59158 68081
rect 59084 68013 59158 68047
rect 59084 67979 59104 68013
rect 59138 67979 59158 68013
rect 59084 67945 59158 67979
rect 59084 67911 59104 67945
rect 59138 67911 59158 67945
rect 59084 67877 59158 67911
rect 59084 67843 59104 67877
rect 59138 67843 59158 67877
rect 59084 67809 59158 67843
rect 59084 67775 59104 67809
rect 59138 67775 59158 67809
rect 59084 67741 59158 67775
rect 59084 67707 59104 67741
rect 59138 67707 59158 67741
rect 59084 67673 59158 67707
rect 59084 67639 59104 67673
rect 59138 67639 59158 67673
rect 59084 67605 59158 67639
rect 59084 67571 59104 67605
rect 59138 67571 59158 67605
rect 59084 67537 59158 67571
rect 59084 67503 59104 67537
rect 59138 67503 59158 67537
rect 59084 67469 59158 67503
rect 59084 67435 59104 67469
rect 59138 67435 59158 67469
rect 59084 67401 59158 67435
rect 59084 67367 59104 67401
rect 59138 67367 59158 67401
rect 59084 67333 59158 67367
rect 59084 67299 59104 67333
rect 59138 67299 59158 67333
rect 59084 67265 59158 67299
rect 59084 67231 59104 67265
rect 59138 67231 59158 67265
rect 59084 67197 59158 67231
rect 59084 67163 59104 67197
rect 59138 67163 59158 67197
rect 59084 67129 59158 67163
rect 59084 67095 59104 67129
rect 59138 67095 59158 67129
rect 59084 67061 59158 67095
rect 59084 67027 59104 67061
rect 59138 67027 59158 67061
rect 59084 66993 59158 67027
rect 59084 66959 59104 66993
rect 59138 66959 59158 66993
rect 59084 66925 59158 66959
rect 59084 66891 59104 66925
rect 59138 66891 59158 66925
rect 59084 66857 59158 66891
rect 59084 66823 59104 66857
rect 59138 66823 59158 66857
rect 59084 66789 59158 66823
rect 59084 66755 59104 66789
rect 59138 66755 59158 66789
rect 59084 66721 59158 66755
rect 59084 66687 59104 66721
rect 59138 66687 59158 66721
rect 59084 66653 59158 66687
rect 59084 66619 59104 66653
rect 59138 66619 59158 66653
rect 59084 66585 59158 66619
rect 59084 66551 59104 66585
rect 59138 66551 59158 66585
rect 59084 66517 59158 66551
rect 59084 66483 59104 66517
rect 59138 66483 59158 66517
rect 59084 66449 59158 66483
rect 59084 66415 59104 66449
rect 59138 66415 59158 66449
rect 59084 66381 59158 66415
rect 59084 66347 59104 66381
rect 59138 66347 59158 66381
rect 59084 66313 59158 66347
rect 59084 66279 59104 66313
rect 59138 66279 59158 66313
rect 59084 66245 59158 66279
rect 59084 66211 59104 66245
rect 59138 66211 59158 66245
rect 59084 66177 59158 66211
rect 59084 66143 59104 66177
rect 59138 66143 59158 66177
rect 59084 66109 59158 66143
rect 59084 66075 59104 66109
rect 59138 66075 59158 66109
rect 59084 66041 59158 66075
rect 59084 66007 59104 66041
rect 59138 66007 59158 66041
rect 59084 65973 59158 66007
rect 59084 65939 59104 65973
rect 59138 65939 59158 65973
rect 59084 65905 59158 65939
rect 59084 65871 59104 65905
rect 59138 65871 59158 65905
rect 59084 65837 59158 65871
rect 59084 65803 59104 65837
rect 59138 65803 59158 65837
rect 59084 65769 59158 65803
rect 59084 65735 59104 65769
rect 59138 65735 59158 65769
rect 59084 65701 59158 65735
rect 59084 65667 59104 65701
rect 59138 65667 59158 65701
rect 59084 65633 59158 65667
rect 59084 65599 59104 65633
rect 59138 65599 59158 65633
rect 59084 65565 59158 65599
rect 59084 65531 59104 65565
rect 59138 65531 59158 65565
rect 59084 65497 59158 65531
rect 59084 65463 59104 65497
rect 59138 65463 59158 65497
rect 59084 65429 59158 65463
rect 59084 65395 59104 65429
rect 59138 65395 59158 65429
rect 59084 65361 59158 65395
rect 59084 65327 59104 65361
rect 59138 65327 59158 65361
rect 59084 65293 59158 65327
rect 59084 65259 59104 65293
rect 59138 65259 59158 65293
rect 59084 65225 59158 65259
rect 59084 65191 59104 65225
rect 59138 65191 59158 65225
rect 59084 65157 59158 65191
rect 59084 65123 59104 65157
rect 59138 65123 59158 65157
rect 59084 65089 59158 65123
rect 59084 65055 59104 65089
rect 59138 65055 59158 65089
rect 59084 65021 59158 65055
rect 59084 64987 59104 65021
rect 59138 64987 59158 65021
rect 59084 64953 59158 64987
rect 59084 64919 59104 64953
rect 59138 64919 59158 64953
rect 59084 64885 59158 64919
rect 59084 64851 59104 64885
rect 59138 64851 59158 64885
rect 59084 64817 59158 64851
rect 59084 64783 59104 64817
rect 59138 64783 59158 64817
rect 59084 64749 59158 64783
rect 59084 64715 59104 64749
rect 59138 64715 59158 64749
rect 59084 64681 59158 64715
rect 59084 64647 59104 64681
rect 59138 64647 59158 64681
rect 59084 64613 59158 64647
rect 59084 64579 59104 64613
rect 59138 64579 59158 64613
rect 59084 64545 59158 64579
rect 59084 64511 59104 64545
rect 59138 64511 59158 64545
rect 59084 64477 59158 64511
rect 59084 64443 59104 64477
rect 59138 64443 59158 64477
rect 59084 64409 59158 64443
rect 59084 64375 59104 64409
rect 59138 64375 59158 64409
rect 59084 64341 59158 64375
rect 59084 64307 59104 64341
rect 59138 64307 59158 64341
rect 59084 64273 59158 64307
rect 59084 64239 59104 64273
rect 59138 64239 59158 64273
rect 59084 64205 59158 64239
rect 59084 64171 59104 64205
rect 59138 64171 59158 64205
rect 59084 64137 59158 64171
rect 59084 64103 59104 64137
rect 59138 64103 59158 64137
rect 59084 64069 59158 64103
rect 59084 64035 59104 64069
rect 59138 64035 59158 64069
rect 59084 64001 59158 64035
rect 59084 63967 59104 64001
rect 59138 63967 59158 64001
rect 59084 63933 59158 63967
rect 59084 63899 59104 63933
rect 59138 63899 59158 63933
rect 59084 63865 59158 63899
rect 59084 63831 59104 63865
rect 59138 63831 59158 63865
rect 59084 63797 59158 63831
rect 59084 63763 59104 63797
rect 59138 63763 59158 63797
rect 59084 63729 59158 63763
rect 59084 63695 59104 63729
rect 59138 63695 59158 63729
rect 59084 63661 59158 63695
rect 59084 63627 59104 63661
rect 59138 63627 59158 63661
rect 59084 63593 59158 63627
rect 59084 63559 59104 63593
rect 59138 63559 59158 63593
rect 59084 63525 59158 63559
rect 59084 63491 59104 63525
rect 59138 63491 59158 63525
rect 59084 63457 59158 63491
rect 59084 63423 59104 63457
rect 59138 63423 59158 63457
rect 59084 63389 59158 63423
rect 59084 63355 59104 63389
rect 59138 63355 59158 63389
rect 59084 63321 59158 63355
rect 59084 63287 59104 63321
rect 59138 63287 59158 63321
rect 59084 63253 59158 63287
rect 59084 63219 59104 63253
rect 59138 63219 59158 63253
rect 59084 63185 59158 63219
rect 59084 63151 59104 63185
rect 59138 63151 59158 63185
rect 59084 63117 59158 63151
rect 59084 63083 59104 63117
rect 59138 63083 59158 63117
rect 59084 63049 59158 63083
rect 59084 63015 59104 63049
rect 59138 63015 59158 63049
rect 59084 62981 59158 63015
rect 59084 62947 59104 62981
rect 59138 62947 59158 62981
rect 59084 62913 59158 62947
rect 59084 62879 59104 62913
rect 59138 62879 59158 62913
rect 59084 62845 59158 62879
rect 59084 62811 59104 62845
rect 59138 62811 59158 62845
rect 59084 62777 59158 62811
rect 59084 62743 59104 62777
rect 59138 62743 59158 62777
rect 59084 62709 59158 62743
rect 59084 62675 59104 62709
rect 59138 62675 59158 62709
rect 59084 62641 59158 62675
rect 59084 62607 59104 62641
rect 59138 62607 59158 62641
rect 59084 62573 59158 62607
rect 59084 62539 59104 62573
rect 59138 62539 59158 62573
rect 59084 62505 59158 62539
rect 59084 62471 59104 62505
rect 59138 62471 59158 62505
rect 59084 62437 59158 62471
rect 59084 62403 59104 62437
rect 59138 62403 59158 62437
rect 59084 62369 59158 62403
rect 59084 62335 59104 62369
rect 59138 62335 59158 62369
rect 59084 62301 59158 62335
rect 59084 62267 59104 62301
rect 59138 62267 59158 62301
rect 59084 62233 59158 62267
rect 59084 62199 59104 62233
rect 59138 62199 59158 62233
rect 59084 62165 59158 62199
rect 59084 62131 59104 62165
rect 59138 62131 59158 62165
rect 59084 62097 59158 62131
rect 59084 62063 59104 62097
rect 59138 62063 59158 62097
rect -3738 62014 -3718 62048
rect -3684 62014 -3664 62048
rect -3738 61980 -3664 62014
rect -3738 61946 -3718 61980
rect -3684 61946 -3664 61980
rect -3738 61912 -3664 61946
rect -3738 61878 -3718 61912
rect -3684 61878 -3664 61912
rect -3738 61844 -3664 61878
rect -3738 61810 -3718 61844
rect -3684 61810 -3664 61844
rect -3738 61776 -3664 61810
rect -3738 61742 -3718 61776
rect -3684 61742 -3664 61776
rect -3738 61708 -3664 61742
rect -3738 61674 -3718 61708
rect -3684 61674 -3664 61708
rect -3738 61640 -3664 61674
rect -3738 61606 -3718 61640
rect -3684 61606 -3664 61640
rect -3738 61572 -3664 61606
rect -3738 61538 -3718 61572
rect -3684 61538 -3664 61572
rect -3738 61504 -3664 61538
rect -3738 61470 -3718 61504
rect -3684 61470 -3664 61504
rect -3738 61436 -3664 61470
rect -3738 61402 -3718 61436
rect -3684 61402 -3664 61436
rect -3738 61368 -3664 61402
rect -3738 61334 -3718 61368
rect -3684 61334 -3664 61368
rect -3738 61300 -3664 61334
rect -3738 61266 -3718 61300
rect -3684 61266 -3664 61300
rect -3738 61232 -3664 61266
rect -3738 61198 -3718 61232
rect -3684 61198 -3664 61232
rect -3738 61164 -3664 61198
rect -3738 61130 -3718 61164
rect -3684 61130 -3664 61164
rect -3738 61096 -3664 61130
rect -3738 61062 -3718 61096
rect -3684 61062 -3664 61096
rect -3738 61028 -3664 61062
rect -3738 60994 -3718 61028
rect -3684 60994 -3664 61028
rect -3738 60960 -3664 60994
rect -3738 60926 -3718 60960
rect -3684 60926 -3664 60960
rect -3738 60892 -3664 60926
rect -3738 60858 -3718 60892
rect -3684 60858 -3664 60892
rect -3738 60824 -3664 60858
rect -3738 60790 -3718 60824
rect -3684 60790 -3664 60824
rect -3738 60756 -3664 60790
rect -3738 60722 -3718 60756
rect -3684 60722 -3664 60756
rect -3738 60688 -3664 60722
rect -3738 60654 -3718 60688
rect -3684 60654 -3664 60688
rect -3738 60620 -3664 60654
rect -3738 60586 -3718 60620
rect -3684 60586 -3664 60620
rect -3738 60552 -3664 60586
rect -3738 60518 -3718 60552
rect -3684 60518 -3664 60552
rect -3738 60484 -3664 60518
rect -3738 60450 -3718 60484
rect -3684 60450 -3664 60484
rect -3738 60416 -3664 60450
rect -3738 60382 -3718 60416
rect -3684 60382 -3664 60416
rect -3738 60348 -3664 60382
rect -3738 60314 -3718 60348
rect -3684 60314 -3664 60348
rect -3738 60280 -3664 60314
rect -3738 60246 -3718 60280
rect -3684 60246 -3664 60280
rect -3738 60212 -3664 60246
rect -3738 60178 -3718 60212
rect -3684 60178 -3664 60212
rect -3738 60144 -3664 60178
rect -3738 60110 -3718 60144
rect -3684 60110 -3664 60144
rect -3738 60076 -3664 60110
rect -3738 60042 -3718 60076
rect -3684 60042 -3664 60076
rect -3738 60008 -3664 60042
rect -3738 59974 -3718 60008
rect -3684 59974 -3664 60008
rect -3738 59940 -3664 59974
rect -3738 59906 -3718 59940
rect -3684 59906 -3664 59940
rect -3738 59872 -3664 59906
rect -3738 59838 -3718 59872
rect -3684 59838 -3664 59872
rect -3738 59804 -3664 59838
rect -3738 59770 -3718 59804
rect -3684 59770 -3664 59804
rect -3738 59736 -3664 59770
rect -3738 59702 -3718 59736
rect -3684 59702 -3664 59736
rect -3738 59668 -3664 59702
rect -3738 59634 -3718 59668
rect -3684 59634 -3664 59668
rect -3738 59600 -3664 59634
rect -3738 59566 -3718 59600
rect -3684 59566 -3664 59600
rect -3738 59532 -3664 59566
rect -3738 59498 -3718 59532
rect -3684 59498 -3664 59532
rect -3738 59464 -3664 59498
rect -3738 59430 -3718 59464
rect -3684 59430 -3664 59464
rect -3738 59396 -3664 59430
rect -3738 59362 -3718 59396
rect -3684 59362 -3664 59396
rect -3738 59328 -3664 59362
rect -3738 59294 -3718 59328
rect -3684 59294 -3664 59328
rect -3738 59260 -3664 59294
rect -3738 59226 -3718 59260
rect -3684 59226 -3664 59260
rect -3738 59192 -3664 59226
rect -3738 59158 -3718 59192
rect -3684 59158 -3664 59192
rect -3738 59124 -3664 59158
rect -3738 59090 -3718 59124
rect -3684 59090 -3664 59124
rect -3738 59056 -3664 59090
rect -3738 59022 -3718 59056
rect -3684 59022 -3664 59056
rect -3738 58988 -3664 59022
rect -3738 58954 -3718 58988
rect -3684 58954 -3664 58988
rect -3738 58920 -3664 58954
rect -3738 58886 -3718 58920
rect -3684 58886 -3664 58920
rect -3738 58852 -3664 58886
rect -3738 58818 -3718 58852
rect -3684 58818 -3664 58852
rect -3738 58784 -3664 58818
rect -3738 58750 -3718 58784
rect -3684 58750 -3664 58784
rect -3738 58716 -3664 58750
rect -3738 58682 -3718 58716
rect -3684 58682 -3664 58716
rect -3738 58648 -3664 58682
rect -3738 58614 -3718 58648
rect -3684 58614 -3664 58648
rect -3738 58580 -3664 58614
rect -3738 58546 -3718 58580
rect -3684 58546 -3664 58580
rect -3738 58512 -3664 58546
rect -3738 58478 -3718 58512
rect -3684 58478 -3664 58512
rect -3738 58444 -3664 58478
rect -3738 58410 -3718 58444
rect -3684 58410 -3664 58444
rect -3738 58376 -3664 58410
rect -3738 58342 -3718 58376
rect -3684 58342 -3664 58376
rect -3738 58308 -3664 58342
rect 50436 62040 56370 62060
rect 50436 62006 50530 62040
rect 50564 62006 50598 62040
rect 50632 62006 50666 62040
rect 50700 62006 50734 62040
rect 50768 62006 50802 62040
rect 50836 62006 50870 62040
rect 50904 62006 50938 62040
rect 50972 62006 51006 62040
rect 51040 62006 51074 62040
rect 51108 62006 51142 62040
rect 51176 62006 51210 62040
rect 51244 62006 51278 62040
rect 51312 62006 51346 62040
rect 51380 62006 51414 62040
rect 51448 62006 51482 62040
rect 51516 62006 51550 62040
rect 51584 62006 51618 62040
rect 51652 62006 51686 62040
rect 51720 62006 51754 62040
rect 51788 62006 51822 62040
rect 51856 62006 51890 62040
rect 51924 62006 51958 62040
rect 51992 62006 52026 62040
rect 52060 62006 52094 62040
rect 52128 62006 52162 62040
rect 52196 62006 52230 62040
rect 52264 62006 52298 62040
rect 52332 62006 52366 62040
rect 52400 62006 52434 62040
rect 52468 62006 52502 62040
rect 52536 62006 52570 62040
rect 52604 62006 52638 62040
rect 52672 62006 52706 62040
rect 52740 62006 52774 62040
rect 52808 62006 52842 62040
rect 52876 62006 52910 62040
rect 52944 62006 52978 62040
rect 53012 62006 53046 62040
rect 53080 62006 53114 62040
rect 53148 62006 53182 62040
rect 53216 62006 53250 62040
rect 53284 62006 53318 62040
rect 53352 62006 53386 62040
rect 53420 62006 53454 62040
rect 53488 62006 53522 62040
rect 53556 62006 53590 62040
rect 53624 62006 53658 62040
rect 53692 62006 53726 62040
rect 53760 62006 53794 62040
rect 53828 62006 53862 62040
rect 53896 62006 53930 62040
rect 53964 62006 53998 62040
rect 54032 62006 54066 62040
rect 54100 62006 54134 62040
rect 54168 62006 54202 62040
rect 54236 62006 54270 62040
rect 54304 62006 54338 62040
rect 54372 62006 54406 62040
rect 54440 62006 54474 62040
rect 54508 62006 54542 62040
rect 54576 62006 54610 62040
rect 54644 62006 54678 62040
rect 54712 62006 54746 62040
rect 54780 62006 54814 62040
rect 54848 62006 54882 62040
rect 54916 62006 54950 62040
rect 54984 62006 55018 62040
rect 55052 62006 55086 62040
rect 55120 62006 55154 62040
rect 55188 62006 55222 62040
rect 55256 62006 55290 62040
rect 55324 62006 55358 62040
rect 55392 62006 55426 62040
rect 55460 62006 55494 62040
rect 55528 62006 55562 62040
rect 55596 62006 55630 62040
rect 55664 62006 55698 62040
rect 55732 62006 55766 62040
rect 55800 62006 55834 62040
rect 55868 62006 55902 62040
rect 55936 62006 55970 62040
rect 56004 62006 56038 62040
rect 56072 62006 56106 62040
rect 56140 62006 56174 62040
rect 56208 62006 56242 62040
rect 56276 62006 56370 62040
rect 50436 61986 56370 62006
rect 50436 61976 50510 61986
rect 50436 61942 50456 61976
rect 50490 61942 50510 61976
rect 50436 61908 50510 61942
rect 50436 61874 50456 61908
rect 50490 61874 50510 61908
rect 50436 61840 50510 61874
rect 50436 61806 50456 61840
rect 50490 61806 50510 61840
rect 50436 61772 50510 61806
rect 50436 61738 50456 61772
rect 50490 61738 50510 61772
rect 50436 61704 50510 61738
rect 50436 61670 50456 61704
rect 50490 61670 50510 61704
rect 50436 61636 50510 61670
rect 50436 61602 50456 61636
rect 50490 61602 50510 61636
rect 50436 61568 50510 61602
rect 50436 61534 50456 61568
rect 50490 61534 50510 61568
rect 50436 61500 50510 61534
rect 50436 61466 50456 61500
rect 50490 61466 50510 61500
rect 50436 61432 50510 61466
rect 50436 61398 50456 61432
rect 50490 61398 50510 61432
rect 50436 61364 50510 61398
rect 50436 61330 50456 61364
rect 50490 61330 50510 61364
rect 50436 61296 50510 61330
rect 50436 61262 50456 61296
rect 50490 61262 50510 61296
rect 50436 61228 50510 61262
rect 50436 61194 50456 61228
rect 50490 61194 50510 61228
rect 50436 61160 50510 61194
rect 50436 61126 50456 61160
rect 50490 61126 50510 61160
rect 50436 61092 50510 61126
rect 50436 61058 50456 61092
rect 50490 61058 50510 61092
rect 50436 61024 50510 61058
rect 50436 60990 50456 61024
rect 50490 60990 50510 61024
rect 50436 60956 50510 60990
rect 50436 60922 50456 60956
rect 50490 60922 50510 60956
rect 50436 60888 50510 60922
rect 50436 60854 50456 60888
rect 50490 60854 50510 60888
rect 50436 60820 50510 60854
rect 50436 60786 50456 60820
rect 50490 60786 50510 60820
rect 50436 60752 50510 60786
rect 50436 60718 50456 60752
rect 50490 60718 50510 60752
rect 50436 60684 50510 60718
rect 50436 60650 50456 60684
rect 50490 60650 50510 60684
rect 50436 60616 50510 60650
rect 50436 60582 50456 60616
rect 50490 60582 50510 60616
rect 50436 60548 50510 60582
rect 50436 60514 50456 60548
rect 50490 60514 50510 60548
rect 50436 60480 50510 60514
rect 50436 60446 50456 60480
rect 50490 60446 50510 60480
rect 50436 60412 50510 60446
rect 50436 60378 50456 60412
rect 50490 60378 50510 60412
rect 50436 60344 50510 60378
rect 50436 60310 50456 60344
rect 50490 60310 50510 60344
rect 50436 60276 50510 60310
rect 50436 60242 50456 60276
rect 50490 60242 50510 60276
rect 50436 60208 50510 60242
rect 50436 60174 50456 60208
rect 50490 60174 50510 60208
rect 50436 60140 50510 60174
rect 50436 60106 50456 60140
rect 50490 60106 50510 60140
rect 50436 60072 50510 60106
rect 50436 60038 50456 60072
rect 50490 60038 50510 60072
rect 50436 60004 50510 60038
rect 50436 59970 50456 60004
rect 50490 59970 50510 60004
rect 50436 59936 50510 59970
rect 50436 59902 50456 59936
rect 50490 59902 50510 59936
rect 50436 59868 50510 59902
rect 50436 59834 50456 59868
rect 50490 59834 50510 59868
rect 50436 59800 50510 59834
rect 50436 59766 50456 59800
rect 50490 59766 50510 59800
rect 50436 59732 50510 59766
rect 50436 59698 50456 59732
rect 50490 59698 50510 59732
rect 50436 59664 50510 59698
rect 50436 59630 50456 59664
rect 50490 59630 50510 59664
rect 50436 59596 50510 59630
rect 50436 59562 50456 59596
rect 50490 59562 50510 59596
rect 50436 59528 50510 59562
rect 50436 59494 50456 59528
rect 50490 59494 50510 59528
rect 50436 59460 50510 59494
rect 50436 59426 50456 59460
rect 50490 59426 50510 59460
rect 50436 59392 50510 59426
rect 50436 59358 50456 59392
rect 50490 59358 50510 59392
rect 50436 59324 50510 59358
rect 50436 59290 50456 59324
rect 50490 59290 50510 59324
rect 50436 59256 50510 59290
rect 50436 59222 50456 59256
rect 50490 59222 50510 59256
rect 50436 59188 50510 59222
rect 50436 59154 50456 59188
rect 50490 59154 50510 59188
rect 50436 59120 50510 59154
rect 50436 59086 50456 59120
rect 50490 59086 50510 59120
rect 50436 59052 50510 59086
rect 50436 59018 50456 59052
rect 50490 59018 50510 59052
rect 50436 58984 50510 59018
rect 50436 58950 50456 58984
rect 50490 58950 50510 58984
rect 50436 58916 50510 58950
rect 50436 58882 50456 58916
rect 50490 58882 50510 58916
rect 50436 58848 50510 58882
rect 50436 58814 50456 58848
rect 50490 58814 50510 58848
rect 50436 58780 50510 58814
rect 50436 58746 50456 58780
rect 50490 58746 50510 58780
rect 50436 58712 50510 58746
rect 50436 58678 50456 58712
rect 50490 58678 50510 58712
rect 50436 58644 50510 58678
rect 50436 58610 50456 58644
rect 50490 58610 50510 58644
rect 50436 58576 50510 58610
rect 50436 58542 50456 58576
rect 50490 58542 50510 58576
rect 50436 58508 50510 58542
rect 50436 58474 50456 58508
rect 50490 58474 50510 58508
rect 50436 58440 50510 58474
rect 50436 58406 50456 58440
rect 50490 58406 50510 58440
rect 50436 58396 50510 58406
rect 56296 61976 56370 61986
rect 56296 61942 56316 61976
rect 56350 61942 56370 61976
rect 56296 61908 56370 61942
rect 56296 61874 56316 61908
rect 56350 61874 56370 61908
rect 56296 61840 56370 61874
rect 56296 61806 56316 61840
rect 56350 61806 56370 61840
rect 56296 61772 56370 61806
rect 56296 61738 56316 61772
rect 56350 61738 56370 61772
rect 56296 61704 56370 61738
rect 56296 61670 56316 61704
rect 56350 61670 56370 61704
rect 56296 61636 56370 61670
rect 56296 61602 56316 61636
rect 56350 61602 56370 61636
rect 56296 61568 56370 61602
rect 56296 61534 56316 61568
rect 56350 61534 56370 61568
rect 56296 61500 56370 61534
rect 56296 61466 56316 61500
rect 56350 61466 56370 61500
rect 56296 61432 56370 61466
rect 56296 61398 56316 61432
rect 56350 61398 56370 61432
rect 56296 61364 56370 61398
rect 56296 61330 56316 61364
rect 56350 61330 56370 61364
rect 56296 61296 56370 61330
rect 56296 61262 56316 61296
rect 56350 61262 56370 61296
rect 56296 61228 56370 61262
rect 56296 61194 56316 61228
rect 56350 61194 56370 61228
rect 56296 61160 56370 61194
rect 56296 61126 56316 61160
rect 56350 61126 56370 61160
rect 56296 61092 56370 61126
rect 56296 61058 56316 61092
rect 56350 61058 56370 61092
rect 56296 61024 56370 61058
rect 56296 60990 56316 61024
rect 56350 60990 56370 61024
rect 56296 60956 56370 60990
rect 56296 60922 56316 60956
rect 56350 60922 56370 60956
rect 56296 60888 56370 60922
rect 56296 60854 56316 60888
rect 56350 60854 56370 60888
rect 56296 60820 56370 60854
rect 56296 60786 56316 60820
rect 56350 60786 56370 60820
rect 56296 60752 56370 60786
rect 56296 60718 56316 60752
rect 56350 60718 56370 60752
rect 56296 60684 56370 60718
rect 56296 60650 56316 60684
rect 56350 60650 56370 60684
rect 56296 60616 56370 60650
rect 56296 60582 56316 60616
rect 56350 60582 56370 60616
rect 56296 60548 56370 60582
rect 56296 60514 56316 60548
rect 56350 60514 56370 60548
rect 56296 60480 56370 60514
rect 56296 60446 56316 60480
rect 56350 60446 56370 60480
rect 56296 60412 56370 60446
rect 56296 60378 56316 60412
rect 56350 60378 56370 60412
rect 56296 60344 56370 60378
rect 56296 60310 56316 60344
rect 56350 60310 56370 60344
rect 56296 60276 56370 60310
rect 56296 60242 56316 60276
rect 56350 60242 56370 60276
rect 56296 60208 56370 60242
rect 56296 60174 56316 60208
rect 56350 60174 56370 60208
rect 56296 60140 56370 60174
rect 56296 60106 56316 60140
rect 56350 60106 56370 60140
rect 56296 60072 56370 60106
rect 56296 60038 56316 60072
rect 56350 60038 56370 60072
rect 56296 60004 56370 60038
rect 56296 59970 56316 60004
rect 56350 59970 56370 60004
rect 56296 59936 56370 59970
rect 56296 59902 56316 59936
rect 56350 59902 56370 59936
rect 56296 59868 56370 59902
rect 56296 59834 56316 59868
rect 56350 59834 56370 59868
rect 56296 59800 56370 59834
rect 56296 59766 56316 59800
rect 56350 59766 56370 59800
rect 56296 59732 56370 59766
rect 56296 59698 56316 59732
rect 56350 59698 56370 59732
rect 56296 59664 56370 59698
rect 56296 59630 56316 59664
rect 56350 59630 56370 59664
rect 56296 59596 56370 59630
rect 56296 59562 56316 59596
rect 56350 59562 56370 59596
rect 56296 59528 56370 59562
rect 56296 59494 56316 59528
rect 56350 59494 56370 59528
rect 56296 59460 56370 59494
rect 56296 59426 56316 59460
rect 56350 59426 56370 59460
rect 56296 59392 56370 59426
rect 56296 59358 56316 59392
rect 56350 59358 56370 59392
rect 56296 59324 56370 59358
rect 56296 59290 56316 59324
rect 56350 59290 56370 59324
rect 56296 59256 56370 59290
rect 56296 59222 56316 59256
rect 56350 59222 56370 59256
rect 56296 59188 56370 59222
rect 56296 59154 56316 59188
rect 56350 59154 56370 59188
rect 56296 59120 56370 59154
rect 56296 59086 56316 59120
rect 56350 59086 56370 59120
rect 56296 59052 56370 59086
rect 56296 59018 56316 59052
rect 56350 59018 56370 59052
rect 56296 58984 56370 59018
rect 56296 58950 56316 58984
rect 56350 58950 56370 58984
rect 56296 58916 56370 58950
rect 56296 58882 56316 58916
rect 56350 58882 56370 58916
rect 56296 58848 56370 58882
rect 56296 58814 56316 58848
rect 56350 58814 56370 58848
rect 56296 58780 56370 58814
rect 56296 58746 56316 58780
rect 56350 58746 56370 58780
rect 56296 58712 56370 58746
rect 56296 58678 56316 58712
rect 56350 58678 56370 58712
rect 56296 58644 56370 58678
rect 56296 58610 56316 58644
rect 56350 58610 56370 58644
rect 56296 58576 56370 58610
rect 56296 58542 56316 58576
rect 56350 58542 56370 58576
rect 56296 58508 56370 58542
rect 56296 58474 56316 58508
rect 56350 58474 56370 58508
rect 56296 58440 56370 58474
rect 56296 58406 56316 58440
rect 56350 58406 56370 58440
rect 56296 58396 56370 58406
rect 50436 58376 56370 58396
rect 50436 58342 50530 58376
rect 50564 58342 50598 58376
rect 50632 58342 50666 58376
rect 50700 58342 50734 58376
rect 50768 58342 50802 58376
rect 50836 58342 50870 58376
rect 50904 58342 50938 58376
rect 50972 58342 51006 58376
rect 51040 58342 51074 58376
rect 51108 58342 51142 58376
rect 51176 58342 51210 58376
rect 51244 58342 51278 58376
rect 51312 58342 51346 58376
rect 51380 58342 51414 58376
rect 51448 58342 51482 58376
rect 51516 58342 51550 58376
rect 51584 58342 51618 58376
rect 51652 58342 51686 58376
rect 51720 58342 51754 58376
rect 51788 58342 51822 58376
rect 51856 58342 51890 58376
rect 51924 58342 51958 58376
rect 51992 58342 52026 58376
rect 52060 58342 52094 58376
rect 52128 58342 52162 58376
rect 52196 58342 52230 58376
rect 52264 58342 52298 58376
rect 52332 58342 52366 58376
rect 52400 58342 52434 58376
rect 52468 58342 52502 58376
rect 52536 58342 52570 58376
rect 52604 58342 52638 58376
rect 52672 58342 52706 58376
rect 52740 58342 52774 58376
rect 52808 58342 52842 58376
rect 52876 58342 52910 58376
rect 52944 58342 52978 58376
rect 53012 58342 53046 58376
rect 53080 58342 53114 58376
rect 53148 58342 53182 58376
rect 53216 58342 53250 58376
rect 53284 58342 53318 58376
rect 53352 58342 53386 58376
rect 53420 58342 53454 58376
rect 53488 58342 53522 58376
rect 53556 58342 53590 58376
rect 53624 58342 53658 58376
rect 53692 58342 53726 58376
rect 53760 58342 53794 58376
rect 53828 58342 53862 58376
rect 53896 58342 53930 58376
rect 53964 58342 53998 58376
rect 54032 58342 54066 58376
rect 54100 58342 54134 58376
rect 54168 58342 54202 58376
rect 54236 58342 54270 58376
rect 54304 58342 54338 58376
rect 54372 58342 54406 58376
rect 54440 58342 54474 58376
rect 54508 58342 54542 58376
rect 54576 58342 54610 58376
rect 54644 58342 54678 58376
rect 54712 58342 54746 58376
rect 54780 58342 54814 58376
rect 54848 58342 54882 58376
rect 54916 58342 54950 58376
rect 54984 58342 55018 58376
rect 55052 58342 55086 58376
rect 55120 58342 55154 58376
rect 55188 58342 55222 58376
rect 55256 58342 55290 58376
rect 55324 58342 55358 58376
rect 55392 58342 55426 58376
rect 55460 58342 55494 58376
rect 55528 58342 55562 58376
rect 55596 58342 55630 58376
rect 55664 58342 55698 58376
rect 55732 58342 55766 58376
rect 55800 58342 55834 58376
rect 55868 58342 55902 58376
rect 55936 58342 55970 58376
rect 56004 58342 56038 58376
rect 56072 58342 56106 58376
rect 56140 58342 56174 58376
rect 56208 58342 56242 58376
rect 56276 58342 56370 58376
rect 50436 58322 56370 58342
rect 59084 62029 59158 62063
rect 59084 61995 59104 62029
rect 59138 61995 59158 62029
rect 59084 61961 59158 61995
rect 59084 61927 59104 61961
rect 59138 61927 59158 61961
rect 59084 61893 59158 61927
rect 59084 61859 59104 61893
rect 59138 61859 59158 61893
rect 59084 61825 59158 61859
rect 59084 61791 59104 61825
rect 59138 61791 59158 61825
rect 59084 61757 59158 61791
rect 59084 61723 59104 61757
rect 59138 61723 59158 61757
rect 59084 61689 59158 61723
rect 59084 61655 59104 61689
rect 59138 61655 59158 61689
rect 59084 61621 59158 61655
rect 59084 61587 59104 61621
rect 59138 61587 59158 61621
rect 59084 61553 59158 61587
rect 59084 61519 59104 61553
rect 59138 61519 59158 61553
rect 59084 61485 59158 61519
rect 59084 61451 59104 61485
rect 59138 61451 59158 61485
rect 59084 61417 59158 61451
rect 59084 61383 59104 61417
rect 59138 61383 59158 61417
rect 59084 61349 59158 61383
rect 59084 61315 59104 61349
rect 59138 61315 59158 61349
rect 59084 61281 59158 61315
rect 59084 61247 59104 61281
rect 59138 61247 59158 61281
rect 59084 61213 59158 61247
rect 59084 61179 59104 61213
rect 59138 61179 59158 61213
rect 59084 61145 59158 61179
rect 59084 61111 59104 61145
rect 59138 61111 59158 61145
rect 59084 61077 59158 61111
rect 59084 61043 59104 61077
rect 59138 61043 59158 61077
rect 59084 61009 59158 61043
rect 59084 60975 59104 61009
rect 59138 60975 59158 61009
rect 59084 60941 59158 60975
rect 59084 60907 59104 60941
rect 59138 60907 59158 60941
rect 59084 60873 59158 60907
rect 59084 60839 59104 60873
rect 59138 60839 59158 60873
rect 59084 60805 59158 60839
rect 59084 60771 59104 60805
rect 59138 60771 59158 60805
rect 59084 60737 59158 60771
rect 59084 60703 59104 60737
rect 59138 60703 59158 60737
rect 59084 60669 59158 60703
rect 59084 60635 59104 60669
rect 59138 60635 59158 60669
rect 59084 60601 59158 60635
rect 59084 60567 59104 60601
rect 59138 60567 59158 60601
rect 59084 60533 59158 60567
rect 59084 60499 59104 60533
rect 59138 60499 59158 60533
rect 59084 60465 59158 60499
rect 59084 60431 59104 60465
rect 59138 60431 59158 60465
rect 59084 60397 59158 60431
rect 59084 60363 59104 60397
rect 59138 60363 59158 60397
rect 59084 60329 59158 60363
rect 59084 60295 59104 60329
rect 59138 60295 59158 60329
rect 59084 60261 59158 60295
rect 59084 60227 59104 60261
rect 59138 60227 59158 60261
rect 59084 60193 59158 60227
rect 59084 60159 59104 60193
rect 59138 60159 59158 60193
rect 59084 60125 59158 60159
rect 59084 60091 59104 60125
rect 59138 60091 59158 60125
rect 59084 60057 59158 60091
rect 59084 60023 59104 60057
rect 59138 60023 59158 60057
rect 59084 59989 59158 60023
rect 59084 59955 59104 59989
rect 59138 59955 59158 59989
rect 59084 59921 59158 59955
rect 59084 59887 59104 59921
rect 59138 59887 59158 59921
rect 59084 59853 59158 59887
rect 59084 59819 59104 59853
rect 59138 59819 59158 59853
rect 59084 59785 59158 59819
rect 59084 59751 59104 59785
rect 59138 59751 59158 59785
rect 59084 59717 59158 59751
rect 59084 59683 59104 59717
rect 59138 59683 59158 59717
rect 59084 59649 59158 59683
rect 59084 59615 59104 59649
rect 59138 59615 59158 59649
rect 59084 59581 59158 59615
rect 59084 59547 59104 59581
rect 59138 59547 59158 59581
rect 59084 59513 59158 59547
rect 59084 59479 59104 59513
rect 59138 59479 59158 59513
rect 59084 59445 59158 59479
rect 59084 59411 59104 59445
rect 59138 59411 59158 59445
rect 59084 59377 59158 59411
rect 59084 59343 59104 59377
rect 59138 59343 59158 59377
rect 59084 59309 59158 59343
rect 59084 59275 59104 59309
rect 59138 59275 59158 59309
rect 59084 59241 59158 59275
rect 59084 59207 59104 59241
rect 59138 59207 59158 59241
rect 59084 59173 59158 59207
rect 59084 59139 59104 59173
rect 59138 59139 59158 59173
rect 59084 59105 59158 59139
rect 59084 59071 59104 59105
rect 59138 59071 59158 59105
rect 59084 59037 59158 59071
rect 59084 59003 59104 59037
rect 59138 59003 59158 59037
rect 59084 58969 59158 59003
rect 59084 58935 59104 58969
rect 59138 58935 59158 58969
rect 59084 58901 59158 58935
rect 59084 58867 59104 58901
rect 59138 58867 59158 58901
rect 59084 58833 59158 58867
rect 59084 58799 59104 58833
rect 59138 58799 59158 58833
rect 59084 58765 59158 58799
rect 59084 58731 59104 58765
rect 59138 58731 59158 58765
rect 59084 58697 59158 58731
rect 59084 58663 59104 58697
rect 59138 58663 59158 58697
rect 59084 58629 59158 58663
rect 59084 58595 59104 58629
rect 59138 58595 59158 58629
rect 59084 58561 59158 58595
rect 59084 58527 59104 58561
rect 59138 58527 59158 58561
rect 59084 58493 59158 58527
rect 59084 58459 59104 58493
rect 59138 58459 59158 58493
rect 59084 58425 59158 58459
rect 59084 58391 59104 58425
rect 59138 58391 59158 58425
rect 59084 58357 59158 58391
rect 59084 58323 59104 58357
rect 59138 58323 59158 58357
rect -3738 58274 -3718 58308
rect -3684 58274 -3664 58308
rect -3738 58240 -3664 58274
rect -3738 58206 -3718 58240
rect -3684 58206 -3664 58240
rect -3738 58172 -3664 58206
rect -3738 58138 -3718 58172
rect -3684 58138 -3664 58172
rect -3738 58104 -3664 58138
rect -3738 58070 -3718 58104
rect -3684 58070 -3664 58104
rect -3738 58036 -3664 58070
rect -3738 58002 -3718 58036
rect -3684 58002 -3664 58036
rect -3738 57968 -3664 58002
rect -3738 57934 -3718 57968
rect -3684 57934 -3664 57968
rect -3738 57900 -3664 57934
rect -3738 57866 -3718 57900
rect -3684 57866 -3664 57900
rect -3738 57832 -3664 57866
rect -3738 57798 -3718 57832
rect -3684 57798 -3664 57832
rect -3738 57764 -3664 57798
rect -3738 57730 -3718 57764
rect -3684 57730 -3664 57764
rect -3738 57696 -3664 57730
rect -3738 57662 -3718 57696
rect -3684 57662 -3664 57696
rect -3738 57628 -3664 57662
rect -3738 57594 -3718 57628
rect -3684 57594 -3664 57628
rect -3738 57560 -3664 57594
rect -3738 57526 -3718 57560
rect -3684 57526 -3664 57560
rect -3738 57492 -3664 57526
rect -3738 57458 -3718 57492
rect -3684 57458 -3664 57492
rect -3738 57424 -3664 57458
rect -3738 57390 -3718 57424
rect -3684 57390 -3664 57424
rect -3738 57356 -3664 57390
rect -3738 57322 -3718 57356
rect -3684 57322 -3664 57356
rect -3738 57288 -3664 57322
rect -3738 57254 -3718 57288
rect -3684 57254 -3664 57288
rect -3738 57220 -3664 57254
rect -3738 57186 -3718 57220
rect -3684 57186 -3664 57220
rect -3738 57152 -3664 57186
rect -3738 57118 -3718 57152
rect -3684 57118 -3664 57152
rect -3738 57084 -3664 57118
rect -3738 57050 -3718 57084
rect -3684 57050 -3664 57084
rect -3738 57016 -3664 57050
rect -3738 56982 -3718 57016
rect -3684 56982 -3664 57016
rect -3738 56948 -3664 56982
rect -3738 56914 -3718 56948
rect -3684 56914 -3664 56948
rect -3738 56880 -3664 56914
rect -3738 56846 -3718 56880
rect -3684 56846 -3664 56880
rect -3738 56812 -3664 56846
rect -3738 56778 -3718 56812
rect -3684 56778 -3664 56812
rect -3738 56744 -3664 56778
rect -3738 56710 -3718 56744
rect -3684 56710 -3664 56744
rect -3738 56676 -3664 56710
rect -3738 56642 -3718 56676
rect -3684 56642 -3664 56676
rect -3738 56608 -3664 56642
rect -3738 56574 -3718 56608
rect -3684 56574 -3664 56608
rect -3738 56540 -3664 56574
rect -3738 56506 -3718 56540
rect -3684 56506 -3664 56540
rect -3738 56472 -3664 56506
rect -3738 56438 -3718 56472
rect -3684 56438 -3664 56472
rect -3738 56404 -3664 56438
rect -3738 56370 -3718 56404
rect -3684 56370 -3664 56404
rect -3738 56336 -3664 56370
rect -3738 56302 -3718 56336
rect -3684 56302 -3664 56336
rect -3738 56268 -3664 56302
rect -10719 56245 -10645 56250
rect -10719 56211 -10699 56245
rect -10665 56211 -10645 56245
rect -10719 56177 -10645 56211
rect -10719 56143 -10699 56177
rect -10665 56143 -10645 56177
rect -10719 56109 -10645 56143
rect -10719 56075 -10699 56109
rect -10665 56075 -10645 56109
rect -10719 56041 -10645 56075
rect -10719 56007 -10699 56041
rect -10665 56007 -10645 56041
rect -10719 55973 -10645 56007
rect -10719 55939 -10699 55973
rect -10665 55939 -10645 55973
rect -10719 55905 -10645 55939
rect -10719 55871 -10699 55905
rect -10665 55871 -10645 55905
rect -10719 55837 -10645 55871
rect -10719 55803 -10699 55837
rect -10665 55803 -10645 55837
rect -10719 55769 -10645 55803
rect -10719 55735 -10699 55769
rect -10665 55735 -10645 55769
rect -10719 55701 -10645 55735
rect -10719 55667 -10699 55701
rect -10665 55667 -10645 55701
rect -10719 55633 -10645 55667
rect -10719 55599 -10699 55633
rect -10665 55599 -10645 55633
rect -10719 55565 -10645 55599
rect -10719 55531 -10699 55565
rect -10665 55531 -10645 55565
rect -10719 55497 -10645 55531
rect -10719 55463 -10699 55497
rect -10665 55463 -10645 55497
rect -10719 55429 -10645 55463
rect -10719 55395 -10699 55429
rect -10665 55395 -10645 55429
rect -10719 55361 -10645 55395
rect -10719 55327 -10699 55361
rect -10665 55327 -10645 55361
rect -10719 55293 -10645 55327
rect -10719 55259 -10699 55293
rect -10665 55259 -10645 55293
rect -10719 55225 -10645 55259
rect -10719 55191 -10699 55225
rect -10665 55191 -10645 55225
rect -10719 55157 -10645 55191
rect -10719 55123 -10699 55157
rect -10665 55123 -10645 55157
rect -10719 55089 -10645 55123
rect -10719 55055 -10699 55089
rect -10665 55055 -10645 55089
rect -10719 55021 -10645 55055
rect -10719 54987 -10699 55021
rect -10665 54987 -10645 55021
rect -10719 54953 -10645 54987
rect -10719 54919 -10699 54953
rect -10665 54919 -10645 54953
rect -10719 54885 -10645 54919
rect -10719 54851 -10699 54885
rect -10665 54851 -10645 54885
rect -10719 54817 -10645 54851
rect -10719 54783 -10699 54817
rect -10665 54783 -10645 54817
rect -10719 54749 -10645 54783
rect -10719 54715 -10699 54749
rect -10665 54715 -10645 54749
rect -10719 54681 -10645 54715
rect -10719 54647 -10699 54681
rect -10665 54647 -10645 54681
rect -10719 54613 -10645 54647
rect -10719 54579 -10699 54613
rect -10665 54579 -10645 54613
rect -10719 54545 -10645 54579
rect -10719 54511 -10699 54545
rect -10665 54511 -10645 54545
rect -10719 54477 -10645 54511
rect -10719 54443 -10699 54477
rect -10665 54443 -10645 54477
rect -10719 54409 -10645 54443
rect -10719 54375 -10699 54409
rect -10665 54375 -10645 54409
rect -10719 54341 -10645 54375
rect -10719 54307 -10699 54341
rect -10665 54307 -10645 54341
rect -10719 54273 -10645 54307
rect -10719 54239 -10699 54273
rect -10665 54239 -10645 54273
rect -10719 54205 -10645 54239
rect -10719 54171 -10699 54205
rect -10665 54171 -10645 54205
rect -10719 54137 -10645 54171
rect -10719 54103 -10699 54137
rect -10665 54103 -10645 54137
rect -10719 54069 -10645 54103
rect -10719 54035 -10699 54069
rect -10665 54035 -10645 54069
rect -10719 54001 -10645 54035
rect -10719 53967 -10699 54001
rect -10665 53967 -10645 54001
rect -10719 53933 -10645 53967
rect -10719 53899 -10699 53933
rect -10665 53899 -10645 53933
rect -10719 53865 -10645 53899
rect -10719 53831 -10699 53865
rect -10665 53831 -10645 53865
rect -10719 53797 -10645 53831
rect -10719 53763 -10699 53797
rect -10665 53763 -10645 53797
rect -10719 53729 -10645 53763
rect -10719 53695 -10699 53729
rect -10665 53695 -10645 53729
rect -10719 53661 -10645 53695
rect -10719 53627 -10699 53661
rect -10665 53627 -10645 53661
rect -10719 53593 -10645 53627
rect -10719 53559 -10699 53593
rect -10665 53559 -10645 53593
rect -10719 53525 -10645 53559
rect -10719 53491 -10699 53525
rect -10665 53491 -10645 53525
rect -10719 53457 -10645 53491
rect -10719 53423 -10699 53457
rect -10665 53423 -10645 53457
rect -10719 53389 -10645 53423
rect -10719 53355 -10699 53389
rect -10665 53355 -10645 53389
rect -10719 53321 -10645 53355
rect -10719 53287 -10699 53321
rect -10665 53287 -10645 53321
rect -10719 53253 -10645 53287
rect -10719 53219 -10699 53253
rect -10665 53219 -10645 53253
rect -10719 53185 -10645 53219
rect -10719 53151 -10699 53185
rect -10665 53151 -10645 53185
rect -10719 53117 -10645 53151
rect -10719 53083 -10699 53117
rect -10665 53083 -10645 53117
rect -10719 53049 -10645 53083
rect -10719 53015 -10699 53049
rect -10665 53015 -10645 53049
rect -10719 52981 -10645 53015
rect -10719 52947 -10699 52981
rect -10665 52947 -10645 52981
rect -10719 52913 -10645 52947
rect -10719 52879 -10699 52913
rect -10665 52879 -10645 52913
rect -10719 52845 -10645 52879
rect -10719 52811 -10699 52845
rect -10665 52811 -10645 52845
rect -10719 52777 -10645 52811
rect -10719 52743 -10699 52777
rect -10665 52743 -10645 52777
rect -10719 52709 -10645 52743
rect -10719 52675 -10699 52709
rect -10665 52675 -10645 52709
rect -10719 52641 -10645 52675
rect -10719 52607 -10699 52641
rect -10665 52607 -10645 52641
rect -10719 52573 -10645 52607
rect -10719 52539 -10699 52573
rect -10665 52539 -10645 52573
rect -10719 52505 -10645 52539
rect -10719 52471 -10699 52505
rect -10665 52471 -10645 52505
rect -10719 52437 -10645 52471
rect -10719 52403 -10699 52437
rect -10665 52403 -10645 52437
rect -10719 52369 -10645 52403
rect -10719 52335 -10699 52369
rect -10665 52335 -10645 52369
rect -10719 52301 -10645 52335
rect -10719 52267 -10699 52301
rect -10665 52267 -10645 52301
rect -10719 52233 -10645 52267
rect -10719 52199 -10699 52233
rect -10665 52199 -10645 52233
rect -10719 52165 -10645 52199
rect -10719 52131 -10699 52165
rect -10665 52131 -10645 52165
rect -10719 52097 -10645 52131
rect -10719 52063 -10699 52097
rect -10665 52063 -10645 52097
rect -10719 52029 -10645 52063
rect -10719 51995 -10699 52029
rect -10665 51995 -10645 52029
rect -10719 51961 -10645 51995
rect -10719 51927 -10699 51961
rect -10665 51927 -10645 51961
rect -10719 51893 -10645 51927
rect -10719 51859 -10699 51893
rect -10665 51859 -10645 51893
rect -10719 51825 -10645 51859
rect -10719 51791 -10699 51825
rect -10665 51791 -10645 51825
rect -10719 51757 -10645 51791
rect -10719 51723 -10699 51757
rect -10665 51723 -10645 51757
rect -10719 51689 -10645 51723
rect -10719 51655 -10699 51689
rect -10665 51655 -10645 51689
rect -10719 51621 -10645 51655
rect -10719 51587 -10699 51621
rect -10665 51587 -10645 51621
rect -10719 51553 -10645 51587
rect -10719 51519 -10699 51553
rect -10665 51519 -10645 51553
rect -10719 51485 -10645 51519
rect -10719 51451 -10699 51485
rect -10665 51451 -10645 51485
rect -10719 51417 -10645 51451
rect -10719 51383 -10699 51417
rect -10665 51383 -10645 51417
rect -10719 51349 -10645 51383
rect -10719 51315 -10699 51349
rect -10665 51315 -10645 51349
rect -10719 51281 -10645 51315
rect -10719 51247 -10699 51281
rect -10665 51247 -10645 51281
rect -10719 51213 -10645 51247
rect -10719 51179 -10699 51213
rect -10665 51179 -10645 51213
rect -10719 51145 -10645 51179
rect -10719 51111 -10699 51145
rect -10665 51111 -10645 51145
rect -10719 51077 -10645 51111
rect -10719 51043 -10699 51077
rect -10665 51043 -10645 51077
rect -10719 51009 -10645 51043
rect -10719 50975 -10699 51009
rect -10665 50975 -10645 51009
rect -10719 50941 -10645 50975
rect -10719 50907 -10699 50941
rect -10665 50907 -10645 50941
rect -10719 50873 -10645 50907
rect -10719 50839 -10699 50873
rect -10665 50839 -10645 50873
rect -10719 50805 -10645 50839
rect -10719 50771 -10699 50805
rect -10665 50771 -10645 50805
rect -10719 50737 -10645 50771
rect -10719 50703 -10699 50737
rect -10665 50703 -10645 50737
rect -10719 50669 -10645 50703
rect -10719 50635 -10699 50669
rect -10665 50635 -10645 50669
rect -10719 50601 -10645 50635
rect -10719 50567 -10699 50601
rect -10665 50567 -10645 50601
rect -10719 50533 -10645 50567
rect -10719 50499 -10699 50533
rect -10665 50499 -10645 50533
rect -10719 50465 -10645 50499
rect -10719 50431 -10699 50465
rect -10665 50431 -10645 50465
rect -10719 50397 -10645 50431
rect -10719 50363 -10699 50397
rect -10665 50363 -10645 50397
rect -10719 50329 -10645 50363
rect -10719 50295 -10699 50329
rect -10665 50295 -10645 50329
rect -10719 50261 -10645 50295
rect -10719 50227 -10699 50261
rect -10665 50227 -10645 50261
rect -10719 50193 -10645 50227
rect -10719 50159 -10699 50193
rect -10665 50159 -10645 50193
rect -10719 50125 -10645 50159
rect -10719 50091 -10699 50125
rect -10665 50091 -10645 50125
rect -10719 50057 -10645 50091
rect -10719 50023 -10699 50057
rect -10665 50023 -10645 50057
rect -10719 49989 -10645 50023
rect -10719 49955 -10699 49989
rect -10665 49955 -10645 49989
rect -10719 49921 -10645 49955
rect -10719 49887 -10699 49921
rect -10665 49887 -10645 49921
rect -10719 49853 -10645 49887
rect -10719 49819 -10699 49853
rect -10665 49819 -10645 49853
rect -10719 49785 -10645 49819
rect -10719 49751 -10699 49785
rect -10665 49751 -10645 49785
rect -10719 49717 -10645 49751
rect -10719 49683 -10699 49717
rect -10665 49683 -10645 49717
rect -10719 49649 -10645 49683
rect -10719 49615 -10699 49649
rect -10665 49615 -10645 49649
rect -10719 49581 -10645 49615
rect -10719 49547 -10699 49581
rect -10665 49547 -10645 49581
rect -10719 49513 -10645 49547
rect -10719 49479 -10699 49513
rect -10665 49479 -10645 49513
rect -10719 49445 -10645 49479
rect -10719 49411 -10699 49445
rect -10665 49411 -10645 49445
rect -10719 49377 -10645 49411
rect -10719 49343 -10699 49377
rect -10665 49343 -10645 49377
rect -10719 49309 -10645 49343
rect -10719 49275 -10699 49309
rect -10665 49275 -10645 49309
rect -10719 49241 -10645 49275
rect -10719 49207 -10699 49241
rect -10665 49207 -10645 49241
rect -10719 49173 -10645 49207
rect -10719 49139 -10699 49173
rect -10665 49139 -10645 49173
rect -10719 49105 -10645 49139
rect -10719 49071 -10699 49105
rect -10665 49071 -10645 49105
rect -10719 49037 -10645 49071
rect -10719 49003 -10699 49037
rect -10665 49003 -10645 49037
rect -10719 48969 -10645 49003
rect -10719 48935 -10699 48969
rect -10665 48935 -10645 48969
rect -10719 48901 -10645 48935
rect -10719 48867 -10699 48901
rect -10665 48867 -10645 48901
rect -10719 48833 -10645 48867
rect -10719 48799 -10699 48833
rect -10665 48799 -10645 48833
rect -10719 48765 -10645 48799
rect -10719 48731 -10699 48765
rect -10665 48731 -10645 48765
rect -10719 48697 -10645 48731
rect -10719 48663 -10699 48697
rect -10665 48663 -10645 48697
rect -10719 48629 -10645 48663
rect -10719 48595 -10699 48629
rect -10665 48595 -10645 48629
rect -10719 48561 -10645 48595
rect -10719 48527 -10699 48561
rect -10665 48527 -10645 48561
rect -10719 48493 -10645 48527
rect -10719 48459 -10699 48493
rect -10665 48459 -10645 48493
rect -10719 48425 -10645 48459
rect -10719 48391 -10699 48425
rect -10665 48391 -10645 48425
rect -10719 48357 -10645 48391
rect -10719 48323 -10699 48357
rect -10665 48323 -10645 48357
rect -10719 48289 -10645 48323
rect -10719 48255 -10699 48289
rect -10665 48255 -10645 48289
rect -10719 48221 -10645 48255
rect -10719 48187 -10699 48221
rect -10665 48187 -10645 48221
rect -10719 48153 -10645 48187
rect -10719 48119 -10699 48153
rect -10665 48119 -10645 48153
rect -10719 48085 -10645 48119
rect -10719 48051 -10699 48085
rect -10665 48051 -10645 48085
rect -10719 48017 -10645 48051
rect -10719 47983 -10699 48017
rect -10665 47983 -10645 48017
rect -10719 47949 -10645 47983
rect -10719 47915 -10699 47949
rect -10665 47915 -10645 47949
rect -10719 47881 -10645 47915
rect -10719 47847 -10699 47881
rect -10665 47847 -10645 47881
rect -10719 47813 -10645 47847
rect -10719 47779 -10699 47813
rect -10665 47779 -10645 47813
rect -10719 47745 -10645 47779
rect -10719 47711 -10699 47745
rect -10665 47711 -10645 47745
rect -10719 47677 -10645 47711
rect -10719 47643 -10699 47677
rect -10665 47643 -10645 47677
rect -10719 47609 -10645 47643
rect -10719 47575 -10699 47609
rect -10665 47575 -10645 47609
rect -10719 47541 -10645 47575
rect -10719 47507 -10699 47541
rect -10665 47507 -10645 47541
rect -10719 47473 -10645 47507
rect -10719 47439 -10699 47473
rect -10665 47439 -10645 47473
rect -10719 47405 -10645 47439
rect -10719 47371 -10699 47405
rect -10665 47371 -10645 47405
rect -10719 47337 -10645 47371
rect -10719 47303 -10699 47337
rect -10665 47303 -10645 47337
rect -10719 47269 -10645 47303
rect -10719 47235 -10699 47269
rect -10665 47235 -10645 47269
rect -10719 47201 -10645 47235
rect -10719 47167 -10699 47201
rect -10665 47167 -10645 47201
rect -10719 47133 -10645 47167
rect -10719 47099 -10699 47133
rect -10665 47099 -10645 47133
rect -10719 47065 -10645 47099
rect -10719 47031 -10699 47065
rect -10665 47031 -10645 47065
rect -10719 46997 -10645 47031
rect -10719 46963 -10699 46997
rect -10665 46963 -10645 46997
rect -10719 46929 -10645 46963
rect -10719 46895 -10699 46929
rect -10665 46895 -10645 46929
rect -10719 46861 -10645 46895
rect -10719 46827 -10699 46861
rect -10665 46827 -10645 46861
rect -10719 46793 -10645 46827
rect -10719 46759 -10699 46793
rect -10665 46759 -10645 46793
rect -10719 46725 -10645 46759
rect -10719 46691 -10699 46725
rect -10665 46691 -10645 46725
rect -10719 46657 -10645 46691
rect -10719 46623 -10699 46657
rect -10665 46623 -10645 46657
rect -10719 46589 -10645 46623
rect -10719 46555 -10699 46589
rect -10665 46555 -10645 46589
rect -10719 46521 -10645 46555
rect -10719 46487 -10699 46521
rect -10665 46487 -10645 46521
rect -10719 46453 -10645 46487
rect -10719 46419 -10699 46453
rect -10665 46419 -10645 46453
rect -10719 46385 -10645 46419
rect -10719 46351 -10699 46385
rect -10665 46351 -10645 46385
rect -10719 46317 -10645 46351
rect -10719 46283 -10699 46317
rect -10665 46283 -10645 46317
rect -10719 46249 -10645 46283
rect -10719 46215 -10699 46249
rect -10665 46215 -10645 46249
rect -10719 46181 -10645 46215
rect -10719 46147 -10699 46181
rect -10665 46147 -10645 46181
rect -10719 46113 -10645 46147
rect -10719 46079 -10699 46113
rect -10665 46079 -10645 46113
rect -10719 46045 -10645 46079
rect -10719 46011 -10699 46045
rect -10665 46011 -10645 46045
rect -10719 45977 -10645 46011
rect -10719 45943 -10699 45977
rect -10665 45943 -10645 45977
rect -10719 45909 -10645 45943
rect -10719 45875 -10699 45909
rect -10665 45875 -10645 45909
rect -10719 45841 -10645 45875
rect -10719 45807 -10699 45841
rect -10665 45807 -10645 45841
rect -10719 45773 -10645 45807
rect -10719 45739 -10699 45773
rect -10665 45739 -10645 45773
rect -10719 45705 -10645 45739
rect -10719 45671 -10699 45705
rect -10665 45671 -10645 45705
rect -10719 45637 -10645 45671
rect -10719 45603 -10699 45637
rect -10665 45603 -10645 45637
rect -10719 45569 -10645 45603
rect -10719 45535 -10699 45569
rect -10665 45535 -10645 45569
rect -10719 45501 -10645 45535
rect -10719 45467 -10699 45501
rect -10665 45467 -10645 45501
rect -10719 45433 -10645 45467
rect -10719 45399 -10699 45433
rect -10665 45399 -10645 45433
rect -10719 45365 -10645 45399
rect -10719 45331 -10699 45365
rect -10665 45331 -10645 45365
rect -10719 45297 -10645 45331
rect -10719 45263 -10699 45297
rect -10665 45263 -10645 45297
rect -10719 45229 -10645 45263
rect -10719 45195 -10699 45229
rect -10665 45195 -10645 45229
rect -10719 45161 -10645 45195
rect -10719 45127 -10699 45161
rect -10665 45127 -10645 45161
rect -10719 45093 -10645 45127
rect -10719 45059 -10699 45093
rect -10665 45059 -10645 45093
rect -10719 45025 -10645 45059
rect -10719 44991 -10699 45025
rect -10665 44991 -10645 45025
rect -10719 44957 -10645 44991
rect -10719 44923 -10699 44957
rect -10665 44923 -10645 44957
rect -10719 44889 -10645 44923
rect -10719 44855 -10699 44889
rect -10665 44855 -10645 44889
rect -10719 44821 -10645 44855
rect -10719 44787 -10699 44821
rect -10665 44787 -10645 44821
rect -10719 44753 -10645 44787
rect -10719 44719 -10699 44753
rect -10665 44719 -10645 44753
rect -10719 44685 -10645 44719
rect -10719 44651 -10699 44685
rect -10665 44651 -10645 44685
rect -10719 44617 -10645 44651
rect -10719 44583 -10699 44617
rect -10665 44583 -10645 44617
rect -10719 44549 -10645 44583
rect -10719 44515 -10699 44549
rect -10665 44515 -10645 44549
rect -10719 44481 -10645 44515
rect -10719 44447 -10699 44481
rect -10665 44447 -10645 44481
rect -10719 44413 -10645 44447
rect -10719 44379 -10699 44413
rect -10665 44379 -10645 44413
rect -10719 44345 -10645 44379
rect -10719 44311 -10699 44345
rect -10665 44311 -10645 44345
rect -10719 44300 -10645 44311
rect -3738 56234 -3718 56268
rect -3684 56234 -3664 56268
rect -3738 56200 -3664 56234
rect -3738 56166 -3718 56200
rect -3684 56166 -3664 56200
rect -3738 56132 -3664 56166
rect -3738 56098 -3718 56132
rect -3684 56098 -3664 56132
rect -3738 56064 -3664 56098
rect -3738 56030 -3718 56064
rect -3684 56030 -3664 56064
rect -3738 55996 -3664 56030
rect -3738 55962 -3718 55996
rect -3684 55962 -3664 55996
rect -3738 55928 -3664 55962
rect -3738 55894 -3718 55928
rect -3684 55894 -3664 55928
rect -3738 55860 -3664 55894
rect -3738 55826 -3718 55860
rect -3684 55826 -3664 55860
rect -3738 55792 -3664 55826
rect -3738 55758 -3718 55792
rect -3684 55758 -3664 55792
rect -3738 55724 -3664 55758
rect -3738 55690 -3718 55724
rect -3684 55690 -3664 55724
rect -3738 55656 -3664 55690
rect -3738 55622 -3718 55656
rect -3684 55622 -3664 55656
rect -3738 55588 -3664 55622
rect -3738 55554 -3718 55588
rect -3684 55554 -3664 55588
rect -3738 55520 -3664 55554
rect -3738 55486 -3718 55520
rect -3684 55486 -3664 55520
rect -3738 55452 -3664 55486
rect -3738 55418 -3718 55452
rect -3684 55418 -3664 55452
rect -3738 55384 -3664 55418
rect -3738 55350 -3718 55384
rect -3684 55350 -3664 55384
rect -3738 55316 -3664 55350
rect -3738 55282 -3718 55316
rect -3684 55282 -3664 55316
rect -3738 55248 -3664 55282
rect -3738 55214 -3718 55248
rect -3684 55214 -3664 55248
rect -3738 55180 -3664 55214
rect -3738 55146 -3718 55180
rect -3684 55146 -3664 55180
rect -3738 55112 -3664 55146
rect -3738 55078 -3718 55112
rect -3684 55078 -3664 55112
rect -3738 55044 -3664 55078
rect -3738 55010 -3718 55044
rect -3684 55010 -3664 55044
rect -3738 54976 -3664 55010
rect -3738 54942 -3718 54976
rect -3684 54942 -3664 54976
rect -3738 54908 -3664 54942
rect -3738 54874 -3718 54908
rect -3684 54874 -3664 54908
rect -3738 54840 -3664 54874
rect -3738 54806 -3718 54840
rect -3684 54806 -3664 54840
rect -3738 54772 -3664 54806
rect -3738 54738 -3718 54772
rect -3684 54738 -3664 54772
rect -3738 54704 -3664 54738
rect -3738 54670 -3718 54704
rect -3684 54670 -3664 54704
rect -3738 54636 -3664 54670
rect -3738 54602 -3718 54636
rect -3684 54602 -3664 54636
rect -3738 54568 -3664 54602
rect -3738 54534 -3718 54568
rect -3684 54534 -3664 54568
rect -3738 54500 -3664 54534
rect -3738 54466 -3718 54500
rect -3684 54466 -3664 54500
rect -3738 54432 -3664 54466
rect -3738 54398 -3718 54432
rect -3684 54398 -3664 54432
rect -3738 54364 -3664 54398
rect -3738 54330 -3718 54364
rect -3684 54330 -3664 54364
rect -3738 54296 -3664 54330
rect -3738 54262 -3718 54296
rect -3684 54262 -3664 54296
rect -3738 54228 -3664 54262
rect -3738 54194 -3718 54228
rect -3684 54194 -3664 54228
rect -3738 54160 -3664 54194
rect -3738 54126 -3718 54160
rect -3684 54126 -3664 54160
rect -3738 54092 -3664 54126
rect -3738 54058 -3718 54092
rect -3684 54058 -3664 54092
rect -3738 54024 -3664 54058
rect -3738 53990 -3718 54024
rect -3684 53990 -3664 54024
rect -3738 53956 -3664 53990
rect -3738 53922 -3718 53956
rect -3684 53922 -3664 53956
rect -3738 53888 -3664 53922
rect -3738 53854 -3718 53888
rect -3684 53854 -3664 53888
rect -3738 53820 -3664 53854
rect -3738 53786 -3718 53820
rect -3684 53786 -3664 53820
rect -3738 53752 -3664 53786
rect -3738 53718 -3718 53752
rect -3684 53718 -3664 53752
rect -3738 53684 -3664 53718
rect -3738 53650 -3718 53684
rect -3684 53650 -3664 53684
rect -3738 53616 -3664 53650
rect -3738 53582 -3718 53616
rect -3684 53582 -3664 53616
rect -3738 53548 -3664 53582
rect -3738 53514 -3718 53548
rect -3684 53514 -3664 53548
rect -3738 53480 -3664 53514
rect -3738 53446 -3718 53480
rect -3684 53446 -3664 53480
rect -3738 53412 -3664 53446
rect -3738 53378 -3718 53412
rect -3684 53378 -3664 53412
rect -3738 53344 -3664 53378
rect -3738 53310 -3718 53344
rect -3684 53310 -3664 53344
rect -3738 53276 -3664 53310
rect -3738 53242 -3718 53276
rect -3684 53242 -3664 53276
rect -3738 53208 -3664 53242
rect -3738 53174 -3718 53208
rect -3684 53174 -3664 53208
rect -3738 53140 -3664 53174
rect -3738 53106 -3718 53140
rect -3684 53106 -3664 53140
rect -3738 53072 -3664 53106
rect -3738 53038 -3718 53072
rect -3684 53038 -3664 53072
rect -3738 53004 -3664 53038
rect -3738 52970 -3718 53004
rect -3684 52970 -3664 53004
rect -3738 52936 -3664 52970
rect -3738 52902 -3718 52936
rect -3684 52902 -3664 52936
rect -3738 52868 -3664 52902
rect -3738 52834 -3718 52868
rect -3684 52834 -3664 52868
rect -3738 52800 -3664 52834
rect -3738 52766 -3718 52800
rect -3684 52766 -3664 52800
rect -3738 52732 -3664 52766
rect -3738 52698 -3718 52732
rect -3684 52698 -3664 52732
rect -3738 52664 -3664 52698
rect -3738 52630 -3718 52664
rect -3684 52630 -3664 52664
rect -3738 52596 -3664 52630
rect -3738 52562 -3718 52596
rect -3684 52562 -3664 52596
rect -3738 52528 -3664 52562
rect -3738 52494 -3718 52528
rect -3684 52494 -3664 52528
rect -3738 52460 -3664 52494
rect -3738 52426 -3718 52460
rect -3684 52426 -3664 52460
rect -3738 52392 -3664 52426
rect -3738 52358 -3718 52392
rect -3684 52358 -3664 52392
rect -3738 52324 -3664 52358
rect -3738 52290 -3718 52324
rect -3684 52290 -3664 52324
rect -3738 52256 -3664 52290
rect -3738 52222 -3718 52256
rect -3684 52222 -3664 52256
rect -3738 52188 -3664 52222
rect -3738 52154 -3718 52188
rect -3684 52154 -3664 52188
rect -3738 52120 -3664 52154
rect -3738 52086 -3718 52120
rect -3684 52086 -3664 52120
rect -3738 52052 -3664 52086
rect -3738 52018 -3718 52052
rect -3684 52018 -3664 52052
rect -3738 51984 -3664 52018
rect -3738 51950 -3718 51984
rect -3684 51950 -3664 51984
rect -3738 51916 -3664 51950
rect -3738 51882 -3718 51916
rect -3684 51882 -3664 51916
rect -3738 51848 -3664 51882
rect -3738 51814 -3718 51848
rect -3684 51814 -3664 51848
rect -3738 51780 -3664 51814
rect -3738 51746 -3718 51780
rect -3684 51746 -3664 51780
rect -3738 51712 -3664 51746
rect -3738 51678 -3718 51712
rect -3684 51678 -3664 51712
rect -3738 51644 -3664 51678
rect -3738 51610 -3718 51644
rect -3684 51610 -3664 51644
rect -3738 51576 -3664 51610
rect -3738 51542 -3718 51576
rect -3684 51542 -3664 51576
rect -3738 51508 -3664 51542
rect -3738 51474 -3718 51508
rect -3684 51474 -3664 51508
rect -3738 51440 -3664 51474
rect -3738 51406 -3718 51440
rect -3684 51406 -3664 51440
rect -3738 51372 -3664 51406
rect -3738 51338 -3718 51372
rect -3684 51338 -3664 51372
rect -3738 51304 -3664 51338
rect -3738 51270 -3718 51304
rect -3684 51270 -3664 51304
rect -3738 51236 -3664 51270
rect -3738 51202 -3718 51236
rect -3684 51202 -3664 51236
rect -3738 51168 -3664 51202
rect -3738 51134 -3718 51168
rect -3684 51134 -3664 51168
rect -3738 51100 -3664 51134
rect -3738 51066 -3718 51100
rect -3684 51066 -3664 51100
rect -3738 51032 -3664 51066
rect -3738 50998 -3718 51032
rect -3684 50998 -3664 51032
rect -3738 50964 -3664 50998
rect -3738 50930 -3718 50964
rect -3684 50930 -3664 50964
rect -3738 50896 -3664 50930
rect -3738 50862 -3718 50896
rect -3684 50862 -3664 50896
rect -3738 50828 -3664 50862
rect -3738 50794 -3718 50828
rect -3684 50794 -3664 50828
rect -3738 50760 -3664 50794
rect -3738 50726 -3718 50760
rect -3684 50726 -3664 50760
rect -3738 50692 -3664 50726
rect -3738 50658 -3718 50692
rect -3684 50658 -3664 50692
rect -3738 50624 -3664 50658
rect -3738 50590 -3718 50624
rect -3684 50590 -3664 50624
rect -3738 50556 -3664 50590
rect -3738 50522 -3718 50556
rect -3684 50522 -3664 50556
rect -3738 50488 -3664 50522
rect -3738 50454 -3718 50488
rect -3684 50454 -3664 50488
rect -3738 50420 -3664 50454
rect -3738 50386 -3718 50420
rect -3684 50386 -3664 50420
rect -3738 50352 -3664 50386
rect -3738 50318 -3718 50352
rect -3684 50318 -3664 50352
rect -3738 50284 -3664 50318
rect -3738 50250 -3718 50284
rect -3684 50250 -3664 50284
rect -3738 50216 -3664 50250
rect -3738 50182 -3718 50216
rect -3684 50182 -3664 50216
rect -3738 50148 -3664 50182
rect -3738 50114 -3718 50148
rect -3684 50114 -3664 50148
rect -3738 50080 -3664 50114
rect -3738 50046 -3718 50080
rect -3684 50046 -3664 50080
rect -3738 50012 -3664 50046
rect -3738 49978 -3718 50012
rect -3684 49978 -3664 50012
rect -3738 49944 -3664 49978
rect -3738 49910 -3718 49944
rect -3684 49910 -3664 49944
rect -3738 49876 -3664 49910
rect -3738 49842 -3718 49876
rect -3684 49842 -3664 49876
rect -3738 49808 -3664 49842
rect -3738 49774 -3718 49808
rect -3684 49774 -3664 49808
rect -3738 49740 -3664 49774
rect -3738 49706 -3718 49740
rect -3684 49706 -3664 49740
rect -3738 49672 -3664 49706
rect -3738 49638 -3718 49672
rect -3684 49638 -3664 49672
rect -3738 49604 -3664 49638
rect -3738 49570 -3718 49604
rect -3684 49570 -3664 49604
rect -3738 49536 -3664 49570
rect -3738 49502 -3718 49536
rect -3684 49502 -3664 49536
rect -3738 49468 -3664 49502
rect -3738 49434 -3718 49468
rect -3684 49434 -3664 49468
rect -3738 49400 -3664 49434
rect -3738 49366 -3718 49400
rect -3684 49366 -3664 49400
rect -3738 49332 -3664 49366
rect -3738 49298 -3718 49332
rect -3684 49298 -3664 49332
rect -3738 49264 -3664 49298
rect -3738 49230 -3718 49264
rect -3684 49230 -3664 49264
rect -3738 49196 -3664 49230
rect -3738 49162 -3718 49196
rect -3684 49162 -3664 49196
rect -3738 49128 -3664 49162
rect -3738 49094 -3718 49128
rect -3684 49094 -3664 49128
rect -3738 49060 -3664 49094
rect -3738 49026 -3718 49060
rect -3684 49026 -3664 49060
rect -3738 48992 -3664 49026
rect -3738 48958 -3718 48992
rect -3684 48958 -3664 48992
rect -3738 48924 -3664 48958
rect -3738 48890 -3718 48924
rect -3684 48890 -3664 48924
rect -3738 48856 -3664 48890
rect -3738 48822 -3718 48856
rect -3684 48822 -3664 48856
rect -3738 48788 -3664 48822
rect -3738 48754 -3718 48788
rect -3684 48754 -3664 48788
rect -3738 48720 -3664 48754
rect -3738 48686 -3718 48720
rect -3684 48686 -3664 48720
rect -3738 48652 -3664 48686
rect -3738 48618 -3718 48652
rect -3684 48618 -3664 48652
rect -3738 48584 -3664 48618
rect -3738 48550 -3718 48584
rect -3684 48550 -3664 48584
rect -3738 48516 -3664 48550
rect -3738 48482 -3718 48516
rect -3684 48482 -3664 48516
rect -3738 48448 -3664 48482
rect -3738 48414 -3718 48448
rect -3684 48414 -3664 48448
rect -3738 48380 -3664 48414
rect -3738 48346 -3718 48380
rect -3684 48346 -3664 48380
rect -3738 48312 -3664 48346
rect -3738 48278 -3718 48312
rect -3684 48278 -3664 48312
rect -3738 48244 -3664 48278
rect -3738 48210 -3718 48244
rect -3684 48210 -3664 48244
rect -3738 48176 -3664 48210
rect -3738 48142 -3718 48176
rect -3684 48142 -3664 48176
rect -3738 48108 -3664 48142
rect -3738 48074 -3718 48108
rect -3684 48074 -3664 48108
rect -3738 48040 -3664 48074
rect -3738 48006 -3718 48040
rect -3684 48006 -3664 48040
rect -3738 47972 -3664 48006
rect -3738 47938 -3718 47972
rect -3684 47938 -3664 47972
rect -3738 47904 -3664 47938
rect -3738 47870 -3718 47904
rect -3684 47870 -3664 47904
rect -3738 47836 -3664 47870
rect -3738 47802 -3718 47836
rect -3684 47802 -3664 47836
rect -3738 47768 -3664 47802
rect -3738 47734 -3718 47768
rect -3684 47734 -3664 47768
rect -3738 47700 -3664 47734
rect -3738 47666 -3718 47700
rect -3684 47666 -3664 47700
rect -3738 47632 -3664 47666
rect -3738 47598 -3718 47632
rect -3684 47598 -3664 47632
rect -3738 47564 -3664 47598
rect -3738 47530 -3718 47564
rect -3684 47530 -3664 47564
rect -3738 47496 -3664 47530
rect -3738 47462 -3718 47496
rect -3684 47462 -3664 47496
rect -3738 47428 -3664 47462
rect -3738 47394 -3718 47428
rect -3684 47394 -3664 47428
rect -3738 47360 -3664 47394
rect -3738 47326 -3718 47360
rect -3684 47326 -3664 47360
rect -3738 47292 -3664 47326
rect -3738 47258 -3718 47292
rect -3684 47258 -3664 47292
rect -3738 47224 -3664 47258
rect -3738 47190 -3718 47224
rect -3684 47190 -3664 47224
rect -3738 47156 -3664 47190
rect -3738 47122 -3718 47156
rect -3684 47122 -3664 47156
rect -3738 47088 -3664 47122
rect -3738 47054 -3718 47088
rect -3684 47054 -3664 47088
rect -3738 47020 -3664 47054
rect -3738 46986 -3718 47020
rect -3684 46986 -3664 47020
rect -3738 46952 -3664 46986
rect -3738 46918 -3718 46952
rect -3684 46918 -3664 46952
rect -3738 46884 -3664 46918
rect -3738 46850 -3718 46884
rect -3684 46850 -3664 46884
rect -3738 46816 -3664 46850
rect -3738 46782 -3718 46816
rect -3684 46782 -3664 46816
rect -3738 46748 -3664 46782
rect -3738 46714 -3718 46748
rect -3684 46714 -3664 46748
rect -3738 46680 -3664 46714
rect -3738 46646 -3718 46680
rect -3684 46646 -3664 46680
rect -3738 46612 -3664 46646
rect -3738 46578 -3718 46612
rect -3684 46578 -3664 46612
rect -3738 46544 -3664 46578
rect -3738 46510 -3718 46544
rect -3684 46510 -3664 46544
rect -3738 46476 -3664 46510
rect -3738 46442 -3718 46476
rect -3684 46442 -3664 46476
rect -3738 46408 -3664 46442
rect -3738 46374 -3718 46408
rect -3684 46374 -3664 46408
rect -3738 46340 -3664 46374
rect -3738 46306 -3718 46340
rect -3684 46306 -3664 46340
rect -3738 46272 -3664 46306
rect -3738 46238 -3718 46272
rect -3684 46238 -3664 46272
rect -3738 46204 -3664 46238
rect -3738 46170 -3718 46204
rect -3684 46170 -3664 46204
rect -3738 46136 -3664 46170
rect -3738 46102 -3718 46136
rect -3684 46102 -3664 46136
rect -3738 46068 -3664 46102
rect -3738 46034 -3718 46068
rect -3684 46034 -3664 46068
rect -3738 46000 -3664 46034
rect -3738 45966 -3718 46000
rect -3684 45966 -3664 46000
rect -3738 45932 -3664 45966
rect -3738 45898 -3718 45932
rect -3684 45898 -3664 45932
rect -3738 45864 -3664 45898
rect 59084 58289 59158 58323
rect 59084 58255 59104 58289
rect 59138 58255 59158 58289
rect 59084 58221 59158 58255
rect 59084 58187 59104 58221
rect 59138 58187 59158 58221
rect 59084 58153 59158 58187
rect 59084 58119 59104 58153
rect 59138 58119 59158 58153
rect 59084 58085 59158 58119
rect 59084 58051 59104 58085
rect 59138 58051 59158 58085
rect 59084 58017 59158 58051
rect 59084 57983 59104 58017
rect 59138 57983 59158 58017
rect 59084 57949 59158 57983
rect 59084 57915 59104 57949
rect 59138 57915 59158 57949
rect 59084 57881 59158 57915
rect 59084 57847 59104 57881
rect 59138 57847 59158 57881
rect 59084 57813 59158 57847
rect 59084 57779 59104 57813
rect 59138 57779 59158 57813
rect 59084 57745 59158 57779
rect 59084 57711 59104 57745
rect 59138 57711 59158 57745
rect 59084 57677 59158 57711
rect 59084 57643 59104 57677
rect 59138 57643 59158 57677
rect 59084 57609 59158 57643
rect 59084 57575 59104 57609
rect 59138 57575 59158 57609
rect 59084 57541 59158 57575
rect 59084 57507 59104 57541
rect 59138 57507 59158 57541
rect 59084 57473 59158 57507
rect 59084 57439 59104 57473
rect 59138 57439 59158 57473
rect 59084 57405 59158 57439
rect 59084 57371 59104 57405
rect 59138 57371 59158 57405
rect 59084 57337 59158 57371
rect 59084 57303 59104 57337
rect 59138 57303 59158 57337
rect 59084 57269 59158 57303
rect 59084 57235 59104 57269
rect 59138 57235 59158 57269
rect 59084 57201 59158 57235
rect 59084 57167 59104 57201
rect 59138 57167 59158 57201
rect 59084 57133 59158 57167
rect 59084 57099 59104 57133
rect 59138 57099 59158 57133
rect 59084 57065 59158 57099
rect 59084 57031 59104 57065
rect 59138 57031 59158 57065
rect 59084 56997 59158 57031
rect 59084 56963 59104 56997
rect 59138 56963 59158 56997
rect 59084 56929 59158 56963
rect 59084 56895 59104 56929
rect 59138 56895 59158 56929
rect 59084 56861 59158 56895
rect 59084 56827 59104 56861
rect 59138 56827 59158 56861
rect 59084 56793 59158 56827
rect 59084 56759 59104 56793
rect 59138 56759 59158 56793
rect 59084 56725 59158 56759
rect 59084 56691 59104 56725
rect 59138 56691 59158 56725
rect 59084 56657 59158 56691
rect 59084 56623 59104 56657
rect 59138 56623 59158 56657
rect 59084 56589 59158 56623
rect 59084 56555 59104 56589
rect 59138 56555 59158 56589
rect 59084 56521 59158 56555
rect 59084 56487 59104 56521
rect 59138 56487 59158 56521
rect 59084 56453 59158 56487
rect 59084 56419 59104 56453
rect 59138 56419 59158 56453
rect 59084 56385 59158 56419
rect 59084 56351 59104 56385
rect 59138 56351 59158 56385
rect 59084 56317 59158 56351
rect 59084 56283 59104 56317
rect 59138 56283 59158 56317
rect 59084 56249 59158 56283
rect 59084 56215 59104 56249
rect 59138 56215 59158 56249
rect 59084 56181 59158 56215
rect 59084 56147 59104 56181
rect 59138 56147 59158 56181
rect 59084 56113 59158 56147
rect 59084 56079 59104 56113
rect 59138 56079 59158 56113
rect 59084 56045 59158 56079
rect 59084 56011 59104 56045
rect 59138 56011 59158 56045
rect 59084 55977 59158 56011
rect 59084 55943 59104 55977
rect 59138 55943 59158 55977
rect 59084 55909 59158 55943
rect 59084 55875 59104 55909
rect 59138 55875 59158 55909
rect 59084 55841 59158 55875
rect 59084 55807 59104 55841
rect 59138 55807 59158 55841
rect 59084 55773 59158 55807
rect 59084 55739 59104 55773
rect 59138 55739 59158 55773
rect 59084 55705 59158 55739
rect 59084 55671 59104 55705
rect 59138 55671 59158 55705
rect 59084 55637 59158 55671
rect 59084 55603 59104 55637
rect 59138 55603 59158 55637
rect 59084 55569 59158 55603
rect 59084 55535 59104 55569
rect 59138 55535 59158 55569
rect 59084 55501 59158 55535
rect 59084 55467 59104 55501
rect 59138 55467 59158 55501
rect 59084 55433 59158 55467
rect 59084 55399 59104 55433
rect 59138 55399 59158 55433
rect 59084 55365 59158 55399
rect 59084 55331 59104 55365
rect 59138 55331 59158 55365
rect 59084 55297 59158 55331
rect 59084 55263 59104 55297
rect 59138 55263 59158 55297
rect 59084 55229 59158 55263
rect 59084 55195 59104 55229
rect 59138 55195 59158 55229
rect 59084 55161 59158 55195
rect 59084 55127 59104 55161
rect 59138 55127 59158 55161
rect 59084 55093 59158 55127
rect 59084 55059 59104 55093
rect 59138 55059 59158 55093
rect 59084 55025 59158 55059
rect 59084 54991 59104 55025
rect 59138 54991 59158 55025
rect 59084 54957 59158 54991
rect 59084 54923 59104 54957
rect 59138 54923 59158 54957
rect 59084 54889 59158 54923
rect 59084 54855 59104 54889
rect 59138 54855 59158 54889
rect 59084 54821 59158 54855
rect 59084 54787 59104 54821
rect 59138 54787 59158 54821
rect 59084 54753 59158 54787
rect 59084 54719 59104 54753
rect 59138 54719 59158 54753
rect 59084 54685 59158 54719
rect 59084 54651 59104 54685
rect 59138 54651 59158 54685
rect 59084 54617 59158 54651
rect 59084 54583 59104 54617
rect 59138 54583 59158 54617
rect 59084 54549 59158 54583
rect 59084 54515 59104 54549
rect 59138 54515 59158 54549
rect 59084 54481 59158 54515
rect 59084 54447 59104 54481
rect 59138 54447 59158 54481
rect 59084 54413 59158 54447
rect 59084 54379 59104 54413
rect 59138 54379 59158 54413
rect 59084 54345 59158 54379
rect 59084 54311 59104 54345
rect 59138 54311 59158 54345
rect 59084 54277 59158 54311
rect 59084 54243 59104 54277
rect 59138 54243 59158 54277
rect 59084 54209 59158 54243
rect 59084 54175 59104 54209
rect 59138 54175 59158 54209
rect 59084 54141 59158 54175
rect 59084 54107 59104 54141
rect 59138 54107 59158 54141
rect 59084 54073 59158 54107
rect 59084 54039 59104 54073
rect 59138 54039 59158 54073
rect 59084 54005 59158 54039
rect 59084 53971 59104 54005
rect 59138 53971 59158 54005
rect 59084 53937 59158 53971
rect 59084 53903 59104 53937
rect 59138 53903 59158 53937
rect 59084 53869 59158 53903
rect 59084 53835 59104 53869
rect 59138 53835 59158 53869
rect 59084 53801 59158 53835
rect 59084 53767 59104 53801
rect 59138 53767 59158 53801
rect 59084 53733 59158 53767
rect 59084 53699 59104 53733
rect 59138 53699 59158 53733
rect 59084 53665 59158 53699
rect 59084 53631 59104 53665
rect 59138 53631 59158 53665
rect 59084 53597 59158 53631
rect 59084 53563 59104 53597
rect 59138 53563 59158 53597
rect 59084 53529 59158 53563
rect 59084 53495 59104 53529
rect 59138 53495 59158 53529
rect 59084 53461 59158 53495
rect 59084 53427 59104 53461
rect 59138 53427 59158 53461
rect 59084 53393 59158 53427
rect 59084 53359 59104 53393
rect 59138 53359 59158 53393
rect 59084 53325 59158 53359
rect 59084 53291 59104 53325
rect 59138 53291 59158 53325
rect 59084 53257 59158 53291
rect 59084 53223 59104 53257
rect 59138 53223 59158 53257
rect 59084 53189 59158 53223
rect 59084 53155 59104 53189
rect 59138 53155 59158 53189
rect 59084 53121 59158 53155
rect 59084 53087 59104 53121
rect 59138 53087 59158 53121
rect 59084 53053 59158 53087
rect 59084 53019 59104 53053
rect 59138 53019 59158 53053
rect 59084 52985 59158 53019
rect 59084 52951 59104 52985
rect 59138 52951 59158 52985
rect 59084 52917 59158 52951
rect 59084 52883 59104 52917
rect 59138 52883 59158 52917
rect 59084 52849 59158 52883
rect 59084 52815 59104 52849
rect 59138 52815 59158 52849
rect 59084 52781 59158 52815
rect 59084 52747 59104 52781
rect 59138 52747 59158 52781
rect 59084 52713 59158 52747
rect 59084 52679 59104 52713
rect 59138 52679 59158 52713
rect 59084 52645 59158 52679
rect 59084 52611 59104 52645
rect 59138 52611 59158 52645
rect 59084 52577 59158 52611
rect 59084 52543 59104 52577
rect 59138 52543 59158 52577
rect 59084 52509 59158 52543
rect 59084 52475 59104 52509
rect 59138 52475 59158 52509
rect 59084 52441 59158 52475
rect 59084 52407 59104 52441
rect 59138 52407 59158 52441
rect 59084 52373 59158 52407
rect 59084 52339 59104 52373
rect 59138 52339 59158 52373
rect 59084 52305 59158 52339
rect 59084 52271 59104 52305
rect 59138 52271 59158 52305
rect 59084 52237 59158 52271
rect 59084 52203 59104 52237
rect 59138 52203 59158 52237
rect 59084 52169 59158 52203
rect 59084 52135 59104 52169
rect 59138 52135 59158 52169
rect 59084 52101 59158 52135
rect 59084 52067 59104 52101
rect 59138 52067 59158 52101
rect 59084 52033 59158 52067
rect 59084 51999 59104 52033
rect 59138 51999 59158 52033
rect 59084 51965 59158 51999
rect 59084 51931 59104 51965
rect 59138 51931 59158 51965
rect 59084 51897 59158 51931
rect 59084 51863 59104 51897
rect 59138 51863 59158 51897
rect 59084 51829 59158 51863
rect 59084 51795 59104 51829
rect 59138 51795 59158 51829
rect 59084 51761 59158 51795
rect 59084 51727 59104 51761
rect 59138 51727 59158 51761
rect 59084 51693 59158 51727
rect 59084 51659 59104 51693
rect 59138 51659 59158 51693
rect 59084 51625 59158 51659
rect 59084 51591 59104 51625
rect 59138 51591 59158 51625
rect 59084 51557 59158 51591
rect 59084 51523 59104 51557
rect 59138 51523 59158 51557
rect 59084 51489 59158 51523
rect 59084 51455 59104 51489
rect 59138 51455 59158 51489
rect 59084 51421 59158 51455
rect 59084 51387 59104 51421
rect 59138 51387 59158 51421
rect 59084 51353 59158 51387
rect 59084 51319 59104 51353
rect 59138 51319 59158 51353
rect 59084 51285 59158 51319
rect 59084 51251 59104 51285
rect 59138 51251 59158 51285
rect 59084 51217 59158 51251
rect 59084 51183 59104 51217
rect 59138 51183 59158 51217
rect 59084 51149 59158 51183
rect 59084 51115 59104 51149
rect 59138 51115 59158 51149
rect 59084 51081 59158 51115
rect 59084 51047 59104 51081
rect 59138 51047 59158 51081
rect 59084 51013 59158 51047
rect 59084 50979 59104 51013
rect 59138 50979 59158 51013
rect 59084 50945 59158 50979
rect 59084 50911 59104 50945
rect 59138 50911 59158 50945
rect 59084 50877 59158 50911
rect 59084 50843 59104 50877
rect 59138 50843 59158 50877
rect 59084 50809 59158 50843
rect 59084 50775 59104 50809
rect 59138 50775 59158 50809
rect 59084 50741 59158 50775
rect 59084 50707 59104 50741
rect 59138 50707 59158 50741
rect 59084 50673 59158 50707
rect 59084 50639 59104 50673
rect 59138 50639 59158 50673
rect 59084 50605 59158 50639
rect 59084 50571 59104 50605
rect 59138 50571 59158 50605
rect 59084 50537 59158 50571
rect 59084 50503 59104 50537
rect 59138 50503 59158 50537
rect 59084 50469 59158 50503
rect 59084 50435 59104 50469
rect 59138 50435 59158 50469
rect 59084 50401 59158 50435
rect 59084 50367 59104 50401
rect 59138 50367 59158 50401
rect 59084 50333 59158 50367
rect 59084 50299 59104 50333
rect 59138 50299 59158 50333
rect 59084 50265 59158 50299
rect 59084 50231 59104 50265
rect 59138 50231 59158 50265
rect 59084 50197 59158 50231
rect 59084 50163 59104 50197
rect 59138 50163 59158 50197
rect 59084 50129 59158 50163
rect 59084 50095 59104 50129
rect 59138 50095 59158 50129
rect 59084 50061 59158 50095
rect 59084 50027 59104 50061
rect 59138 50027 59158 50061
rect 59084 49993 59158 50027
rect 59084 49959 59104 49993
rect 59138 49959 59158 49993
rect 59084 49925 59158 49959
rect 59084 49891 59104 49925
rect 59138 49891 59158 49925
rect 59084 49857 59158 49891
rect 59084 49823 59104 49857
rect 59138 49823 59158 49857
rect 59084 49789 59158 49823
rect 59084 49755 59104 49789
rect 59138 49755 59158 49789
rect 59084 49721 59158 49755
rect 59084 49687 59104 49721
rect 59138 49687 59158 49721
rect 59084 49653 59158 49687
rect 59084 49619 59104 49653
rect 59138 49619 59158 49653
rect 59084 49585 59158 49619
rect 59084 49551 59104 49585
rect 59138 49551 59158 49585
rect 59084 49517 59158 49551
rect 59084 49483 59104 49517
rect 59138 49483 59158 49517
rect 59084 49449 59158 49483
rect 59084 49415 59104 49449
rect 59138 49415 59158 49449
rect 59084 49381 59158 49415
rect 59084 49347 59104 49381
rect 59138 49347 59158 49381
rect 59084 49313 59158 49347
rect 59084 49279 59104 49313
rect 59138 49279 59158 49313
rect 59084 49245 59158 49279
rect 59084 49211 59104 49245
rect 59138 49211 59158 49245
rect 59084 49177 59158 49211
rect 59084 49143 59104 49177
rect 59138 49143 59158 49177
rect 59084 49109 59158 49143
rect 59084 49075 59104 49109
rect 59138 49075 59158 49109
rect 59084 49041 59158 49075
rect 59084 49007 59104 49041
rect 59138 49007 59158 49041
rect 59084 48973 59158 49007
rect 59084 48939 59104 48973
rect 59138 48939 59158 48973
rect 59084 48905 59158 48939
rect 59084 48871 59104 48905
rect 59138 48871 59158 48905
rect 59084 48837 59158 48871
rect 59084 48803 59104 48837
rect 59138 48803 59158 48837
rect 59084 48769 59158 48803
rect 59084 48735 59104 48769
rect 59138 48735 59158 48769
rect 59084 48701 59158 48735
rect 59084 48667 59104 48701
rect 59138 48667 59158 48701
rect 59084 48633 59158 48667
rect 59084 48599 59104 48633
rect 59138 48599 59158 48633
rect 59084 48565 59158 48599
rect 59084 48531 59104 48565
rect 59138 48531 59158 48565
rect 59084 48497 59158 48531
rect 59084 48463 59104 48497
rect 59138 48463 59158 48497
rect 59084 48429 59158 48463
rect 59084 48395 59104 48429
rect 59138 48395 59158 48429
rect 59084 48361 59158 48395
rect 59084 48327 59104 48361
rect 59138 48327 59158 48361
rect 59084 48293 59158 48327
rect 59084 48259 59104 48293
rect 59138 48259 59158 48293
rect 59084 48225 59158 48259
rect 59084 48191 59104 48225
rect 59138 48191 59158 48225
rect 59084 48157 59158 48191
rect 59084 48123 59104 48157
rect 59138 48123 59158 48157
rect 59084 48089 59158 48123
rect 59084 48055 59104 48089
rect 59138 48055 59158 48089
rect 59084 48021 59158 48055
rect 59084 47987 59104 48021
rect 59138 47987 59158 48021
rect 59084 47953 59158 47987
rect 59084 47919 59104 47953
rect 59138 47919 59158 47953
rect 59084 47885 59158 47919
rect 59084 47851 59104 47885
rect 59138 47851 59158 47885
rect 59084 47817 59158 47851
rect 59084 47783 59104 47817
rect 59138 47783 59158 47817
rect 59084 47749 59158 47783
rect 59084 47715 59104 47749
rect 59138 47715 59158 47749
rect 59084 47681 59158 47715
rect 59084 47647 59104 47681
rect 59138 47647 59158 47681
rect 59084 47613 59158 47647
rect 59084 47579 59104 47613
rect 59138 47579 59158 47613
rect 59084 47545 59158 47579
rect 59084 47511 59104 47545
rect 59138 47511 59158 47545
rect 59084 47477 59158 47511
rect 59084 47443 59104 47477
rect 59138 47443 59158 47477
rect 59084 47409 59158 47443
rect 59084 47375 59104 47409
rect 59138 47375 59158 47409
rect 59084 47341 59158 47375
rect 59084 47307 59104 47341
rect 59138 47307 59158 47341
rect 59084 47273 59158 47307
rect 59084 47239 59104 47273
rect 59138 47239 59158 47273
rect 59084 47205 59158 47239
rect 59084 47171 59104 47205
rect 59138 47171 59158 47205
rect 59084 47137 59158 47171
rect 59084 47103 59104 47137
rect 59138 47103 59158 47137
rect 59084 47069 59158 47103
rect 59084 47035 59104 47069
rect 59138 47035 59158 47069
rect 59084 47001 59158 47035
rect 59084 46967 59104 47001
rect 59138 46967 59158 47001
rect 59084 46933 59158 46967
rect 59084 46899 59104 46933
rect 59138 46899 59158 46933
rect 59084 46865 59158 46899
rect 59084 46831 59104 46865
rect 59138 46831 59158 46865
rect 59084 46797 59158 46831
rect 59084 46763 59104 46797
rect 59138 46763 59158 46797
rect 59084 46729 59158 46763
rect 59084 46695 59104 46729
rect 59138 46695 59158 46729
rect 59084 46661 59158 46695
rect 59084 46627 59104 46661
rect 59138 46627 59158 46661
rect 59084 46593 59158 46627
rect 59084 46559 59104 46593
rect 59138 46559 59158 46593
rect 59084 46525 59158 46559
rect 59084 46491 59104 46525
rect 59138 46491 59158 46525
rect 59084 46457 59158 46491
rect 59084 46423 59104 46457
rect 59138 46423 59158 46457
rect 59084 46389 59158 46423
rect 59084 46355 59104 46389
rect 59138 46355 59158 46389
rect 59084 46321 59158 46355
rect 59084 46287 59104 46321
rect 59138 46287 59158 46321
rect 59084 46253 59158 46287
rect 59084 46219 59104 46253
rect 59138 46219 59158 46253
rect 59084 46185 59158 46219
rect 59084 46151 59104 46185
rect 59138 46151 59158 46185
rect 59084 46117 59158 46151
rect 59084 46083 59104 46117
rect 59138 46083 59158 46117
rect 59084 46049 59158 46083
rect 59084 46015 59104 46049
rect 59138 46015 59158 46049
rect 59084 45981 59158 46015
rect 59084 45947 59104 45981
rect 59138 45947 59158 45981
rect 59084 45940 59158 45947
rect 70818 74745 70892 74752
rect 70818 74711 70838 74745
rect 70872 74711 70892 74745
rect 70818 74677 70892 74711
rect 70818 74643 70838 74677
rect 70872 74643 70892 74677
rect 70818 74609 70892 74643
rect 70818 74575 70838 74609
rect 70872 74575 70892 74609
rect 70818 74541 70892 74575
rect 70818 74507 70838 74541
rect 70872 74507 70892 74541
rect 70818 74473 70892 74507
rect 70818 74439 70838 74473
rect 70872 74439 70892 74473
rect 70818 74405 70892 74439
rect 70818 74371 70838 74405
rect 70872 74371 70892 74405
rect 70818 74337 70892 74371
rect 70818 74303 70838 74337
rect 70872 74303 70892 74337
rect 70818 74269 70892 74303
rect 70818 74235 70838 74269
rect 70872 74235 70892 74269
rect 70818 74201 70892 74235
rect 70818 74167 70838 74201
rect 70872 74167 70892 74201
rect 70818 74133 70892 74167
rect 70818 74099 70838 74133
rect 70872 74099 70892 74133
rect 70818 74065 70892 74099
rect 70818 74031 70838 74065
rect 70872 74031 70892 74065
rect 70818 73997 70892 74031
rect 70818 73963 70838 73997
rect 70872 73963 70892 73997
rect 70818 73929 70892 73963
rect 70818 73895 70838 73929
rect 70872 73895 70892 73929
rect 70818 73861 70892 73895
rect 70818 73827 70838 73861
rect 70872 73827 70892 73861
rect 70818 73793 70892 73827
rect 70818 73759 70838 73793
rect 70872 73759 70892 73793
rect 70818 73725 70892 73759
rect 70818 73691 70838 73725
rect 70872 73691 70892 73725
rect 70818 73657 70892 73691
rect 70818 73623 70838 73657
rect 70872 73623 70892 73657
rect 70818 73589 70892 73623
rect 70818 73555 70838 73589
rect 70872 73555 70892 73589
rect 70818 73521 70892 73555
rect 70818 73487 70838 73521
rect 70872 73487 70892 73521
rect 70818 73453 70892 73487
rect 70818 73419 70838 73453
rect 70872 73419 70892 73453
rect 70818 73385 70892 73419
rect 70818 73351 70838 73385
rect 70872 73351 70892 73385
rect 70818 73317 70892 73351
rect 70818 73283 70838 73317
rect 70872 73283 70892 73317
rect 70818 73249 70892 73283
rect 70818 73215 70838 73249
rect 70872 73215 70892 73249
rect 70818 73181 70892 73215
rect 70818 73147 70838 73181
rect 70872 73147 70892 73181
rect 70818 73113 70892 73147
rect 70818 73079 70838 73113
rect 70872 73079 70892 73113
rect 70818 73045 70892 73079
rect 70818 73011 70838 73045
rect 70872 73011 70892 73045
rect 70818 72977 70892 73011
rect 70818 72943 70838 72977
rect 70872 72943 70892 72977
rect 70818 72909 70892 72943
rect 70818 72875 70838 72909
rect 70872 72875 70892 72909
rect 70818 72841 70892 72875
rect 70818 72807 70838 72841
rect 70872 72807 70892 72841
rect 70818 72773 70892 72807
rect 70818 72739 70838 72773
rect 70872 72739 70892 72773
rect 70818 72705 70892 72739
rect 70818 72671 70838 72705
rect 70872 72671 70892 72705
rect 70818 72637 70892 72671
rect 70818 72603 70838 72637
rect 70872 72603 70892 72637
rect 70818 72569 70892 72603
rect 70818 72535 70838 72569
rect 70872 72535 70892 72569
rect 70818 72501 70892 72535
rect 70818 72467 70838 72501
rect 70872 72467 70892 72501
rect 70818 72433 70892 72467
rect 70818 72399 70838 72433
rect 70872 72399 70892 72433
rect 70818 72365 70892 72399
rect 70818 72331 70838 72365
rect 70872 72331 70892 72365
rect 70818 72297 70892 72331
rect 70818 72263 70838 72297
rect 70872 72263 70892 72297
rect 70818 72229 70892 72263
rect 70818 72195 70838 72229
rect 70872 72195 70892 72229
rect 70818 72161 70892 72195
rect 70818 72127 70838 72161
rect 70872 72127 70892 72161
rect 70818 72093 70892 72127
rect 70818 72059 70838 72093
rect 70872 72059 70892 72093
rect 70818 72025 70892 72059
rect 70818 71991 70838 72025
rect 70872 71991 70892 72025
rect 70818 71957 70892 71991
rect 70818 71923 70838 71957
rect 70872 71923 70892 71957
rect 70818 71889 70892 71923
rect 70818 71855 70838 71889
rect 70872 71855 70892 71889
rect 70818 71821 70892 71855
rect 70818 71787 70838 71821
rect 70872 71787 70892 71821
rect 70818 71753 70892 71787
rect 70818 71719 70838 71753
rect 70872 71719 70892 71753
rect 70818 71685 70892 71719
rect 70818 71651 70838 71685
rect 70872 71651 70892 71685
rect 70818 71617 70892 71651
rect 70818 71583 70838 71617
rect 70872 71583 70892 71617
rect 70818 71549 70892 71583
rect 70818 71515 70838 71549
rect 70872 71515 70892 71549
rect 70818 71481 70892 71515
rect 70818 71447 70838 71481
rect 70872 71447 70892 71481
rect 70818 71413 70892 71447
rect 70818 71379 70838 71413
rect 70872 71379 70892 71413
rect 70818 71345 70892 71379
rect 70818 71311 70838 71345
rect 70872 71311 70892 71345
rect 70818 71277 70892 71311
rect 70818 71243 70838 71277
rect 70872 71243 70892 71277
rect 70818 71209 70892 71243
rect 70818 71175 70838 71209
rect 70872 71175 70892 71209
rect 70818 71141 70892 71175
rect 70818 71107 70838 71141
rect 70872 71107 70892 71141
rect 70818 71073 70892 71107
rect 70818 71039 70838 71073
rect 70872 71039 70892 71073
rect 70818 71005 70892 71039
rect 70818 70971 70838 71005
rect 70872 70971 70892 71005
rect 70818 70937 70892 70971
rect 70818 70903 70838 70937
rect 70872 70903 70892 70937
rect 70818 70869 70892 70903
rect 70818 70835 70838 70869
rect 70872 70835 70892 70869
rect 70818 70801 70892 70835
rect 70818 70767 70838 70801
rect 70872 70767 70892 70801
rect 70818 70733 70892 70767
rect 70818 70699 70838 70733
rect 70872 70699 70892 70733
rect 70818 70665 70892 70699
rect 70818 70631 70838 70665
rect 70872 70631 70892 70665
rect 70818 70597 70892 70631
rect 70818 70563 70838 70597
rect 70872 70563 70892 70597
rect 70818 70529 70892 70563
rect 70818 70495 70838 70529
rect 70872 70495 70892 70529
rect 70818 70461 70892 70495
rect 70818 70427 70838 70461
rect 70872 70427 70892 70461
rect 70818 70393 70892 70427
rect 70818 70359 70838 70393
rect 70872 70359 70892 70393
rect 70818 70325 70892 70359
rect 70818 70291 70838 70325
rect 70872 70291 70892 70325
rect 70818 70257 70892 70291
rect 70818 70223 70838 70257
rect 70872 70223 70892 70257
rect 70818 70189 70892 70223
rect 70818 70155 70838 70189
rect 70872 70155 70892 70189
rect 70818 70121 70892 70155
rect 70818 70087 70838 70121
rect 70872 70087 70892 70121
rect 70818 70053 70892 70087
rect 70818 70019 70838 70053
rect 70872 70019 70892 70053
rect 70818 69985 70892 70019
rect 70818 69951 70838 69985
rect 70872 69951 70892 69985
rect 70818 69917 70892 69951
rect 70818 69883 70838 69917
rect 70872 69883 70892 69917
rect 70818 69849 70892 69883
rect 70818 69815 70838 69849
rect 70872 69815 70892 69849
rect 70818 69781 70892 69815
rect 70818 69747 70838 69781
rect 70872 69747 70892 69781
rect 70818 69713 70892 69747
rect 70818 69679 70838 69713
rect 70872 69679 70892 69713
rect 70818 69645 70892 69679
rect 70818 69611 70838 69645
rect 70872 69611 70892 69645
rect 70818 69577 70892 69611
rect 70818 69543 70838 69577
rect 70872 69543 70892 69577
rect 70818 69509 70892 69543
rect 70818 69475 70838 69509
rect 70872 69475 70892 69509
rect 70818 69441 70892 69475
rect 70818 69407 70838 69441
rect 70872 69407 70892 69441
rect 70818 69373 70892 69407
rect 70818 69339 70838 69373
rect 70872 69339 70892 69373
rect 70818 69305 70892 69339
rect 70818 69271 70838 69305
rect 70872 69271 70892 69305
rect 70818 69237 70892 69271
rect 70818 69203 70838 69237
rect 70872 69203 70892 69237
rect 70818 69169 70892 69203
rect 70818 69135 70838 69169
rect 70872 69135 70892 69169
rect 70818 69101 70892 69135
rect 70818 69067 70838 69101
rect 70872 69067 70892 69101
rect 70818 69033 70892 69067
rect 70818 68999 70838 69033
rect 70872 68999 70892 69033
rect 70818 68965 70892 68999
rect 70818 68931 70838 68965
rect 70872 68931 70892 68965
rect 70818 68897 70892 68931
rect 70818 68863 70838 68897
rect 70872 68863 70892 68897
rect 70818 68829 70892 68863
rect 70818 68795 70838 68829
rect 70872 68795 70892 68829
rect 70818 68761 70892 68795
rect 70818 68727 70838 68761
rect 70872 68727 70892 68761
rect 70818 68693 70892 68727
rect 70818 68659 70838 68693
rect 70872 68659 70892 68693
rect 70818 68625 70892 68659
rect 70818 68591 70838 68625
rect 70872 68591 70892 68625
rect 70818 68557 70892 68591
rect 70818 68523 70838 68557
rect 70872 68523 70892 68557
rect 70818 68489 70892 68523
rect 70818 68455 70838 68489
rect 70872 68455 70892 68489
rect 70818 68421 70892 68455
rect 70818 68387 70838 68421
rect 70872 68387 70892 68421
rect 70818 68353 70892 68387
rect 70818 68319 70838 68353
rect 70872 68319 70892 68353
rect 70818 68285 70892 68319
rect 70818 68251 70838 68285
rect 70872 68251 70892 68285
rect 70818 68217 70892 68251
rect 70818 68183 70838 68217
rect 70872 68183 70892 68217
rect 70818 68149 70892 68183
rect 70818 68115 70838 68149
rect 70872 68115 70892 68149
rect 70818 68081 70892 68115
rect 70818 68047 70838 68081
rect 70872 68047 70892 68081
rect 70818 68013 70892 68047
rect 70818 67979 70838 68013
rect 70872 67979 70892 68013
rect 70818 67945 70892 67979
rect 70818 67911 70838 67945
rect 70872 67911 70892 67945
rect 70818 67877 70892 67911
rect 70818 67843 70838 67877
rect 70872 67843 70892 67877
rect 70818 67809 70892 67843
rect 70818 67775 70838 67809
rect 70872 67775 70892 67809
rect 70818 67741 70892 67775
rect 70818 67707 70838 67741
rect 70872 67707 70892 67741
rect 70818 67673 70892 67707
rect 70818 67639 70838 67673
rect 70872 67639 70892 67673
rect 70818 67605 70892 67639
rect 70818 67571 70838 67605
rect 70872 67571 70892 67605
rect 70818 67537 70892 67571
rect 70818 67503 70838 67537
rect 70872 67503 70892 67537
rect 70818 67469 70892 67503
rect 70818 67435 70838 67469
rect 70872 67435 70892 67469
rect 70818 67401 70892 67435
rect 70818 67367 70838 67401
rect 70872 67367 70892 67401
rect 70818 67333 70892 67367
rect 70818 67299 70838 67333
rect 70872 67299 70892 67333
rect 70818 67265 70892 67299
rect 70818 67231 70838 67265
rect 70872 67231 70892 67265
rect 70818 67197 70892 67231
rect 70818 67163 70838 67197
rect 70872 67163 70892 67197
rect 70818 67129 70892 67163
rect 70818 67095 70838 67129
rect 70872 67095 70892 67129
rect 70818 67061 70892 67095
rect 70818 67027 70838 67061
rect 70872 67027 70892 67061
rect 70818 66993 70892 67027
rect 70818 66959 70838 66993
rect 70872 66959 70892 66993
rect 70818 66925 70892 66959
rect 70818 66891 70838 66925
rect 70872 66891 70892 66925
rect 70818 66857 70892 66891
rect 70818 66823 70838 66857
rect 70872 66823 70892 66857
rect 70818 66789 70892 66823
rect 70818 66755 70838 66789
rect 70872 66755 70892 66789
rect 70818 66721 70892 66755
rect 70818 66687 70838 66721
rect 70872 66687 70892 66721
rect 70818 66653 70892 66687
rect 70818 66619 70838 66653
rect 70872 66619 70892 66653
rect 70818 66585 70892 66619
rect 70818 66551 70838 66585
rect 70872 66551 70892 66585
rect 70818 66517 70892 66551
rect 70818 66483 70838 66517
rect 70872 66483 70892 66517
rect 70818 66449 70892 66483
rect 70818 66415 70838 66449
rect 70872 66415 70892 66449
rect 70818 66381 70892 66415
rect 70818 66347 70838 66381
rect 70872 66347 70892 66381
rect 70818 66313 70892 66347
rect 70818 66279 70838 66313
rect 70872 66279 70892 66313
rect 70818 66245 70892 66279
rect 70818 66211 70838 66245
rect 70872 66211 70892 66245
rect 70818 66177 70892 66211
rect 70818 66143 70838 66177
rect 70872 66143 70892 66177
rect 70818 66109 70892 66143
rect 70818 66075 70838 66109
rect 70872 66075 70892 66109
rect 70818 66041 70892 66075
rect 70818 66007 70838 66041
rect 70872 66007 70892 66041
rect 70818 65973 70892 66007
rect 70818 65939 70838 65973
rect 70872 65939 70892 65973
rect 70818 65905 70892 65939
rect 70818 65871 70838 65905
rect 70872 65871 70892 65905
rect 70818 65837 70892 65871
rect 70818 65803 70838 65837
rect 70872 65803 70892 65837
rect 70818 65769 70892 65803
rect 70818 65735 70838 65769
rect 70872 65735 70892 65769
rect 70818 65701 70892 65735
rect 70818 65667 70838 65701
rect 70872 65667 70892 65701
rect 70818 65633 70892 65667
rect 70818 65599 70838 65633
rect 70872 65599 70892 65633
rect 70818 65565 70892 65599
rect 70818 65531 70838 65565
rect 70872 65531 70892 65565
rect 70818 65497 70892 65531
rect 70818 65463 70838 65497
rect 70872 65463 70892 65497
rect 70818 65429 70892 65463
rect 70818 65395 70838 65429
rect 70872 65395 70892 65429
rect 70818 65361 70892 65395
rect 70818 65327 70838 65361
rect 70872 65327 70892 65361
rect 70818 65293 70892 65327
rect 70818 65259 70838 65293
rect 70872 65259 70892 65293
rect 70818 65225 70892 65259
rect 70818 65191 70838 65225
rect 70872 65191 70892 65225
rect 70818 65157 70892 65191
rect 70818 65123 70838 65157
rect 70872 65123 70892 65157
rect 70818 65089 70892 65123
rect 70818 65055 70838 65089
rect 70872 65055 70892 65089
rect 70818 65021 70892 65055
rect 70818 64987 70838 65021
rect 70872 64987 70892 65021
rect 70818 64953 70892 64987
rect 70818 64919 70838 64953
rect 70872 64919 70892 64953
rect 70818 64885 70892 64919
rect 70818 64851 70838 64885
rect 70872 64851 70892 64885
rect 70818 64817 70892 64851
rect 70818 64783 70838 64817
rect 70872 64783 70892 64817
rect 70818 64749 70892 64783
rect 70818 64715 70838 64749
rect 70872 64715 70892 64749
rect 70818 64681 70892 64715
rect 70818 64647 70838 64681
rect 70872 64647 70892 64681
rect 70818 64613 70892 64647
rect 70818 64579 70838 64613
rect 70872 64579 70892 64613
rect 70818 64545 70892 64579
rect 70818 64511 70838 64545
rect 70872 64511 70892 64545
rect 70818 64477 70892 64511
rect 70818 64443 70838 64477
rect 70872 64443 70892 64477
rect 70818 64409 70892 64443
rect 70818 64375 70838 64409
rect 70872 64375 70892 64409
rect 70818 64341 70892 64375
rect 70818 64307 70838 64341
rect 70872 64307 70892 64341
rect 70818 64273 70892 64307
rect 70818 64239 70838 64273
rect 70872 64239 70892 64273
rect 70818 64205 70892 64239
rect 70818 64171 70838 64205
rect 70872 64171 70892 64205
rect 70818 64137 70892 64171
rect 70818 64103 70838 64137
rect 70872 64103 70892 64137
rect 70818 64069 70892 64103
rect 70818 64035 70838 64069
rect 70872 64035 70892 64069
rect 70818 64001 70892 64035
rect 70818 63967 70838 64001
rect 70872 63967 70892 64001
rect 70818 63933 70892 63967
rect 70818 63899 70838 63933
rect 70872 63899 70892 63933
rect 70818 63865 70892 63899
rect 70818 63831 70838 63865
rect 70872 63831 70892 63865
rect 70818 63797 70892 63831
rect 70818 63763 70838 63797
rect 70872 63763 70892 63797
rect 70818 63729 70892 63763
rect 70818 63695 70838 63729
rect 70872 63695 70892 63729
rect 70818 63661 70892 63695
rect 70818 63627 70838 63661
rect 70872 63627 70892 63661
rect 70818 63593 70892 63627
rect 70818 63559 70838 63593
rect 70872 63559 70892 63593
rect 70818 63525 70892 63559
rect 70818 63491 70838 63525
rect 70872 63491 70892 63525
rect 70818 63457 70892 63491
rect 70818 63423 70838 63457
rect 70872 63423 70892 63457
rect 70818 63389 70892 63423
rect 70818 63355 70838 63389
rect 70872 63355 70892 63389
rect 70818 63321 70892 63355
rect 70818 63287 70838 63321
rect 70872 63287 70892 63321
rect 70818 63253 70892 63287
rect 70818 63219 70838 63253
rect 70872 63219 70892 63253
rect 70818 63185 70892 63219
rect 70818 63151 70838 63185
rect 70872 63151 70892 63185
rect 70818 63117 70892 63151
rect 70818 63083 70838 63117
rect 70872 63083 70892 63117
rect 70818 63049 70892 63083
rect 70818 63015 70838 63049
rect 70872 63015 70892 63049
rect 70818 62981 70892 63015
rect 70818 62947 70838 62981
rect 70872 62947 70892 62981
rect 70818 62913 70892 62947
rect 70818 62879 70838 62913
rect 70872 62879 70892 62913
rect 70818 62845 70892 62879
rect 70818 62811 70838 62845
rect 70872 62811 70892 62845
rect 70818 62777 70892 62811
rect 70818 62743 70838 62777
rect 70872 62743 70892 62777
rect 70818 62709 70892 62743
rect 70818 62675 70838 62709
rect 70872 62675 70892 62709
rect 70818 62641 70892 62675
rect 70818 62607 70838 62641
rect 70872 62607 70892 62641
rect 70818 62573 70892 62607
rect 70818 62539 70838 62573
rect 70872 62539 70892 62573
rect 70818 62505 70892 62539
rect 70818 62471 70838 62505
rect 70872 62471 70892 62505
rect 70818 62437 70892 62471
rect 70818 62403 70838 62437
rect 70872 62403 70892 62437
rect 70818 62369 70892 62403
rect 70818 62335 70838 62369
rect 70872 62335 70892 62369
rect 70818 62301 70892 62335
rect 70818 62267 70838 62301
rect 70872 62267 70892 62301
rect 70818 62233 70892 62267
rect 70818 62199 70838 62233
rect 70872 62199 70892 62233
rect 70818 62165 70892 62199
rect 70818 62131 70838 62165
rect 70872 62131 70892 62165
rect 70818 62097 70892 62131
rect 70818 62063 70838 62097
rect 70872 62063 70892 62097
rect 70818 62029 70892 62063
rect 70818 61995 70838 62029
rect 70872 61995 70892 62029
rect 70818 61961 70892 61995
rect 70818 61927 70838 61961
rect 70872 61927 70892 61961
rect 70818 61893 70892 61927
rect 70818 61859 70838 61893
rect 70872 61859 70892 61893
rect 70818 61825 70892 61859
rect 70818 61791 70838 61825
rect 70872 61791 70892 61825
rect 70818 61757 70892 61791
rect 70818 61723 70838 61757
rect 70872 61723 70892 61757
rect 70818 61689 70892 61723
rect 70818 61655 70838 61689
rect 70872 61655 70892 61689
rect 70818 61621 70892 61655
rect 70818 61587 70838 61621
rect 70872 61587 70892 61621
rect 70818 61553 70892 61587
rect 70818 61519 70838 61553
rect 70872 61519 70892 61553
rect 70818 61485 70892 61519
rect 70818 61451 70838 61485
rect 70872 61451 70892 61485
rect 70818 61417 70892 61451
rect 70818 61383 70838 61417
rect 70872 61383 70892 61417
rect 70818 61349 70892 61383
rect 70818 61315 70838 61349
rect 70872 61315 70892 61349
rect 70818 61281 70892 61315
rect 70818 61247 70838 61281
rect 70872 61247 70892 61281
rect 70818 61213 70892 61247
rect 70818 61179 70838 61213
rect 70872 61179 70892 61213
rect 70818 61145 70892 61179
rect 70818 61111 70838 61145
rect 70872 61111 70892 61145
rect 70818 61077 70892 61111
rect 70818 61043 70838 61077
rect 70872 61043 70892 61077
rect 70818 61009 70892 61043
rect 70818 60975 70838 61009
rect 70872 60975 70892 61009
rect 70818 60941 70892 60975
rect 70818 60907 70838 60941
rect 70872 60907 70892 60941
rect 70818 60873 70892 60907
rect 70818 60839 70838 60873
rect 70872 60839 70892 60873
rect 70818 60805 70892 60839
rect 70818 60771 70838 60805
rect 70872 60771 70892 60805
rect 70818 60737 70892 60771
rect 70818 60703 70838 60737
rect 70872 60703 70892 60737
rect 70818 60669 70892 60703
rect 70818 60635 70838 60669
rect 70872 60635 70892 60669
rect 70818 60601 70892 60635
rect 70818 60567 70838 60601
rect 70872 60567 70892 60601
rect 70818 60533 70892 60567
rect 70818 60499 70838 60533
rect 70872 60499 70892 60533
rect 70818 60465 70892 60499
rect 70818 60431 70838 60465
rect 70872 60431 70892 60465
rect 70818 60397 70892 60431
rect 70818 60363 70838 60397
rect 70872 60363 70892 60397
rect 70818 60329 70892 60363
rect 70818 60295 70838 60329
rect 70872 60295 70892 60329
rect 70818 60261 70892 60295
rect 70818 60227 70838 60261
rect 70872 60227 70892 60261
rect 70818 60193 70892 60227
rect 70818 60159 70838 60193
rect 70872 60159 70892 60193
rect 70818 60125 70892 60159
rect 70818 60091 70838 60125
rect 70872 60091 70892 60125
rect 70818 60057 70892 60091
rect 70818 60023 70838 60057
rect 70872 60023 70892 60057
rect 70818 59989 70892 60023
rect 70818 59955 70838 59989
rect 70872 59955 70892 59989
rect 70818 59921 70892 59955
rect 70818 59887 70838 59921
rect 70872 59887 70892 59921
rect 70818 59853 70892 59887
rect 70818 59819 70838 59853
rect 70872 59819 70892 59853
rect 70818 59785 70892 59819
rect 70818 59751 70838 59785
rect 70872 59751 70892 59785
rect 70818 59717 70892 59751
rect 70818 59683 70838 59717
rect 70872 59683 70892 59717
rect 70818 59649 70892 59683
rect 70818 59615 70838 59649
rect 70872 59615 70892 59649
rect 70818 59581 70892 59615
rect 70818 59547 70838 59581
rect 70872 59547 70892 59581
rect 70818 59513 70892 59547
rect 70818 59479 70838 59513
rect 70872 59479 70892 59513
rect 70818 59445 70892 59479
rect 70818 59411 70838 59445
rect 70872 59411 70892 59445
rect 70818 59377 70892 59411
rect 70818 59343 70838 59377
rect 70872 59343 70892 59377
rect 70818 59309 70892 59343
rect 70818 59275 70838 59309
rect 70872 59275 70892 59309
rect 70818 59241 70892 59275
rect 70818 59207 70838 59241
rect 70872 59207 70892 59241
rect 70818 59173 70892 59207
rect 70818 59139 70838 59173
rect 70872 59139 70892 59173
rect 70818 59105 70892 59139
rect 70818 59071 70838 59105
rect 70872 59071 70892 59105
rect 70818 59037 70892 59071
rect 70818 59003 70838 59037
rect 70872 59003 70892 59037
rect 70818 58969 70892 59003
rect 70818 58935 70838 58969
rect 70872 58935 70892 58969
rect 70818 58901 70892 58935
rect 70818 58867 70838 58901
rect 70872 58867 70892 58901
rect 70818 58833 70892 58867
rect 70818 58799 70838 58833
rect 70872 58799 70892 58833
rect 70818 58765 70892 58799
rect 70818 58731 70838 58765
rect 70872 58731 70892 58765
rect 70818 58697 70892 58731
rect 70818 58663 70838 58697
rect 70872 58663 70892 58697
rect 70818 58629 70892 58663
rect 70818 58595 70838 58629
rect 70872 58595 70892 58629
rect 70818 58561 70892 58595
rect 70818 58527 70838 58561
rect 70872 58527 70892 58561
rect 70818 58493 70892 58527
rect 70818 58459 70838 58493
rect 70872 58459 70892 58493
rect 70818 58425 70892 58459
rect 70818 58391 70838 58425
rect 70872 58391 70892 58425
rect 70818 58357 70892 58391
rect 70818 58323 70838 58357
rect 70872 58323 70892 58357
rect 70818 58289 70892 58323
rect 70818 58255 70838 58289
rect 70872 58255 70892 58289
rect 70818 58221 70892 58255
rect 70818 58187 70838 58221
rect 70872 58187 70892 58221
rect 70818 58153 70892 58187
rect 70818 58119 70838 58153
rect 70872 58119 70892 58153
rect 70818 58085 70892 58119
rect 70818 58051 70838 58085
rect 70872 58051 70892 58085
rect 70818 58017 70892 58051
rect 70818 57983 70838 58017
rect 70872 57983 70892 58017
rect 70818 57949 70892 57983
rect 70818 57915 70838 57949
rect 70872 57915 70892 57949
rect 70818 57881 70892 57915
rect 70818 57847 70838 57881
rect 70872 57847 70892 57881
rect 70818 57813 70892 57847
rect 70818 57779 70838 57813
rect 70872 57779 70892 57813
rect 70818 57745 70892 57779
rect 70818 57711 70838 57745
rect 70872 57711 70892 57745
rect 70818 57677 70892 57711
rect 70818 57643 70838 57677
rect 70872 57643 70892 57677
rect 70818 57609 70892 57643
rect 70818 57575 70838 57609
rect 70872 57575 70892 57609
rect 70818 57541 70892 57575
rect 70818 57507 70838 57541
rect 70872 57507 70892 57541
rect 70818 57473 70892 57507
rect 70818 57439 70838 57473
rect 70872 57439 70892 57473
rect 70818 57405 70892 57439
rect 70818 57371 70838 57405
rect 70872 57371 70892 57405
rect 70818 57337 70892 57371
rect 70818 57303 70838 57337
rect 70872 57303 70892 57337
rect 70818 57269 70892 57303
rect 70818 57235 70838 57269
rect 70872 57235 70892 57269
rect 70818 57201 70892 57235
rect 70818 57167 70838 57201
rect 70872 57167 70892 57201
rect 70818 57133 70892 57167
rect 70818 57099 70838 57133
rect 70872 57099 70892 57133
rect 70818 57065 70892 57099
rect 70818 57031 70838 57065
rect 70872 57031 70892 57065
rect 70818 56997 70892 57031
rect 70818 56963 70838 56997
rect 70872 56963 70892 56997
rect 70818 56929 70892 56963
rect 70818 56895 70838 56929
rect 70872 56895 70892 56929
rect 70818 56861 70892 56895
rect 70818 56827 70838 56861
rect 70872 56827 70892 56861
rect 70818 56793 70892 56827
rect 70818 56759 70838 56793
rect 70872 56759 70892 56793
rect 70818 56725 70892 56759
rect 70818 56691 70838 56725
rect 70872 56691 70892 56725
rect 70818 56657 70892 56691
rect 70818 56623 70838 56657
rect 70872 56623 70892 56657
rect 70818 56589 70892 56623
rect 70818 56555 70838 56589
rect 70872 56555 70892 56589
rect 70818 56521 70892 56555
rect 70818 56487 70838 56521
rect 70872 56487 70892 56521
rect 70818 56453 70892 56487
rect 70818 56419 70838 56453
rect 70872 56419 70892 56453
rect 70818 56385 70892 56419
rect 70818 56351 70838 56385
rect 70872 56351 70892 56385
rect 70818 56317 70892 56351
rect 70818 56283 70838 56317
rect 70872 56283 70892 56317
rect 70818 56249 70892 56283
rect 70818 56215 70838 56249
rect 70872 56215 70892 56249
rect 70818 56181 70892 56215
rect 70818 56147 70838 56181
rect 70872 56147 70892 56181
rect 70818 56113 70892 56147
rect 70818 56079 70838 56113
rect 70872 56079 70892 56113
rect 70818 56045 70892 56079
rect 70818 56011 70838 56045
rect 70872 56011 70892 56045
rect 70818 55977 70892 56011
rect 70818 55943 70838 55977
rect 70872 55943 70892 55977
rect 70818 55909 70892 55943
rect 70818 55875 70838 55909
rect 70872 55875 70892 55909
rect 70818 55841 70892 55875
rect 70818 55807 70838 55841
rect 70872 55807 70892 55841
rect 70818 55773 70892 55807
rect 70818 55739 70838 55773
rect 70872 55739 70892 55773
rect 70818 55705 70892 55739
rect 70818 55671 70838 55705
rect 70872 55671 70892 55705
rect 70818 55637 70892 55671
rect 70818 55603 70838 55637
rect 70872 55603 70892 55637
rect 70818 55569 70892 55603
rect 70818 55535 70838 55569
rect 70872 55535 70892 55569
rect 70818 55501 70892 55535
rect 70818 55467 70838 55501
rect 70872 55467 70892 55501
rect 70818 55433 70892 55467
rect 70818 55399 70838 55433
rect 70872 55399 70892 55433
rect 70818 55365 70892 55399
rect 70818 55331 70838 55365
rect 70872 55331 70892 55365
rect 70818 55297 70892 55331
rect 70818 55263 70838 55297
rect 70872 55263 70892 55297
rect 70818 55229 70892 55263
rect 70818 55195 70838 55229
rect 70872 55195 70892 55229
rect 70818 55161 70892 55195
rect 70818 55127 70838 55161
rect 70872 55127 70892 55161
rect 70818 55093 70892 55127
rect 70818 55059 70838 55093
rect 70872 55059 70892 55093
rect 70818 55025 70892 55059
rect 70818 54991 70838 55025
rect 70872 54991 70892 55025
rect 70818 54957 70892 54991
rect 70818 54923 70838 54957
rect 70872 54923 70892 54957
rect 70818 54889 70892 54923
rect 70818 54855 70838 54889
rect 70872 54855 70892 54889
rect 70818 54821 70892 54855
rect 70818 54787 70838 54821
rect 70872 54787 70892 54821
rect 70818 54753 70892 54787
rect 70818 54719 70838 54753
rect 70872 54719 70892 54753
rect 70818 54685 70892 54719
rect 70818 54651 70838 54685
rect 70872 54651 70892 54685
rect 70818 54617 70892 54651
rect 70818 54583 70838 54617
rect 70872 54583 70892 54617
rect 70818 54549 70892 54583
rect 70818 54515 70838 54549
rect 70872 54515 70892 54549
rect 70818 54481 70892 54515
rect 70818 54447 70838 54481
rect 70872 54447 70892 54481
rect 70818 54413 70892 54447
rect 70818 54379 70838 54413
rect 70872 54379 70892 54413
rect 70818 54345 70892 54379
rect 70818 54311 70838 54345
rect 70872 54311 70892 54345
rect 70818 54277 70892 54311
rect 70818 54243 70838 54277
rect 70872 54243 70892 54277
rect 70818 54209 70892 54243
rect 70818 54175 70838 54209
rect 70872 54175 70892 54209
rect 70818 54141 70892 54175
rect 70818 54107 70838 54141
rect 70872 54107 70892 54141
rect 70818 54073 70892 54107
rect 70818 54039 70838 54073
rect 70872 54039 70892 54073
rect 70818 54005 70892 54039
rect 70818 53971 70838 54005
rect 70872 53971 70892 54005
rect 70818 53937 70892 53971
rect 70818 53903 70838 53937
rect 70872 53903 70892 53937
rect 70818 53869 70892 53903
rect 70818 53835 70838 53869
rect 70872 53835 70892 53869
rect 70818 53801 70892 53835
rect 70818 53767 70838 53801
rect 70872 53767 70892 53801
rect 70818 53733 70892 53767
rect 70818 53699 70838 53733
rect 70872 53699 70892 53733
rect 70818 53665 70892 53699
rect 70818 53631 70838 53665
rect 70872 53631 70892 53665
rect 70818 53597 70892 53631
rect 70818 53563 70838 53597
rect 70872 53563 70892 53597
rect 70818 53529 70892 53563
rect 70818 53495 70838 53529
rect 70872 53495 70892 53529
rect 70818 53461 70892 53495
rect 70818 53427 70838 53461
rect 70872 53427 70892 53461
rect 70818 53393 70892 53427
rect 70818 53359 70838 53393
rect 70872 53359 70892 53393
rect 70818 53325 70892 53359
rect 70818 53291 70838 53325
rect 70872 53291 70892 53325
rect 70818 53257 70892 53291
rect 70818 53223 70838 53257
rect 70872 53223 70892 53257
rect 70818 53189 70892 53223
rect 70818 53155 70838 53189
rect 70872 53155 70892 53189
rect 70818 53121 70892 53155
rect 70818 53087 70838 53121
rect 70872 53087 70892 53121
rect 70818 53053 70892 53087
rect 70818 53019 70838 53053
rect 70872 53019 70892 53053
rect 70818 52985 70892 53019
rect 70818 52951 70838 52985
rect 70872 52951 70892 52985
rect 70818 52917 70892 52951
rect 70818 52883 70838 52917
rect 70872 52883 70892 52917
rect 70818 52849 70892 52883
rect 70818 52815 70838 52849
rect 70872 52815 70892 52849
rect 70818 52781 70892 52815
rect 70818 52747 70838 52781
rect 70872 52747 70892 52781
rect 70818 52713 70892 52747
rect 70818 52679 70838 52713
rect 70872 52679 70892 52713
rect 70818 52645 70892 52679
rect 70818 52611 70838 52645
rect 70872 52611 70892 52645
rect 70818 52577 70892 52611
rect 70818 52543 70838 52577
rect 70872 52543 70892 52577
rect 70818 52509 70892 52543
rect 70818 52475 70838 52509
rect 70872 52475 70892 52509
rect 70818 52441 70892 52475
rect 70818 52407 70838 52441
rect 70872 52407 70892 52441
rect 70818 52373 70892 52407
rect 70818 52339 70838 52373
rect 70872 52339 70892 52373
rect 70818 52305 70892 52339
rect 70818 52271 70838 52305
rect 70872 52271 70892 52305
rect 70818 52237 70892 52271
rect 70818 52203 70838 52237
rect 70872 52203 70892 52237
rect 70818 52169 70892 52203
rect 70818 52135 70838 52169
rect 70872 52135 70892 52169
rect 70818 52101 70892 52135
rect 70818 52067 70838 52101
rect 70872 52067 70892 52101
rect 70818 52033 70892 52067
rect 70818 51999 70838 52033
rect 70872 51999 70892 52033
rect 70818 51965 70892 51999
rect 70818 51931 70838 51965
rect 70872 51931 70892 51965
rect 70818 51897 70892 51931
rect 70818 51863 70838 51897
rect 70872 51863 70892 51897
rect 70818 51829 70892 51863
rect 70818 51795 70838 51829
rect 70872 51795 70892 51829
rect 70818 51761 70892 51795
rect 70818 51727 70838 51761
rect 70872 51727 70892 51761
rect 70818 51693 70892 51727
rect 70818 51659 70838 51693
rect 70872 51659 70892 51693
rect 70818 51625 70892 51659
rect 70818 51591 70838 51625
rect 70872 51591 70892 51625
rect 70818 51557 70892 51591
rect 70818 51523 70838 51557
rect 70872 51523 70892 51557
rect 70818 51489 70892 51523
rect 70818 51455 70838 51489
rect 70872 51455 70892 51489
rect 70818 51421 70892 51455
rect 70818 51387 70838 51421
rect 70872 51387 70892 51421
rect 70818 51353 70892 51387
rect 70818 51319 70838 51353
rect 70872 51319 70892 51353
rect 70818 51285 70892 51319
rect 70818 51251 70838 51285
rect 70872 51251 70892 51285
rect 70818 51217 70892 51251
rect 70818 51183 70838 51217
rect 70872 51183 70892 51217
rect 70818 51149 70892 51183
rect 70818 51115 70838 51149
rect 70872 51115 70892 51149
rect 70818 51081 70892 51115
rect 70818 51047 70838 51081
rect 70872 51047 70892 51081
rect 70818 51013 70892 51047
rect 70818 50979 70838 51013
rect 70872 50979 70892 51013
rect 70818 50945 70892 50979
rect 70818 50911 70838 50945
rect 70872 50911 70892 50945
rect 70818 50877 70892 50911
rect 70818 50843 70838 50877
rect 70872 50843 70892 50877
rect 70818 50809 70892 50843
rect 70818 50775 70838 50809
rect 70872 50775 70892 50809
rect 70818 50741 70892 50775
rect 70818 50707 70838 50741
rect 70872 50707 70892 50741
rect 70818 50673 70892 50707
rect 70818 50639 70838 50673
rect 70872 50639 70892 50673
rect 70818 50605 70892 50639
rect 70818 50571 70838 50605
rect 70872 50571 70892 50605
rect 70818 50537 70892 50571
rect 70818 50503 70838 50537
rect 70872 50503 70892 50537
rect 70818 50469 70892 50503
rect 70818 50435 70838 50469
rect 70872 50435 70892 50469
rect 70818 50401 70892 50435
rect 70818 50367 70838 50401
rect 70872 50367 70892 50401
rect 70818 50333 70892 50367
rect 70818 50299 70838 50333
rect 70872 50299 70892 50333
rect 70818 50265 70892 50299
rect 70818 50231 70838 50265
rect 70872 50231 70892 50265
rect 70818 50197 70892 50231
rect 70818 50163 70838 50197
rect 70872 50163 70892 50197
rect 70818 50129 70892 50163
rect 70818 50095 70838 50129
rect 70872 50095 70892 50129
rect 70818 50061 70892 50095
rect 70818 50027 70838 50061
rect 70872 50027 70892 50061
rect 70818 49993 70892 50027
rect 70818 49959 70838 49993
rect 70872 49959 70892 49993
rect 70818 49925 70892 49959
rect 70818 49891 70838 49925
rect 70872 49891 70892 49925
rect 70818 49857 70892 49891
rect 70818 49823 70838 49857
rect 70872 49823 70892 49857
rect 70818 49789 70892 49823
rect 70818 49755 70838 49789
rect 70872 49755 70892 49789
rect 70818 49721 70892 49755
rect 70818 49687 70838 49721
rect 70872 49687 70892 49721
rect 70818 49653 70892 49687
rect 70818 49619 70838 49653
rect 70872 49619 70892 49653
rect 70818 49585 70892 49619
rect 70818 49551 70838 49585
rect 70872 49551 70892 49585
rect 70818 49517 70892 49551
rect 70818 49483 70838 49517
rect 70872 49483 70892 49517
rect 70818 49449 70892 49483
rect 70818 49415 70838 49449
rect 70872 49415 70892 49449
rect 70818 49381 70892 49415
rect 70818 49347 70838 49381
rect 70872 49347 70892 49381
rect 70818 49313 70892 49347
rect 70818 49279 70838 49313
rect 70872 49279 70892 49313
rect 70818 49245 70892 49279
rect 70818 49211 70838 49245
rect 70872 49211 70892 49245
rect 70818 49177 70892 49211
rect 70818 49143 70838 49177
rect 70872 49143 70892 49177
rect 70818 49109 70892 49143
rect 70818 49075 70838 49109
rect 70872 49075 70892 49109
rect 70818 49041 70892 49075
rect 70818 49007 70838 49041
rect 70872 49007 70892 49041
rect 70818 48973 70892 49007
rect 70818 48939 70838 48973
rect 70872 48939 70892 48973
rect 70818 48905 70892 48939
rect 70818 48871 70838 48905
rect 70872 48871 70892 48905
rect 70818 48837 70892 48871
rect 70818 48803 70838 48837
rect 70872 48803 70892 48837
rect 70818 48769 70892 48803
rect 70818 48735 70838 48769
rect 70872 48735 70892 48769
rect 70818 48701 70892 48735
rect 70818 48667 70838 48701
rect 70872 48667 70892 48701
rect 70818 48633 70892 48667
rect 70818 48599 70838 48633
rect 70872 48599 70892 48633
rect 70818 48565 70892 48599
rect 70818 48531 70838 48565
rect 70872 48531 70892 48565
rect 70818 48497 70892 48531
rect 70818 48463 70838 48497
rect 70872 48463 70892 48497
rect 70818 48429 70892 48463
rect 70818 48395 70838 48429
rect 70872 48395 70892 48429
rect 70818 48361 70892 48395
rect 70818 48327 70838 48361
rect 70872 48327 70892 48361
rect 70818 48293 70892 48327
rect 70818 48259 70838 48293
rect 70872 48259 70892 48293
rect 70818 48225 70892 48259
rect 70818 48191 70838 48225
rect 70872 48191 70892 48225
rect 70818 48157 70892 48191
rect 70818 48123 70838 48157
rect 70872 48123 70892 48157
rect 70818 48089 70892 48123
rect 70818 48055 70838 48089
rect 70872 48055 70892 48089
rect 70818 48021 70892 48055
rect 70818 47987 70838 48021
rect 70872 47987 70892 48021
rect 70818 47953 70892 47987
rect 70818 47919 70838 47953
rect 70872 47919 70892 47953
rect 70818 47885 70892 47919
rect 70818 47851 70838 47885
rect 70872 47851 70892 47885
rect 70818 47817 70892 47851
rect 70818 47783 70838 47817
rect 70872 47783 70892 47817
rect 70818 47749 70892 47783
rect 70818 47715 70838 47749
rect 70872 47715 70892 47749
rect 70818 47681 70892 47715
rect 70818 47647 70838 47681
rect 70872 47647 70892 47681
rect 70818 47613 70892 47647
rect 70818 47579 70838 47613
rect 70872 47579 70892 47613
rect 70818 47545 70892 47579
rect 70818 47511 70838 47545
rect 70872 47511 70892 47545
rect 70818 47477 70892 47511
rect 70818 47443 70838 47477
rect 70872 47443 70892 47477
rect 70818 47409 70892 47443
rect 70818 47375 70838 47409
rect 70872 47375 70892 47409
rect 70818 47341 70892 47375
rect 70818 47307 70838 47341
rect 70872 47307 70892 47341
rect 70818 47273 70892 47307
rect 70818 47239 70838 47273
rect 70872 47239 70892 47273
rect 70818 47205 70892 47239
rect 70818 47171 70838 47205
rect 70872 47171 70892 47205
rect 70818 47137 70892 47171
rect 70818 47103 70838 47137
rect 70872 47103 70892 47137
rect 70818 47069 70892 47103
rect 70818 47035 70838 47069
rect 70872 47035 70892 47069
rect 70818 47001 70892 47035
rect 70818 46967 70838 47001
rect 70872 46967 70892 47001
rect 70818 46933 70892 46967
rect 70818 46899 70838 46933
rect 70872 46899 70892 46933
rect 70818 46865 70892 46899
rect 70818 46831 70838 46865
rect 70872 46831 70892 46865
rect 70818 46797 70892 46831
rect 70818 46763 70838 46797
rect 70872 46763 70892 46797
rect 70818 46729 70892 46763
rect 70818 46695 70838 46729
rect 70872 46695 70892 46729
rect 70818 46661 70892 46695
rect 70818 46627 70838 46661
rect 70872 46627 70892 46661
rect 70818 46593 70892 46627
rect 70818 46559 70838 46593
rect 70872 46559 70892 46593
rect 70818 46525 70892 46559
rect 70818 46491 70838 46525
rect 70872 46491 70892 46525
rect 70818 46457 70892 46491
rect 70818 46423 70838 46457
rect 70872 46423 70892 46457
rect 70818 46389 70892 46423
rect 70818 46355 70838 46389
rect 70872 46355 70892 46389
rect 70818 46321 70892 46355
rect 70818 46287 70838 46321
rect 70872 46287 70892 46321
rect 70818 46253 70892 46287
rect 70818 46219 70838 46253
rect 70872 46219 70892 46253
rect 70818 46185 70892 46219
rect 70818 46151 70838 46185
rect 70872 46151 70892 46185
rect 70818 46117 70892 46151
rect 70818 46083 70838 46117
rect 70872 46083 70892 46117
rect 70818 46049 70892 46083
rect 70818 46015 70838 46049
rect 70872 46015 70892 46049
rect 70818 45981 70892 46015
rect 70818 45947 70838 45981
rect 70872 45947 70892 45981
rect 70818 45940 70892 45947
rect 59084 45920 70892 45940
rect 59084 45886 59191 45920
rect 59225 45886 59259 45920
rect 59293 45886 59327 45920
rect 59361 45886 59395 45920
rect 59429 45886 59463 45920
rect 59497 45886 59531 45920
rect 59565 45886 59599 45920
rect 59633 45886 59667 45920
rect 59701 45886 59735 45920
rect 59769 45886 59803 45920
rect 59837 45886 59871 45920
rect 59905 45886 59939 45920
rect 59973 45886 60007 45920
rect 60041 45886 60075 45920
rect 60109 45886 60143 45920
rect 60177 45886 60211 45920
rect 60245 45886 60279 45920
rect 60313 45886 60347 45920
rect 60381 45886 60415 45920
rect 60449 45886 60483 45920
rect 60517 45886 60551 45920
rect 60585 45886 60619 45920
rect 60653 45886 60687 45920
rect 60721 45886 60755 45920
rect 60789 45886 60823 45920
rect 60857 45886 60891 45920
rect 60925 45886 60959 45920
rect 60993 45886 61027 45920
rect 61061 45886 61095 45920
rect 61129 45886 61163 45920
rect 61197 45886 61231 45920
rect 61265 45886 61299 45920
rect 61333 45886 61367 45920
rect 61401 45886 61435 45920
rect 61469 45886 61503 45920
rect 61537 45886 61571 45920
rect 61605 45886 61639 45920
rect 61673 45886 61707 45920
rect 61741 45886 61775 45920
rect 61809 45886 61843 45920
rect 61877 45886 61911 45920
rect 61945 45886 61979 45920
rect 62013 45886 62047 45920
rect 62081 45886 62115 45920
rect 62149 45886 62183 45920
rect 62217 45886 62251 45920
rect 62285 45886 62319 45920
rect 62353 45886 62387 45920
rect 62421 45886 62455 45920
rect 62489 45886 62523 45920
rect 62557 45886 62591 45920
rect 62625 45886 62659 45920
rect 62693 45886 62727 45920
rect 62761 45886 62795 45920
rect 62829 45886 62863 45920
rect 62897 45886 62931 45920
rect 62965 45886 62999 45920
rect 63033 45886 63067 45920
rect 63101 45886 63135 45920
rect 63169 45886 63203 45920
rect 63237 45886 63271 45920
rect 63305 45886 63339 45920
rect 63373 45886 63407 45920
rect 63441 45886 63475 45920
rect 63509 45886 63543 45920
rect 63577 45886 63611 45920
rect 63645 45886 63679 45920
rect 63713 45886 63747 45920
rect 63781 45886 63815 45920
rect 63849 45886 63883 45920
rect 63917 45886 63951 45920
rect 63985 45886 64019 45920
rect 64053 45886 64087 45920
rect 64121 45886 64155 45920
rect 64189 45886 64223 45920
rect 64257 45886 64291 45920
rect 64325 45886 64359 45920
rect 64393 45886 64427 45920
rect 64461 45886 64495 45920
rect 64529 45886 64563 45920
rect 64597 45886 64631 45920
rect 64665 45886 64699 45920
rect 64733 45886 64767 45920
rect 64801 45886 64835 45920
rect 64869 45886 64903 45920
rect 64937 45886 64971 45920
rect 65005 45886 65039 45920
rect 65073 45886 65107 45920
rect 65141 45886 65175 45920
rect 65209 45886 65243 45920
rect 65277 45886 65311 45920
rect 65345 45886 65379 45920
rect 65413 45886 65447 45920
rect 65481 45886 65515 45920
rect 65549 45886 65583 45920
rect 65617 45886 65651 45920
rect 65685 45886 65719 45920
rect 65753 45886 65787 45920
rect 65821 45886 65855 45920
rect 65889 45886 65923 45920
rect 65957 45886 65991 45920
rect 66025 45886 66059 45920
rect 66093 45886 66127 45920
rect 66161 45886 66195 45920
rect 66229 45886 66263 45920
rect 66297 45886 66331 45920
rect 66365 45886 66399 45920
rect 66433 45886 66467 45920
rect 66501 45886 66535 45920
rect 66569 45886 66603 45920
rect 66637 45886 66671 45920
rect 66705 45886 66739 45920
rect 66773 45886 66807 45920
rect 66841 45886 66875 45920
rect 66909 45886 66943 45920
rect 66977 45886 67011 45920
rect 67045 45886 67079 45920
rect 67113 45886 67147 45920
rect 67181 45886 67215 45920
rect 67249 45886 67283 45920
rect 67317 45886 67351 45920
rect 67385 45886 67419 45920
rect 67453 45886 67487 45920
rect 67521 45886 67555 45920
rect 67589 45886 67623 45920
rect 67657 45886 67691 45920
rect 67725 45886 67759 45920
rect 67793 45886 67827 45920
rect 67861 45886 67895 45920
rect 67929 45886 67963 45920
rect 67997 45886 68031 45920
rect 68065 45886 68099 45920
rect 68133 45886 68167 45920
rect 68201 45886 68235 45920
rect 68269 45886 68303 45920
rect 68337 45886 68371 45920
rect 68405 45886 68439 45920
rect 68473 45886 68507 45920
rect 68541 45886 68575 45920
rect 68609 45886 68643 45920
rect 68677 45886 68711 45920
rect 68745 45886 68779 45920
rect 68813 45886 68847 45920
rect 68881 45886 68915 45920
rect 68949 45886 68983 45920
rect 69017 45886 69051 45920
rect 69085 45886 69119 45920
rect 69153 45886 69187 45920
rect 69221 45886 69255 45920
rect 69289 45886 69323 45920
rect 69357 45886 69391 45920
rect 69425 45886 69459 45920
rect 69493 45886 69527 45920
rect 69561 45886 69595 45920
rect 69629 45886 69663 45920
rect 69697 45886 69731 45920
rect 69765 45886 69799 45920
rect 69833 45886 69867 45920
rect 69901 45886 69935 45920
rect 69969 45886 70003 45920
rect 70037 45886 70071 45920
rect 70105 45886 70139 45920
rect 70173 45886 70207 45920
rect 70241 45886 70275 45920
rect 70309 45886 70343 45920
rect 70377 45886 70411 45920
rect 70445 45886 70479 45920
rect 70513 45886 70547 45920
rect 70581 45886 70615 45920
rect 70649 45886 70683 45920
rect 70717 45886 70751 45920
rect 70785 45886 70892 45920
rect 59084 45866 70892 45886
rect -3738 45830 -3718 45864
rect -3684 45830 -3664 45864
rect -3738 45796 -3664 45830
rect -3738 45762 -3718 45796
rect -3684 45762 -3664 45796
rect -3738 45728 -3664 45762
rect -3738 45694 -3718 45728
rect -3684 45694 -3664 45728
rect -3738 45660 -3664 45694
rect -3738 45626 -3718 45660
rect -3684 45626 -3664 45660
rect -3738 45592 -3664 45626
rect -3738 45558 -3718 45592
rect -3684 45558 -3664 45592
rect -3738 45524 -3664 45558
rect -3738 45490 -3718 45524
rect -3684 45490 -3664 45524
rect -3738 45456 -3664 45490
rect -3738 45422 -3718 45456
rect -3684 45422 -3664 45456
rect -3738 45388 -3664 45422
rect -3738 45354 -3718 45388
rect -3684 45354 -3664 45388
rect -3738 45320 -3664 45354
rect -3738 45286 -3718 45320
rect -3684 45286 -3664 45320
rect -3738 45252 -3664 45286
rect -3738 45218 -3718 45252
rect -3684 45218 -3664 45252
rect -3738 45184 -3664 45218
rect -3738 45150 -3718 45184
rect -3684 45150 -3664 45184
rect -3738 45116 -3664 45150
rect -3738 45082 -3718 45116
rect -3684 45082 -3664 45116
rect -3738 45048 -3664 45082
rect -3738 45014 -3718 45048
rect -3684 45014 -3664 45048
rect -3738 44980 -3664 45014
rect -3738 44946 -3718 44980
rect -3684 44946 -3664 44980
rect -3738 44912 -3664 44946
rect -3738 44878 -3718 44912
rect -3684 44878 -3664 44912
rect -3738 44844 -3664 44878
rect -3738 44810 -3718 44844
rect -3684 44810 -3664 44844
rect -3738 44776 -3664 44810
rect -3738 44742 -3718 44776
rect -3684 44742 -3664 44776
rect -3738 44708 -3664 44742
rect -3738 44674 -3718 44708
rect -3684 44674 -3664 44708
rect -3738 44640 -3664 44674
rect -3738 44606 -3718 44640
rect -3684 44606 -3664 44640
rect -3738 44572 -3664 44606
rect -3738 44538 -3718 44572
rect -3684 44538 -3664 44572
rect -3738 44504 -3664 44538
rect -3738 44470 -3718 44504
rect -3684 44470 -3664 44504
rect -3738 44436 -3664 44470
rect -3738 44402 -3718 44436
rect -3684 44402 -3664 44436
rect -3738 44368 -3664 44402
rect -3738 44334 -3718 44368
rect -3684 44334 -3664 44368
rect -3738 44300 -3664 44334
rect -10719 44280 -3664 44300
rect -10719 44246 -10609 44280
rect -10575 44246 -10541 44280
rect -10507 44246 -10473 44280
rect -10439 44246 -10405 44280
rect -10371 44246 -10337 44280
rect -10303 44246 -10269 44280
rect -10235 44246 -10201 44280
rect -10167 44246 -10133 44280
rect -10099 44246 -10065 44280
rect -10031 44246 -9997 44280
rect -9963 44246 -9929 44280
rect -9895 44246 -9861 44280
rect -9827 44246 -9793 44280
rect -9759 44246 -9725 44280
rect -9691 44246 -9657 44280
rect -9623 44246 -9589 44280
rect -9555 44246 -9521 44280
rect -9487 44246 -9453 44280
rect -9419 44246 -9385 44280
rect -9351 44246 -9317 44280
rect -9283 44246 -9249 44280
rect -9215 44246 -9181 44280
rect -9147 44246 -9113 44280
rect -9079 44246 -9045 44280
rect -9011 44246 -8977 44280
rect -8943 44246 -8909 44280
rect -8875 44246 -8841 44280
rect -8807 44246 -8773 44280
rect -8739 44246 -8705 44280
rect -8671 44246 -8637 44280
rect -8603 44246 -8569 44280
rect -8535 44246 -8501 44280
rect -8467 44246 -8433 44280
rect -8399 44246 -8365 44280
rect -8331 44246 -8297 44280
rect -8263 44246 -8229 44280
rect -8195 44246 -8161 44280
rect -8127 44246 -8093 44280
rect -8059 44246 -8025 44280
rect -7991 44246 -7957 44280
rect -7923 44246 -7889 44280
rect -7855 44246 -7821 44280
rect -7787 44246 -7753 44280
rect -7719 44246 -7685 44280
rect -7651 44246 -7617 44280
rect -7583 44246 -7549 44280
rect -7515 44246 -7481 44280
rect -7447 44246 -7413 44280
rect -7379 44246 -7345 44280
rect -7311 44246 -7277 44280
rect -7243 44246 -7209 44280
rect -7175 44246 -7141 44280
rect -7107 44246 -7073 44280
rect -7039 44246 -7005 44280
rect -6971 44246 -6937 44280
rect -6903 44246 -6869 44280
rect -6835 44246 -6801 44280
rect -6767 44246 -6733 44280
rect -6699 44246 -6665 44280
rect -6631 44246 -6597 44280
rect -6563 44246 -6529 44280
rect -6495 44246 -6461 44280
rect -6427 44246 -6393 44280
rect -6359 44246 -6325 44280
rect -6291 44246 -6257 44280
rect -6223 44246 -6189 44280
rect -6155 44246 -6121 44280
rect -6087 44246 -6053 44280
rect -6019 44246 -5985 44280
rect -5951 44246 -5917 44280
rect -5883 44246 -5849 44280
rect -5815 44246 -5781 44280
rect -5747 44246 -5713 44280
rect -5679 44246 -5645 44280
rect -5611 44246 -5577 44280
rect -5543 44246 -5509 44280
rect -5475 44246 -5441 44280
rect -5407 44246 -5373 44280
rect -5339 44246 -5305 44280
rect -5271 44246 -5237 44280
rect -5203 44246 -5169 44280
rect -5135 44246 -5101 44280
rect -5067 44246 -5033 44280
rect -4999 44246 -4965 44280
rect -4931 44246 -4897 44280
rect -4863 44246 -4829 44280
rect -4795 44246 -4761 44280
rect -4727 44246 -4693 44280
rect -4659 44246 -4625 44280
rect -4591 44246 -4557 44280
rect -4523 44246 -4489 44280
rect -4455 44246 -4421 44280
rect -4387 44246 -4353 44280
rect -4319 44246 -4285 44280
rect -4251 44246 -4217 44280
rect -4183 44246 -4149 44280
rect -4115 44246 -4081 44280
rect -4047 44246 -4013 44280
rect -3979 44246 -3945 44280
rect -3911 44246 -3877 44280
rect -3843 44246 -3809 44280
rect -3775 44246 -3664 44280
rect -10719 44226 -3664 44246
rect -2416 19521 47250 19541
rect -2416 19487 -2318 19521
rect -2284 19487 -2250 19521
rect -2216 19487 -2182 19521
rect -2148 19487 -2114 19521
rect -2080 19487 -2046 19521
rect -2012 19487 -1978 19521
rect -1944 19487 -1910 19521
rect -1876 19487 -1842 19521
rect -1808 19487 -1774 19521
rect -1740 19487 -1706 19521
rect -1672 19487 -1638 19521
rect -1604 19487 -1570 19521
rect -1536 19487 -1502 19521
rect -1468 19487 -1434 19521
rect -1400 19487 -1366 19521
rect -1332 19487 -1298 19521
rect -1264 19487 -1230 19521
rect -1196 19487 -1162 19521
rect -1128 19487 -1094 19521
rect -1060 19487 -1026 19521
rect -992 19487 -958 19521
rect -924 19487 -890 19521
rect -856 19487 -822 19521
rect -788 19487 -754 19521
rect -720 19487 -686 19521
rect -652 19487 -618 19521
rect -584 19487 -550 19521
rect -516 19487 -482 19521
rect -448 19487 -414 19521
rect -380 19487 -346 19521
rect -312 19487 -278 19521
rect -244 19487 -210 19521
rect -176 19487 -142 19521
rect -108 19487 -74 19521
rect -40 19487 -6 19521
rect 28 19487 62 19521
rect 96 19487 130 19521
rect 164 19487 198 19521
rect 232 19487 266 19521
rect 300 19487 334 19521
rect 368 19487 402 19521
rect 436 19487 470 19521
rect 504 19487 538 19521
rect 572 19487 606 19521
rect 640 19487 674 19521
rect 708 19487 742 19521
rect 776 19487 810 19521
rect 844 19487 878 19521
rect 912 19487 946 19521
rect 980 19487 1014 19521
rect 1048 19487 1082 19521
rect 1116 19487 1150 19521
rect 1184 19487 1218 19521
rect 1252 19487 1286 19521
rect 1320 19487 1354 19521
rect 1388 19487 1422 19521
rect 1456 19487 1490 19521
rect 1524 19487 1558 19521
rect 1592 19487 1626 19521
rect 1660 19487 1694 19521
rect 1728 19487 1762 19521
rect 1796 19487 1830 19521
rect 1864 19487 1898 19521
rect 1932 19487 1966 19521
rect 2000 19487 2034 19521
rect 2068 19487 2102 19521
rect 2136 19487 2170 19521
rect 2204 19487 2238 19521
rect 2272 19487 2306 19521
rect 2340 19487 2374 19521
rect 2408 19487 2442 19521
rect 2476 19487 2510 19521
rect 2544 19487 2578 19521
rect 2612 19487 2646 19521
rect 2680 19487 2714 19521
rect 2748 19487 2782 19521
rect 2816 19487 2850 19521
rect 2884 19487 2918 19521
rect 2952 19487 2986 19521
rect 3020 19487 3054 19521
rect 3088 19487 3122 19521
rect 3156 19487 3190 19521
rect 3224 19487 3258 19521
rect 3292 19487 3326 19521
rect 3360 19487 3394 19521
rect 3428 19487 3462 19521
rect 3496 19487 3530 19521
rect 3564 19487 3598 19521
rect 3632 19487 3666 19521
rect 3700 19487 3734 19521
rect 3768 19487 3802 19521
rect 3836 19487 3870 19521
rect 3904 19487 3938 19521
rect 3972 19487 4006 19521
rect 4040 19487 4074 19521
rect 4108 19487 4142 19521
rect 4176 19487 4210 19521
rect 4244 19487 4278 19521
rect 4312 19487 4346 19521
rect 4380 19487 4414 19521
rect 4448 19487 4482 19521
rect 4516 19487 4550 19521
rect 4584 19487 4618 19521
rect 4652 19487 4686 19521
rect 4720 19487 4754 19521
rect 4788 19487 4822 19521
rect 4856 19487 4890 19521
rect 4924 19487 4958 19521
rect 4992 19487 5026 19521
rect 5060 19487 5094 19521
rect 5128 19487 5162 19521
rect 5196 19487 5230 19521
rect 5264 19487 5298 19521
rect 5332 19487 5366 19521
rect 5400 19487 5434 19521
rect 5468 19487 5502 19521
rect 5536 19487 5570 19521
rect 5604 19487 5638 19521
rect 5672 19487 5706 19521
rect 5740 19487 5774 19521
rect 5808 19487 5842 19521
rect 5876 19487 5910 19521
rect 5944 19487 5978 19521
rect 6012 19487 6046 19521
rect 6080 19487 6114 19521
rect 6148 19487 6182 19521
rect 6216 19487 6250 19521
rect 6284 19487 6318 19521
rect 6352 19487 6386 19521
rect 6420 19487 6454 19521
rect 6488 19487 6522 19521
rect 6556 19487 6590 19521
rect 6624 19487 6658 19521
rect 6692 19487 6726 19521
rect 6760 19487 6794 19521
rect 6828 19487 6862 19521
rect 6896 19487 6930 19521
rect 6964 19487 6998 19521
rect 7032 19487 7066 19521
rect 7100 19487 7134 19521
rect 7168 19487 7202 19521
rect 7236 19487 7270 19521
rect 7304 19487 7338 19521
rect 7372 19487 7406 19521
rect 7440 19487 7474 19521
rect 7508 19487 7542 19521
rect 7576 19487 7610 19521
rect 7644 19487 7678 19521
rect 7712 19487 7746 19521
rect 7780 19487 7814 19521
rect 7848 19487 7882 19521
rect 7916 19487 7950 19521
rect 7984 19487 8018 19521
rect 8052 19487 8086 19521
rect 8120 19487 8154 19521
rect 8188 19487 8222 19521
rect 8256 19487 8290 19521
rect 8324 19487 8358 19521
rect 8392 19487 8426 19521
rect 8460 19487 8494 19521
rect 8528 19487 8562 19521
rect 8596 19487 8630 19521
rect 8664 19487 8698 19521
rect 8732 19487 8766 19521
rect 8800 19487 8834 19521
rect 8868 19487 8902 19521
rect 8936 19487 8970 19521
rect 9004 19487 9038 19521
rect 9072 19487 9106 19521
rect 9140 19487 9174 19521
rect 9208 19487 9242 19521
rect 9276 19487 9310 19521
rect 9344 19487 9378 19521
rect 9412 19487 9446 19521
rect 9480 19487 9514 19521
rect 9548 19487 9582 19521
rect 9616 19487 9650 19521
rect 9684 19487 9718 19521
rect 9752 19487 9786 19521
rect 9820 19487 9854 19521
rect 9888 19487 9922 19521
rect 9956 19487 9990 19521
rect 10024 19487 10058 19521
rect 10092 19487 10126 19521
rect 10160 19487 10194 19521
rect 10228 19487 10262 19521
rect 10296 19487 10330 19521
rect 10364 19487 10398 19521
rect 10432 19487 10466 19521
rect 10500 19487 10534 19521
rect 10568 19487 10602 19521
rect 10636 19487 10670 19521
rect 10704 19487 10738 19521
rect 10772 19487 10806 19521
rect 10840 19487 10874 19521
rect 10908 19487 10942 19521
rect 10976 19487 11010 19521
rect 11044 19487 11078 19521
rect 11112 19487 11146 19521
rect 11180 19487 11214 19521
rect 11248 19487 11282 19521
rect 11316 19487 11350 19521
rect 11384 19487 11418 19521
rect 11452 19487 11486 19521
rect 11520 19487 11554 19521
rect 11588 19487 11622 19521
rect 11656 19487 11690 19521
rect 11724 19487 11758 19521
rect 11792 19487 11826 19521
rect 11860 19487 11894 19521
rect 11928 19487 11962 19521
rect 11996 19487 12030 19521
rect 12064 19487 12098 19521
rect 12132 19487 12166 19521
rect 12200 19487 12234 19521
rect 12268 19487 12302 19521
rect 12336 19487 12370 19521
rect 12404 19487 12438 19521
rect 12472 19487 12506 19521
rect 12540 19487 12574 19521
rect 12608 19487 12642 19521
rect 12676 19487 12710 19521
rect 12744 19487 12778 19521
rect 12812 19487 12846 19521
rect 12880 19487 12914 19521
rect 12948 19487 12982 19521
rect 13016 19487 13050 19521
rect 13084 19487 13118 19521
rect 13152 19487 13186 19521
rect 13220 19487 13254 19521
rect 13288 19487 13322 19521
rect 13356 19487 13390 19521
rect 13424 19487 13458 19521
rect 13492 19487 13526 19521
rect 13560 19487 13594 19521
rect 13628 19487 13662 19521
rect 13696 19487 13730 19521
rect 13764 19487 13798 19521
rect 13832 19487 13866 19521
rect 13900 19487 13934 19521
rect 13968 19487 14002 19521
rect 14036 19487 14070 19521
rect 14104 19487 14138 19521
rect 14172 19487 14206 19521
rect 14240 19487 14274 19521
rect 14308 19487 14342 19521
rect 14376 19487 14410 19521
rect 14444 19487 14478 19521
rect 14512 19487 14546 19521
rect 14580 19487 14614 19521
rect 14648 19487 14682 19521
rect 14716 19487 14750 19521
rect 14784 19487 14818 19521
rect 14852 19487 14886 19521
rect 14920 19487 14954 19521
rect 14988 19487 15022 19521
rect 15056 19487 15090 19521
rect 15124 19487 15158 19521
rect 15192 19487 15226 19521
rect 15260 19487 15294 19521
rect 15328 19487 15362 19521
rect 15396 19487 15430 19521
rect 15464 19487 15498 19521
rect 15532 19487 15566 19521
rect 15600 19487 15634 19521
rect 15668 19487 15702 19521
rect 15736 19487 15770 19521
rect 15804 19487 15838 19521
rect 15872 19487 15906 19521
rect 15940 19487 15974 19521
rect 16008 19487 16042 19521
rect 16076 19487 16110 19521
rect 16144 19487 16178 19521
rect 16212 19487 16246 19521
rect 16280 19487 16314 19521
rect 16348 19487 16382 19521
rect 16416 19487 16450 19521
rect 16484 19487 16518 19521
rect 16552 19487 16586 19521
rect 16620 19487 16654 19521
rect 16688 19487 16722 19521
rect 16756 19487 16790 19521
rect 16824 19487 16858 19521
rect 16892 19487 16926 19521
rect 16960 19487 16994 19521
rect 17028 19487 17062 19521
rect 17096 19487 17130 19521
rect 17164 19487 17198 19521
rect 17232 19487 17266 19521
rect 17300 19487 17334 19521
rect 17368 19487 17402 19521
rect 17436 19487 17470 19521
rect 17504 19487 17538 19521
rect 17572 19487 17606 19521
rect 17640 19487 17674 19521
rect 17708 19487 17742 19521
rect 17776 19487 17810 19521
rect 17844 19487 17878 19521
rect 17912 19487 17946 19521
rect 17980 19487 18014 19521
rect 18048 19487 18082 19521
rect 18116 19487 18150 19521
rect 18184 19487 18218 19521
rect 18252 19487 18286 19521
rect 18320 19487 18354 19521
rect 18388 19487 18422 19521
rect 18456 19487 18490 19521
rect 18524 19487 18558 19521
rect 18592 19487 18626 19521
rect 18660 19487 18694 19521
rect 18728 19487 18762 19521
rect 18796 19487 18830 19521
rect 18864 19487 18898 19521
rect 18932 19487 18966 19521
rect 19000 19487 19034 19521
rect 19068 19487 19102 19521
rect 19136 19487 19170 19521
rect 19204 19487 19238 19521
rect 19272 19487 19306 19521
rect 19340 19487 19374 19521
rect 19408 19487 19442 19521
rect 19476 19487 19510 19521
rect 19544 19487 19578 19521
rect 19612 19487 19646 19521
rect 19680 19487 19714 19521
rect 19748 19487 19782 19521
rect 19816 19487 19850 19521
rect 19884 19487 19918 19521
rect 19952 19487 19986 19521
rect 20020 19487 20054 19521
rect 20088 19487 20122 19521
rect 20156 19487 20190 19521
rect 20224 19487 20258 19521
rect 20292 19487 20326 19521
rect 20360 19487 20394 19521
rect 20428 19487 20462 19521
rect 20496 19487 20530 19521
rect 20564 19487 20598 19521
rect 20632 19487 20666 19521
rect 20700 19487 20734 19521
rect 20768 19487 20802 19521
rect 20836 19487 20870 19521
rect 20904 19487 20938 19521
rect 20972 19487 21006 19521
rect 21040 19487 21074 19521
rect 21108 19487 21142 19521
rect 21176 19487 21210 19521
rect 21244 19487 21278 19521
rect 21312 19487 21346 19521
rect 21380 19487 21414 19521
rect 21448 19487 21482 19521
rect 21516 19487 21550 19521
rect 21584 19487 21618 19521
rect 21652 19487 21686 19521
rect 21720 19487 21754 19521
rect 21788 19487 21822 19521
rect 21856 19487 21890 19521
rect 21924 19487 21958 19521
rect 21992 19487 22026 19521
rect 22060 19487 22094 19521
rect 22128 19487 22162 19521
rect 22196 19487 22230 19521
rect 22264 19487 22298 19521
rect 22332 19487 22366 19521
rect 22400 19487 22434 19521
rect 22468 19487 22502 19521
rect 22536 19487 22570 19521
rect 22604 19487 22638 19521
rect 22672 19487 22706 19521
rect 22740 19487 22774 19521
rect 22808 19487 22842 19521
rect 22876 19487 22910 19521
rect 22944 19487 22978 19521
rect 23012 19487 23046 19521
rect 23080 19487 23114 19521
rect 23148 19487 23182 19521
rect 23216 19487 23250 19521
rect 23284 19487 23318 19521
rect 23352 19487 23386 19521
rect 23420 19487 23454 19521
rect 23488 19487 23522 19521
rect 23556 19487 23590 19521
rect 23624 19487 23658 19521
rect 23692 19487 23726 19521
rect 23760 19487 23794 19521
rect 23828 19487 23862 19521
rect 23896 19487 23930 19521
rect 23964 19487 23998 19521
rect 24032 19487 24066 19521
rect 24100 19487 24134 19521
rect 24168 19487 24202 19521
rect 24236 19487 24270 19521
rect 24304 19487 24338 19521
rect 24372 19487 24406 19521
rect 24440 19487 24474 19521
rect 24508 19487 24542 19521
rect 24576 19487 24610 19521
rect 24644 19487 24678 19521
rect 24712 19487 24746 19521
rect 24780 19487 24814 19521
rect 24848 19487 24882 19521
rect 24916 19487 24950 19521
rect 24984 19487 25018 19521
rect 25052 19487 25086 19521
rect 25120 19487 25154 19521
rect 25188 19487 25222 19521
rect 25256 19487 25290 19521
rect 25324 19487 25358 19521
rect 25392 19487 25426 19521
rect 25460 19487 25494 19521
rect 25528 19487 25562 19521
rect 25596 19487 25630 19521
rect 25664 19487 25698 19521
rect 25732 19487 25766 19521
rect 25800 19487 25834 19521
rect 25868 19487 25902 19521
rect 25936 19487 25970 19521
rect 26004 19487 26038 19521
rect 26072 19487 26106 19521
rect 26140 19487 26174 19521
rect 26208 19487 26242 19521
rect 26276 19487 26310 19521
rect 26344 19487 26378 19521
rect 26412 19487 26446 19521
rect 26480 19487 26514 19521
rect 26548 19487 26582 19521
rect 26616 19487 26650 19521
rect 26684 19487 26718 19521
rect 26752 19487 26786 19521
rect 26820 19487 26854 19521
rect 26888 19487 26922 19521
rect 26956 19487 26990 19521
rect 27024 19487 27058 19521
rect 27092 19487 27126 19521
rect 27160 19487 27194 19521
rect 27228 19487 27262 19521
rect 27296 19487 27330 19521
rect 27364 19487 27398 19521
rect 27432 19487 27466 19521
rect 27500 19487 27534 19521
rect 27568 19487 27602 19521
rect 27636 19487 27670 19521
rect 27704 19487 27738 19521
rect 27772 19487 27806 19521
rect 27840 19487 27874 19521
rect 27908 19487 27942 19521
rect 27976 19487 28010 19521
rect 28044 19487 28078 19521
rect 28112 19487 28146 19521
rect 28180 19487 28214 19521
rect 28248 19487 28282 19521
rect 28316 19487 28350 19521
rect 28384 19487 28418 19521
rect 28452 19487 28486 19521
rect 28520 19487 28554 19521
rect 28588 19487 28622 19521
rect 28656 19487 28690 19521
rect 28724 19487 28758 19521
rect 28792 19487 28826 19521
rect 28860 19487 28894 19521
rect 28928 19487 28962 19521
rect 28996 19487 29030 19521
rect 29064 19487 29098 19521
rect 29132 19487 29166 19521
rect 29200 19487 29234 19521
rect 29268 19487 29302 19521
rect 29336 19487 29370 19521
rect 29404 19487 29438 19521
rect 29472 19487 29506 19521
rect 29540 19487 29574 19521
rect 29608 19487 29642 19521
rect 29676 19487 29710 19521
rect 29744 19487 29778 19521
rect 29812 19487 29846 19521
rect 29880 19487 29914 19521
rect 29948 19487 29982 19521
rect 30016 19487 30050 19521
rect 30084 19487 30118 19521
rect 30152 19487 30186 19521
rect 30220 19487 30254 19521
rect 30288 19487 30322 19521
rect 30356 19487 30390 19521
rect 30424 19487 30458 19521
rect 30492 19487 30526 19521
rect 30560 19487 30594 19521
rect 30628 19487 30662 19521
rect 30696 19487 30730 19521
rect 30764 19487 30798 19521
rect 30832 19487 30866 19521
rect 30900 19487 30934 19521
rect 30968 19487 31002 19521
rect 31036 19487 31070 19521
rect 31104 19487 31138 19521
rect 31172 19487 31206 19521
rect 31240 19487 31274 19521
rect 31308 19487 31342 19521
rect 31376 19487 31410 19521
rect 31444 19487 31478 19521
rect 31512 19487 31546 19521
rect 31580 19487 31614 19521
rect 31648 19487 31682 19521
rect 31716 19487 31750 19521
rect 31784 19487 31818 19521
rect 31852 19487 31886 19521
rect 31920 19487 31954 19521
rect 31988 19487 32022 19521
rect 32056 19487 32090 19521
rect 32124 19487 32158 19521
rect 32192 19487 32226 19521
rect 32260 19487 32294 19521
rect 32328 19487 32362 19521
rect 32396 19487 32430 19521
rect 32464 19487 32498 19521
rect 32532 19487 32566 19521
rect 32600 19487 32634 19521
rect 32668 19487 32702 19521
rect 32736 19487 32770 19521
rect 32804 19487 32838 19521
rect 32872 19487 32906 19521
rect 32940 19487 32974 19521
rect 33008 19487 33042 19521
rect 33076 19487 33110 19521
rect 33144 19487 33178 19521
rect 33212 19487 33246 19521
rect 33280 19487 33314 19521
rect 33348 19487 33382 19521
rect 33416 19487 33450 19521
rect 33484 19487 33518 19521
rect 33552 19487 33586 19521
rect 33620 19487 33654 19521
rect 33688 19487 33722 19521
rect 33756 19487 33790 19521
rect 33824 19487 33858 19521
rect 33892 19487 33926 19521
rect 33960 19487 33994 19521
rect 34028 19487 34062 19521
rect 34096 19487 34130 19521
rect 34164 19487 34198 19521
rect 34232 19487 34266 19521
rect 34300 19487 34334 19521
rect 34368 19487 34402 19521
rect 34436 19487 34470 19521
rect 34504 19487 34538 19521
rect 34572 19487 34606 19521
rect 34640 19487 34674 19521
rect 34708 19487 34742 19521
rect 34776 19487 34810 19521
rect 34844 19487 34878 19521
rect 34912 19487 34946 19521
rect 34980 19487 35014 19521
rect 35048 19487 35082 19521
rect 35116 19487 35150 19521
rect 35184 19487 35218 19521
rect 35252 19487 35286 19521
rect 35320 19487 35354 19521
rect 35388 19487 35422 19521
rect 35456 19487 35490 19521
rect 35524 19487 35558 19521
rect 35592 19487 35626 19521
rect 35660 19487 35694 19521
rect 35728 19487 35762 19521
rect 35796 19487 35830 19521
rect 35864 19487 35898 19521
rect 35932 19487 35966 19521
rect 36000 19487 36034 19521
rect 36068 19487 36102 19521
rect 36136 19487 36170 19521
rect 36204 19487 36238 19521
rect 36272 19487 36306 19521
rect 36340 19487 36374 19521
rect 36408 19487 36442 19521
rect 36476 19487 36510 19521
rect 36544 19487 36578 19521
rect 36612 19487 36646 19521
rect 36680 19487 36714 19521
rect 36748 19487 36782 19521
rect 36816 19487 36850 19521
rect 36884 19487 36918 19521
rect 36952 19487 36986 19521
rect 37020 19487 37054 19521
rect 37088 19487 37122 19521
rect 37156 19487 37190 19521
rect 37224 19487 37258 19521
rect 37292 19487 37326 19521
rect 37360 19487 37394 19521
rect 37428 19487 37462 19521
rect 37496 19487 37530 19521
rect 37564 19487 37598 19521
rect 37632 19487 37666 19521
rect 37700 19487 37734 19521
rect 37768 19487 37802 19521
rect 37836 19487 37870 19521
rect 37904 19487 37938 19521
rect 37972 19487 38006 19521
rect 38040 19487 38074 19521
rect 38108 19487 38142 19521
rect 38176 19487 38210 19521
rect 38244 19487 38278 19521
rect 38312 19487 38346 19521
rect 38380 19487 38414 19521
rect 38448 19487 38482 19521
rect 38516 19487 38550 19521
rect 38584 19487 38618 19521
rect 38652 19487 38686 19521
rect 38720 19487 38754 19521
rect 38788 19487 38822 19521
rect 38856 19487 38890 19521
rect 38924 19487 38958 19521
rect 38992 19487 39026 19521
rect 39060 19487 39094 19521
rect 39128 19487 39162 19521
rect 39196 19487 39230 19521
rect 39264 19487 39298 19521
rect 39332 19487 39366 19521
rect 39400 19487 39434 19521
rect 39468 19487 39502 19521
rect 39536 19487 39570 19521
rect 39604 19487 39638 19521
rect 39672 19487 39706 19521
rect 39740 19487 39774 19521
rect 39808 19487 39842 19521
rect 39876 19487 39910 19521
rect 39944 19487 39978 19521
rect 40012 19487 40046 19521
rect 40080 19487 40114 19521
rect 40148 19487 40182 19521
rect 40216 19487 40250 19521
rect 40284 19487 40318 19521
rect 40352 19487 40386 19521
rect 40420 19487 40454 19521
rect 40488 19487 40522 19521
rect 40556 19487 40590 19521
rect 40624 19487 40658 19521
rect 40692 19487 40726 19521
rect 40760 19487 40794 19521
rect 40828 19487 40862 19521
rect 40896 19487 40930 19521
rect 40964 19487 40998 19521
rect 41032 19487 41066 19521
rect 41100 19487 41134 19521
rect 41168 19487 41202 19521
rect 41236 19487 41270 19521
rect 41304 19487 41338 19521
rect 41372 19487 41406 19521
rect 41440 19487 41474 19521
rect 41508 19487 41542 19521
rect 41576 19487 41610 19521
rect 41644 19487 41678 19521
rect 41712 19487 41746 19521
rect 41780 19487 41814 19521
rect 41848 19487 41882 19521
rect 41916 19487 41950 19521
rect 41984 19487 42018 19521
rect 42052 19487 42086 19521
rect 42120 19487 42154 19521
rect 42188 19487 42222 19521
rect 42256 19487 42290 19521
rect 42324 19487 42358 19521
rect 42392 19487 42426 19521
rect 42460 19487 42494 19521
rect 42528 19487 42562 19521
rect 42596 19487 42630 19521
rect 42664 19487 42698 19521
rect 42732 19487 42766 19521
rect 42800 19487 42834 19521
rect 42868 19487 42902 19521
rect 42936 19487 42970 19521
rect 43004 19487 43038 19521
rect 43072 19487 43106 19521
rect 43140 19487 43174 19521
rect 43208 19487 43242 19521
rect 43276 19487 43310 19521
rect 43344 19487 43378 19521
rect 43412 19487 43446 19521
rect 43480 19487 43514 19521
rect 43548 19487 43582 19521
rect 43616 19487 43650 19521
rect 43684 19487 43718 19521
rect 43752 19487 43786 19521
rect 43820 19487 43854 19521
rect 43888 19487 43922 19521
rect 43956 19487 43990 19521
rect 44024 19487 44058 19521
rect 44092 19487 44126 19521
rect 44160 19487 44194 19521
rect 44228 19487 44262 19521
rect 44296 19487 44330 19521
rect 44364 19487 44398 19521
rect 44432 19487 44466 19521
rect 44500 19487 44534 19521
rect 44568 19487 44602 19521
rect 44636 19487 44670 19521
rect 44704 19487 44738 19521
rect 44772 19487 44806 19521
rect 44840 19487 44874 19521
rect 44908 19487 44942 19521
rect 44976 19487 45010 19521
rect 45044 19487 45078 19521
rect 45112 19487 45146 19521
rect 45180 19487 45214 19521
rect 45248 19487 45282 19521
rect 45316 19487 45350 19521
rect 45384 19487 45418 19521
rect 45452 19487 45486 19521
rect 45520 19487 45554 19521
rect 45588 19487 45622 19521
rect 45656 19487 45690 19521
rect 45724 19487 45758 19521
rect 45792 19487 45826 19521
rect 45860 19487 45894 19521
rect 45928 19487 45962 19521
rect 45996 19487 46030 19521
rect 46064 19487 46098 19521
rect 46132 19487 46166 19521
rect 46200 19487 46234 19521
rect 46268 19487 46302 19521
rect 46336 19487 46370 19521
rect 46404 19487 46438 19521
rect 46472 19487 46506 19521
rect 46540 19487 46574 19521
rect 46608 19487 46642 19521
rect 46676 19487 46710 19521
rect 46744 19487 46778 19521
rect 46812 19487 46846 19521
rect 46880 19487 46914 19521
rect 46948 19487 46982 19521
rect 47016 19487 47050 19521
rect 47084 19487 47118 19521
rect 47152 19487 47250 19521
rect -2416 19467 47250 19487
rect -2416 19434 -2342 19467
rect -2416 19400 -2396 19434
rect -2362 19400 -2342 19434
rect -2416 19366 -2342 19400
rect -2416 19332 -2396 19366
rect -2362 19332 -2342 19366
rect -2416 19298 -2342 19332
rect -2416 19264 -2396 19298
rect -2362 19264 -2342 19298
rect -2416 19230 -2342 19264
rect -2416 19196 -2396 19230
rect -2362 19196 -2342 19230
rect -2416 19162 -2342 19196
rect -2416 19128 -2396 19162
rect -2362 19128 -2342 19162
rect -2416 19094 -2342 19128
rect -2416 19060 -2396 19094
rect -2362 19060 -2342 19094
rect -2416 19026 -2342 19060
rect -2416 18992 -2396 19026
rect -2362 18992 -2342 19026
rect -2416 18958 -2342 18992
rect -2416 18924 -2396 18958
rect -2362 18924 -2342 18958
rect -2416 18890 -2342 18924
rect -2416 18856 -2396 18890
rect -2362 18856 -2342 18890
rect -2416 18822 -2342 18856
rect -2416 18788 -2396 18822
rect -2362 18788 -2342 18822
rect -2416 18754 -2342 18788
rect -2416 18720 -2396 18754
rect -2362 18720 -2342 18754
rect -2416 18686 -2342 18720
rect -2416 18652 -2396 18686
rect -2362 18652 -2342 18686
rect -2416 18618 -2342 18652
rect -2416 18584 -2396 18618
rect -2362 18584 -2342 18618
rect -2416 18550 -2342 18584
rect -2416 18516 -2396 18550
rect -2362 18516 -2342 18550
rect -2416 18482 -2342 18516
rect -2416 18448 -2396 18482
rect -2362 18448 -2342 18482
rect -2416 18414 -2342 18448
rect -2416 18380 -2396 18414
rect -2362 18380 -2342 18414
rect -2416 18346 -2342 18380
rect -2416 18312 -2396 18346
rect -2362 18312 -2342 18346
rect -2416 18278 -2342 18312
rect -2416 18244 -2396 18278
rect -2362 18244 -2342 18278
rect -2416 18210 -2342 18244
rect -2416 18176 -2396 18210
rect -2362 18176 -2342 18210
rect -2416 18142 -2342 18176
rect -2416 18108 -2396 18142
rect -2362 18108 -2342 18142
rect -2416 18074 -2342 18108
rect -2416 18040 -2396 18074
rect -2362 18040 -2342 18074
rect -2416 18006 -2342 18040
rect -2416 17972 -2396 18006
rect -2362 17972 -2342 18006
rect -2416 17938 -2342 17972
rect -2416 17904 -2396 17938
rect -2362 17904 -2342 17938
rect -2416 17870 -2342 17904
rect -2416 17836 -2396 17870
rect -2362 17836 -2342 17870
rect -2416 17802 -2342 17836
rect -2416 17768 -2396 17802
rect -2362 17768 -2342 17802
rect -2416 17734 -2342 17768
rect -2416 17700 -2396 17734
rect -2362 17700 -2342 17734
rect -2416 17666 -2342 17700
rect -2416 17632 -2396 17666
rect -2362 17632 -2342 17666
rect -2416 17598 -2342 17632
rect -2416 17564 -2396 17598
rect -2362 17564 -2342 17598
rect -2416 17530 -2342 17564
rect -2416 17496 -2396 17530
rect -2362 17496 -2342 17530
rect -2416 17462 -2342 17496
rect -2416 17428 -2396 17462
rect -2362 17428 -2342 17462
rect -2416 17394 -2342 17428
rect -2416 17360 -2396 17394
rect -2362 17360 -2342 17394
rect -2416 17326 -2342 17360
rect -2416 17292 -2396 17326
rect -2362 17292 -2342 17326
rect -2416 17258 -2342 17292
rect -2416 17224 -2396 17258
rect -2362 17224 -2342 17258
rect -2416 17190 -2342 17224
rect -2416 17156 -2396 17190
rect -2362 17156 -2342 17190
rect -2416 17122 -2342 17156
rect -2416 17088 -2396 17122
rect -2362 17088 -2342 17122
rect -2416 17054 -2342 17088
rect -2416 17020 -2396 17054
rect -2362 17020 -2342 17054
rect -2416 16986 -2342 17020
rect -2416 16952 -2396 16986
rect -2362 16952 -2342 16986
rect -2416 16918 -2342 16952
rect -2416 16884 -2396 16918
rect -2362 16884 -2342 16918
rect -2416 16850 -2342 16884
rect -2416 16816 -2396 16850
rect -2362 16816 -2342 16850
rect -2416 16782 -2342 16816
rect -2416 16748 -2396 16782
rect -2362 16748 -2342 16782
rect -2416 16714 -2342 16748
rect -2416 16680 -2396 16714
rect -2362 16680 -2342 16714
rect -2416 16646 -2342 16680
rect -2416 16612 -2396 16646
rect -2362 16612 -2342 16646
rect -2416 16578 -2342 16612
rect -2416 16544 -2396 16578
rect -2362 16544 -2342 16578
rect -2416 16510 -2342 16544
rect -2416 16476 -2396 16510
rect -2362 16476 -2342 16510
rect -2416 16442 -2342 16476
rect -2416 16408 -2396 16442
rect -2362 16408 -2342 16442
rect -2416 16374 -2342 16408
rect -2416 16340 -2396 16374
rect -2362 16340 -2342 16374
rect -2416 16306 -2342 16340
rect -2416 16272 -2396 16306
rect -2362 16272 -2342 16306
rect -2416 16238 -2342 16272
rect -2416 16204 -2396 16238
rect -2362 16204 -2342 16238
rect -2416 16170 -2342 16204
rect -2416 16136 -2396 16170
rect -2362 16136 -2342 16170
rect -2416 16102 -2342 16136
rect -2416 16068 -2396 16102
rect -2362 16068 -2342 16102
rect -2416 16034 -2342 16068
rect -2416 16000 -2396 16034
rect -2362 16000 -2342 16034
rect -2416 15966 -2342 16000
rect -2416 15932 -2396 15966
rect -2362 15932 -2342 15966
rect -2416 15898 -2342 15932
rect -2416 15864 -2396 15898
rect -2362 15864 -2342 15898
rect -2416 15830 -2342 15864
rect -2416 15796 -2396 15830
rect -2362 15796 -2342 15830
rect -2416 15762 -2342 15796
rect -2416 15728 -2396 15762
rect -2362 15728 -2342 15762
rect -2416 15694 -2342 15728
rect -2416 15660 -2396 15694
rect -2362 15660 -2342 15694
rect -2416 15626 -2342 15660
rect -2416 15592 -2396 15626
rect -2362 15592 -2342 15626
rect -2416 15558 -2342 15592
rect -2416 15524 -2396 15558
rect -2362 15524 -2342 15558
rect -2416 15490 -2342 15524
rect -2416 15456 -2396 15490
rect -2362 15456 -2342 15490
rect -2416 15422 -2342 15456
rect -2416 15388 -2396 15422
rect -2362 15388 -2342 15422
rect -2416 15354 -2342 15388
rect -2416 15320 -2396 15354
rect -2362 15320 -2342 15354
rect -2416 15286 -2342 15320
rect -2416 15252 -2396 15286
rect -2362 15252 -2342 15286
rect -2416 15218 -2342 15252
rect -2416 15184 -2396 15218
rect -2362 15184 -2342 15218
rect -2416 15150 -2342 15184
rect -2416 15116 -2396 15150
rect -2362 15116 -2342 15150
rect -2416 15082 -2342 15116
rect -2416 15048 -2396 15082
rect -2362 15048 -2342 15082
rect -2416 15014 -2342 15048
rect -2416 14980 -2396 15014
rect -2362 14980 -2342 15014
rect -2416 14946 -2342 14980
rect -2416 14912 -2396 14946
rect -2362 14912 -2342 14946
rect -2416 14878 -2342 14912
rect -2416 14844 -2396 14878
rect -2362 14844 -2342 14878
rect -2416 14810 -2342 14844
rect -2416 14776 -2396 14810
rect -2362 14776 -2342 14810
rect -2416 14742 -2342 14776
rect -2416 14708 -2396 14742
rect -2362 14708 -2342 14742
rect -2416 14674 -2342 14708
rect -2416 14640 -2396 14674
rect -2362 14640 -2342 14674
rect -2416 14606 -2342 14640
rect -2416 14572 -2396 14606
rect -2362 14572 -2342 14606
rect -2416 14538 -2342 14572
rect -2416 14504 -2396 14538
rect -2362 14504 -2342 14538
rect -2416 14470 -2342 14504
rect -2416 14436 -2396 14470
rect -2362 14436 -2342 14470
rect -2416 14402 -2342 14436
rect -2416 14368 -2396 14402
rect -2362 14368 -2342 14402
rect -2416 14334 -2342 14368
rect -2416 14300 -2396 14334
rect -2362 14300 -2342 14334
rect -2416 14266 -2342 14300
rect -2416 14232 -2396 14266
rect -2362 14232 -2342 14266
rect -2416 14198 -2342 14232
rect -2416 14164 -2396 14198
rect -2362 14164 -2342 14198
rect -2416 14130 -2342 14164
rect -2416 14096 -2396 14130
rect -2362 14096 -2342 14130
rect -2416 14062 -2342 14096
rect -2416 14028 -2396 14062
rect -2362 14028 -2342 14062
rect -2416 13994 -2342 14028
rect -2416 13960 -2396 13994
rect -2362 13960 -2342 13994
rect -2416 13926 -2342 13960
rect -2416 13892 -2396 13926
rect -2362 13892 -2342 13926
rect -2416 13858 -2342 13892
rect -2416 13824 -2396 13858
rect -2362 13824 -2342 13858
rect -2416 13790 -2342 13824
rect -2416 13756 -2396 13790
rect -2362 13756 -2342 13790
rect -2416 13722 -2342 13756
rect -2416 13688 -2396 13722
rect -2362 13688 -2342 13722
rect -2416 13654 -2342 13688
rect -2416 13620 -2396 13654
rect -2362 13620 -2342 13654
rect -2416 13586 -2342 13620
rect -2416 13552 -2396 13586
rect -2362 13552 -2342 13586
rect -2416 13518 -2342 13552
rect -2416 13484 -2396 13518
rect -2362 13484 -2342 13518
rect -2416 13450 -2342 13484
rect -2416 13416 -2396 13450
rect -2362 13416 -2342 13450
rect -2416 13382 -2342 13416
rect -2416 13348 -2396 13382
rect -2362 13348 -2342 13382
rect -2416 13314 -2342 13348
rect -2416 13280 -2396 13314
rect -2362 13280 -2342 13314
rect -2416 13246 -2342 13280
rect -2416 13212 -2396 13246
rect -2362 13212 -2342 13246
rect -2416 13178 -2342 13212
rect -2416 13144 -2396 13178
rect -2362 13144 -2342 13178
rect -2416 13110 -2342 13144
rect -2416 13076 -2396 13110
rect -2362 13076 -2342 13110
rect -2416 13042 -2342 13076
rect -2416 13008 -2396 13042
rect -2362 13008 -2342 13042
rect -2416 12974 -2342 13008
rect -2416 12940 -2396 12974
rect -2362 12940 -2342 12974
rect -2416 12906 -2342 12940
rect -2416 12872 -2396 12906
rect -2362 12872 -2342 12906
rect -2416 12838 -2342 12872
rect -2416 12804 -2396 12838
rect -2362 12804 -2342 12838
rect -2416 12770 -2342 12804
rect -2416 12736 -2396 12770
rect -2362 12736 -2342 12770
rect -2416 12702 -2342 12736
rect -2416 12668 -2396 12702
rect -2362 12668 -2342 12702
rect -2416 12634 -2342 12668
rect -2416 12600 -2396 12634
rect -2362 12600 -2342 12634
rect -2416 12566 -2342 12600
rect -2416 12532 -2396 12566
rect -2362 12532 -2342 12566
rect -2416 12498 -2342 12532
rect -2416 12464 -2396 12498
rect -2362 12464 -2342 12498
rect -2416 12430 -2342 12464
rect -2416 12396 -2396 12430
rect -2362 12396 -2342 12430
rect -2416 12362 -2342 12396
rect -2416 12328 -2396 12362
rect -2362 12328 -2342 12362
rect -2416 12294 -2342 12328
rect -2416 12260 -2396 12294
rect -2362 12260 -2342 12294
rect -2416 12226 -2342 12260
rect -2416 12192 -2396 12226
rect -2362 12192 -2342 12226
rect -2416 12158 -2342 12192
rect -2416 12124 -2396 12158
rect -2362 12124 -2342 12158
rect -2416 12090 -2342 12124
rect -2416 12056 -2396 12090
rect -2362 12056 -2342 12090
rect -2416 12022 -2342 12056
rect -2416 11988 -2396 12022
rect -2362 11988 -2342 12022
rect -2416 11954 -2342 11988
rect -2416 11920 -2396 11954
rect -2362 11920 -2342 11954
rect -2416 11886 -2342 11920
rect -2416 11852 -2396 11886
rect -2362 11852 -2342 11886
rect -2416 11818 -2342 11852
rect -2416 11784 -2396 11818
rect -2362 11784 -2342 11818
rect -2416 11750 -2342 11784
rect -2416 11716 -2396 11750
rect -2362 11716 -2342 11750
rect -2416 11682 -2342 11716
rect -2416 11648 -2396 11682
rect -2362 11648 -2342 11682
rect -2416 11614 -2342 11648
rect -2416 11580 -2396 11614
rect -2362 11580 -2342 11614
rect -2416 11546 -2342 11580
rect -2416 11512 -2396 11546
rect -2362 11512 -2342 11546
rect -2416 11478 -2342 11512
rect -2416 11444 -2396 11478
rect -2362 11444 -2342 11478
rect -2416 11410 -2342 11444
rect -2416 11376 -2396 11410
rect -2362 11376 -2342 11410
rect -2416 11342 -2342 11376
rect -2416 11308 -2396 11342
rect -2362 11308 -2342 11342
rect -2416 11274 -2342 11308
rect -2416 11240 -2396 11274
rect -2362 11240 -2342 11274
rect -2416 11206 -2342 11240
rect -2416 11172 -2396 11206
rect -2362 11172 -2342 11206
rect -2416 11138 -2342 11172
rect -2416 11104 -2396 11138
rect -2362 11104 -2342 11138
rect -2416 11070 -2342 11104
rect -2416 11036 -2396 11070
rect -2362 11036 -2342 11070
rect -2416 11002 -2342 11036
rect -2416 10968 -2396 11002
rect -2362 10968 -2342 11002
rect -2416 10934 -2342 10968
rect -2416 10900 -2396 10934
rect -2362 10900 -2342 10934
rect -2416 10866 -2342 10900
rect -2416 10832 -2396 10866
rect -2362 10832 -2342 10866
rect -2416 10798 -2342 10832
rect -2416 10764 -2396 10798
rect -2362 10764 -2342 10798
rect -2416 10730 -2342 10764
rect -2416 10696 -2396 10730
rect -2362 10696 -2342 10730
rect -2416 10662 -2342 10696
rect -2416 10628 -2396 10662
rect -2362 10628 -2342 10662
rect -2416 10594 -2342 10628
rect -2416 10560 -2396 10594
rect -2362 10560 -2342 10594
rect -2416 10526 -2342 10560
rect -2416 10492 -2396 10526
rect -2362 10492 -2342 10526
rect -2416 10458 -2342 10492
rect -2416 10424 -2396 10458
rect -2362 10424 -2342 10458
rect -2416 10390 -2342 10424
rect -2416 10356 -2396 10390
rect -2362 10356 -2342 10390
rect -2416 10322 -2342 10356
rect -2416 10288 -2396 10322
rect -2362 10288 -2342 10322
rect -2416 10254 -2342 10288
rect -2416 10220 -2396 10254
rect -2362 10220 -2342 10254
rect -2416 10186 -2342 10220
rect -2416 10152 -2396 10186
rect -2362 10152 -2342 10186
rect -2416 10118 -2342 10152
rect -2416 10084 -2396 10118
rect -2362 10084 -2342 10118
rect -2416 10050 -2342 10084
rect -2416 10016 -2396 10050
rect -2362 10016 -2342 10050
rect -2416 9982 -2342 10016
rect -2416 9948 -2396 9982
rect -2362 9948 -2342 9982
rect -2416 9914 -2342 9948
rect -2416 9880 -2396 9914
rect -2362 9880 -2342 9914
rect -2416 9846 -2342 9880
rect -2416 9812 -2396 9846
rect -2362 9812 -2342 9846
rect -2416 9778 -2342 9812
rect -2416 9744 -2396 9778
rect -2362 9744 -2342 9778
rect -2416 9710 -2342 9744
rect -2416 9676 -2396 9710
rect -2362 9676 -2342 9710
rect -2416 9642 -2342 9676
rect -2416 9608 -2396 9642
rect -2362 9608 -2342 9642
rect -2416 9574 -2342 9608
rect -2416 9540 -2396 9574
rect -2362 9540 -2342 9574
rect -2416 9506 -2342 9540
rect -2416 9472 -2396 9506
rect -2362 9472 -2342 9506
rect -2416 9438 -2342 9472
rect -2416 9404 -2396 9438
rect -2362 9404 -2342 9438
rect -2416 9370 -2342 9404
rect -2416 9336 -2396 9370
rect -2362 9336 -2342 9370
rect -2416 9302 -2342 9336
rect -2416 9268 -2396 9302
rect -2362 9268 -2342 9302
rect -2416 9234 -2342 9268
rect -2416 9200 -2396 9234
rect -2362 9200 -2342 9234
rect -2416 9166 -2342 9200
rect -2416 9132 -2396 9166
rect -2362 9132 -2342 9166
rect -2416 9098 -2342 9132
rect -2416 9064 -2396 9098
rect -2362 9064 -2342 9098
rect -2416 9030 -2342 9064
rect -2416 8996 -2396 9030
rect -2362 8996 -2342 9030
rect -2416 8962 -2342 8996
rect -2416 8928 -2396 8962
rect -2362 8928 -2342 8962
rect -2416 8894 -2342 8928
rect -2416 8860 -2396 8894
rect -2362 8860 -2342 8894
rect -2416 8826 -2342 8860
rect -2416 8792 -2396 8826
rect -2362 8792 -2342 8826
rect -2416 8758 -2342 8792
rect -2416 8724 -2396 8758
rect -2362 8724 -2342 8758
rect -2416 8690 -2342 8724
rect -2416 8656 -2396 8690
rect -2362 8656 -2342 8690
rect -2416 8622 -2342 8656
rect -2416 8588 -2396 8622
rect -2362 8588 -2342 8622
rect -2416 8554 -2342 8588
rect -2416 8520 -2396 8554
rect -2362 8520 -2342 8554
rect -2416 8486 -2342 8520
rect -2416 8452 -2396 8486
rect -2362 8452 -2342 8486
rect -2416 8418 -2342 8452
rect -2416 8384 -2396 8418
rect -2362 8384 -2342 8418
rect -2416 8350 -2342 8384
rect -2416 8316 -2396 8350
rect -2362 8316 -2342 8350
rect -2416 8282 -2342 8316
rect -2416 8248 -2396 8282
rect -2362 8248 -2342 8282
rect -2416 8214 -2342 8248
rect -2416 8180 -2396 8214
rect -2362 8180 -2342 8214
rect -2416 8146 -2342 8180
rect -2416 8112 -2396 8146
rect -2362 8112 -2342 8146
rect -2416 8078 -2342 8112
rect -2416 8044 -2396 8078
rect -2362 8044 -2342 8078
rect -2416 8010 -2342 8044
rect -2416 7976 -2396 8010
rect -2362 7976 -2342 8010
rect -2416 7942 -2342 7976
rect -2416 7908 -2396 7942
rect -2362 7908 -2342 7942
rect -2416 7874 -2342 7908
rect -2416 7840 -2396 7874
rect -2362 7840 -2342 7874
rect -2416 7806 -2342 7840
rect -2416 7772 -2396 7806
rect -2362 7772 -2342 7806
rect -2416 7738 -2342 7772
rect -2416 7704 -2396 7738
rect -2362 7704 -2342 7738
rect -2416 7670 -2342 7704
rect -2416 7636 -2396 7670
rect -2362 7636 -2342 7670
rect -2416 7602 -2342 7636
rect -2416 7568 -2396 7602
rect -2362 7568 -2342 7602
rect -2416 7534 -2342 7568
rect -2416 7500 -2396 7534
rect -2362 7500 -2342 7534
rect -2416 7466 -2342 7500
rect -2416 7432 -2396 7466
rect -2362 7432 -2342 7466
rect -2416 7398 -2342 7432
rect -2416 7364 -2396 7398
rect -2362 7364 -2342 7398
rect -2416 7330 -2342 7364
rect -2416 7296 -2396 7330
rect -2362 7296 -2342 7330
rect -2416 7262 -2342 7296
rect -2416 7228 -2396 7262
rect -2362 7228 -2342 7262
rect -2416 7194 -2342 7228
rect -2416 7160 -2396 7194
rect -2362 7160 -2342 7194
rect -2416 7126 -2342 7160
rect -2416 7092 -2396 7126
rect -2362 7092 -2342 7126
rect -2416 7058 -2342 7092
rect -2416 7024 -2396 7058
rect -2362 7024 -2342 7058
rect -2416 6990 -2342 7024
rect -2416 6956 -2396 6990
rect -2362 6956 -2342 6990
rect -2416 6922 -2342 6956
rect -2416 6888 -2396 6922
rect -2362 6888 -2342 6922
rect -2416 6854 -2342 6888
rect -2416 6820 -2396 6854
rect -2362 6820 -2342 6854
rect -2416 6786 -2342 6820
rect -2416 6752 -2396 6786
rect -2362 6752 -2342 6786
rect -2416 6718 -2342 6752
rect -2416 6684 -2396 6718
rect -2362 6684 -2342 6718
rect -2416 6650 -2342 6684
rect -2416 6616 -2396 6650
rect -2362 6616 -2342 6650
rect -2416 6582 -2342 6616
rect -2416 6548 -2396 6582
rect -2362 6548 -2342 6582
rect -2416 6514 -2342 6548
rect -2416 6480 -2396 6514
rect -2362 6480 -2342 6514
rect -2416 6446 -2342 6480
rect -2416 6412 -2396 6446
rect -2362 6412 -2342 6446
rect -2416 6378 -2342 6412
rect -2416 6344 -2396 6378
rect -2362 6344 -2342 6378
rect -2416 6310 -2342 6344
rect -2416 6276 -2396 6310
rect -2362 6276 -2342 6310
rect -2416 6242 -2342 6276
rect -2416 6208 -2396 6242
rect -2362 6208 -2342 6242
rect -2416 6174 -2342 6208
rect -2416 6140 -2396 6174
rect -2362 6140 -2342 6174
rect -2416 6106 -2342 6140
rect -2416 6072 -2396 6106
rect -2362 6072 -2342 6106
rect -2416 6038 -2342 6072
rect -2416 6004 -2396 6038
rect -2362 6004 -2342 6038
rect -2416 5970 -2342 6004
rect -2416 5936 -2396 5970
rect -2362 5936 -2342 5970
rect -2416 5902 -2342 5936
rect -2416 5868 -2396 5902
rect -2362 5868 -2342 5902
rect -2416 5834 -2342 5868
rect -2416 5800 -2396 5834
rect -2362 5800 -2342 5834
rect -2416 5766 -2342 5800
rect -2416 5732 -2396 5766
rect -2362 5732 -2342 5766
rect -2416 5698 -2342 5732
rect -2416 5664 -2396 5698
rect -2362 5664 -2342 5698
rect -2416 5630 -2342 5664
rect -2416 5596 -2396 5630
rect -2362 5596 -2342 5630
rect -2416 5562 -2342 5596
rect -2416 5528 -2396 5562
rect -2362 5528 -2342 5562
rect -2416 5494 -2342 5528
rect -2416 5460 -2396 5494
rect -2362 5460 -2342 5494
rect -2416 5426 -2342 5460
rect -2416 5392 -2396 5426
rect -2362 5392 -2342 5426
rect -2416 5358 -2342 5392
rect -2416 5324 -2396 5358
rect -2362 5324 -2342 5358
rect -2416 5290 -2342 5324
rect -2416 5256 -2396 5290
rect -2362 5256 -2342 5290
rect -2416 5222 -2342 5256
rect -2416 5188 -2396 5222
rect -2362 5188 -2342 5222
rect -2416 5154 -2342 5188
rect -2416 5120 -2396 5154
rect -2362 5120 -2342 5154
rect -2416 5086 -2342 5120
rect -2416 5052 -2396 5086
rect -2362 5052 -2342 5086
rect -2416 5018 -2342 5052
rect -2416 4984 -2396 5018
rect -2362 4984 -2342 5018
rect -2416 4950 -2342 4984
rect -2416 4916 -2396 4950
rect -2362 4916 -2342 4950
rect -2416 4882 -2342 4916
rect -2416 4848 -2396 4882
rect -2362 4848 -2342 4882
rect -2416 4814 -2342 4848
rect -2416 4780 -2396 4814
rect -2362 4780 -2342 4814
rect -2416 4746 -2342 4780
rect -2416 4712 -2396 4746
rect -2362 4712 -2342 4746
rect -2416 4678 -2342 4712
rect -2416 4644 -2396 4678
rect -2362 4644 -2342 4678
rect -2416 4610 -2342 4644
rect -2416 4576 -2396 4610
rect -2362 4576 -2342 4610
rect -2416 4542 -2342 4576
rect -2416 4508 -2396 4542
rect -2362 4508 -2342 4542
rect -2416 4474 -2342 4508
rect -2416 4440 -2396 4474
rect -2362 4440 -2342 4474
rect -2416 4406 -2342 4440
rect -2416 4372 -2396 4406
rect -2362 4372 -2342 4406
rect -2416 4338 -2342 4372
rect -2416 4304 -2396 4338
rect -2362 4304 -2342 4338
rect -2416 4270 -2342 4304
rect -2416 4236 -2396 4270
rect -2362 4236 -2342 4270
rect -2416 4202 -2342 4236
rect -2416 4168 -2396 4202
rect -2362 4168 -2342 4202
rect -2416 4134 -2342 4168
rect -2416 4100 -2396 4134
rect -2362 4100 -2342 4134
rect -2416 4066 -2342 4100
rect -2416 4032 -2396 4066
rect -2362 4032 -2342 4066
rect -2416 3998 -2342 4032
rect -2416 3964 -2396 3998
rect -2362 3964 -2342 3998
rect -2416 3930 -2342 3964
rect -2416 3896 -2396 3930
rect -2362 3896 -2342 3930
rect -2416 3862 -2342 3896
rect -2416 3828 -2396 3862
rect -2362 3828 -2342 3862
rect -2416 3794 -2342 3828
rect -2416 3760 -2396 3794
rect -2362 3760 -2342 3794
rect -2416 3726 -2342 3760
rect -2416 3692 -2396 3726
rect -2362 3692 -2342 3726
rect -2416 3660 -2342 3692
rect 47176 19434 47250 19467
rect 47176 19400 47196 19434
rect 47230 19400 47250 19434
rect 47176 19366 47250 19400
rect 47176 19332 47196 19366
rect 47230 19332 47250 19366
rect 47176 19298 47250 19332
rect 47176 19264 47196 19298
rect 47230 19264 47250 19298
rect 47176 19230 47250 19264
rect 47176 19196 47196 19230
rect 47230 19196 47250 19230
rect 47176 19162 47250 19196
rect 47176 19128 47196 19162
rect 47230 19128 47250 19162
rect 47176 19094 47250 19128
rect 47176 19060 47196 19094
rect 47230 19060 47250 19094
rect 47176 19026 47250 19060
rect 47176 18992 47196 19026
rect 47230 18992 47250 19026
rect 47176 18958 47250 18992
rect 47176 18924 47196 18958
rect 47230 18924 47250 18958
rect 47176 18890 47250 18924
rect 47176 18856 47196 18890
rect 47230 18856 47250 18890
rect 47176 18822 47250 18856
rect 47176 18788 47196 18822
rect 47230 18788 47250 18822
rect 47176 18754 47250 18788
rect 47176 18720 47196 18754
rect 47230 18720 47250 18754
rect 47176 18686 47250 18720
rect 47176 18652 47196 18686
rect 47230 18652 47250 18686
rect 47176 18618 47250 18652
rect 47176 18584 47196 18618
rect 47230 18584 47250 18618
rect 47176 18550 47250 18584
rect 47176 18516 47196 18550
rect 47230 18516 47250 18550
rect 47176 18482 47250 18516
rect 47176 18448 47196 18482
rect 47230 18448 47250 18482
rect 47176 18414 47250 18448
rect 47176 18380 47196 18414
rect 47230 18380 47250 18414
rect 47176 18346 47250 18380
rect 47176 18312 47196 18346
rect 47230 18312 47250 18346
rect 47176 18278 47250 18312
rect 47176 18244 47196 18278
rect 47230 18244 47250 18278
rect 47176 18210 47250 18244
rect 47176 18176 47196 18210
rect 47230 18176 47250 18210
rect 47176 18142 47250 18176
rect 47176 18108 47196 18142
rect 47230 18108 47250 18142
rect 47176 18074 47250 18108
rect 47176 18040 47196 18074
rect 47230 18040 47250 18074
rect 47176 18006 47250 18040
rect 47176 17972 47196 18006
rect 47230 17972 47250 18006
rect 47176 17938 47250 17972
rect 47176 17904 47196 17938
rect 47230 17904 47250 17938
rect 47176 17870 47250 17904
rect 47176 17836 47196 17870
rect 47230 17836 47250 17870
rect 47176 17802 47250 17836
rect 47176 17768 47196 17802
rect 47230 17768 47250 17802
rect 47176 17734 47250 17768
rect 47176 17700 47196 17734
rect 47230 17700 47250 17734
rect 47176 17666 47250 17700
rect 47176 17632 47196 17666
rect 47230 17632 47250 17666
rect 47176 17598 47250 17632
rect 47176 17564 47196 17598
rect 47230 17564 47250 17598
rect 47176 17530 47250 17564
rect 47176 17496 47196 17530
rect 47230 17496 47250 17530
rect 47176 17462 47250 17496
rect 47176 17428 47196 17462
rect 47230 17428 47250 17462
rect 47176 17394 47250 17428
rect 47176 17360 47196 17394
rect 47230 17360 47250 17394
rect 47176 17326 47250 17360
rect 47176 17292 47196 17326
rect 47230 17292 47250 17326
rect 47176 17258 47250 17292
rect 47176 17224 47196 17258
rect 47230 17224 47250 17258
rect 47176 17190 47250 17224
rect 47176 17156 47196 17190
rect 47230 17156 47250 17190
rect 47176 17122 47250 17156
rect 47176 17088 47196 17122
rect 47230 17088 47250 17122
rect 47176 17054 47250 17088
rect 47176 17020 47196 17054
rect 47230 17020 47250 17054
rect 47176 16986 47250 17020
rect 47176 16952 47196 16986
rect 47230 16952 47250 16986
rect 47176 16918 47250 16952
rect 47176 16884 47196 16918
rect 47230 16884 47250 16918
rect 47176 16850 47250 16884
rect 47176 16816 47196 16850
rect 47230 16816 47250 16850
rect 47176 16782 47250 16816
rect 47176 16748 47196 16782
rect 47230 16748 47250 16782
rect 47176 16714 47250 16748
rect 47176 16680 47196 16714
rect 47230 16680 47250 16714
rect 47176 16646 47250 16680
rect 47176 16612 47196 16646
rect 47230 16612 47250 16646
rect 47176 16578 47250 16612
rect 47176 16544 47196 16578
rect 47230 16544 47250 16578
rect 47176 16510 47250 16544
rect 47176 16476 47196 16510
rect 47230 16476 47250 16510
rect 47176 16442 47250 16476
rect 47176 16408 47196 16442
rect 47230 16408 47250 16442
rect 47176 16374 47250 16408
rect 47176 16340 47196 16374
rect 47230 16340 47250 16374
rect 47176 16306 47250 16340
rect 47176 16272 47196 16306
rect 47230 16272 47250 16306
rect 47176 16238 47250 16272
rect 47176 16204 47196 16238
rect 47230 16204 47250 16238
rect 47176 16170 47250 16204
rect 47176 16136 47196 16170
rect 47230 16136 47250 16170
rect 47176 16102 47250 16136
rect 47176 16068 47196 16102
rect 47230 16068 47250 16102
rect 47176 16034 47250 16068
rect 47176 16000 47196 16034
rect 47230 16000 47250 16034
rect 47176 15966 47250 16000
rect 47176 15932 47196 15966
rect 47230 15932 47250 15966
rect 47176 15898 47250 15932
rect 47176 15864 47196 15898
rect 47230 15864 47250 15898
rect 47176 15830 47250 15864
rect 47176 15796 47196 15830
rect 47230 15796 47250 15830
rect 47176 15762 47250 15796
rect 47176 15728 47196 15762
rect 47230 15728 47250 15762
rect 47176 15694 47250 15728
rect 47176 15660 47196 15694
rect 47230 15660 47250 15694
rect 47176 15626 47250 15660
rect 47176 15592 47196 15626
rect 47230 15592 47250 15626
rect 47176 15558 47250 15592
rect 47176 15524 47196 15558
rect 47230 15524 47250 15558
rect 47176 15490 47250 15524
rect 47176 15456 47196 15490
rect 47230 15456 47250 15490
rect 47176 15422 47250 15456
rect 47176 15388 47196 15422
rect 47230 15388 47250 15422
rect 47176 15354 47250 15388
rect 47176 15320 47196 15354
rect 47230 15320 47250 15354
rect 47176 15286 47250 15320
rect 47176 15252 47196 15286
rect 47230 15252 47250 15286
rect 47176 15218 47250 15252
rect 47176 15184 47196 15218
rect 47230 15184 47250 15218
rect 47176 15150 47250 15184
rect 47176 15116 47196 15150
rect 47230 15116 47250 15150
rect 47176 15082 47250 15116
rect 47176 15048 47196 15082
rect 47230 15048 47250 15082
rect 47176 15014 47250 15048
rect 47176 14980 47196 15014
rect 47230 14980 47250 15014
rect 47176 14946 47250 14980
rect 47176 14912 47196 14946
rect 47230 14912 47250 14946
rect 47176 14878 47250 14912
rect 47176 14844 47196 14878
rect 47230 14844 47250 14878
rect 47176 14810 47250 14844
rect 47176 14776 47196 14810
rect 47230 14776 47250 14810
rect 47176 14742 47250 14776
rect 47176 14708 47196 14742
rect 47230 14708 47250 14742
rect 47176 14674 47250 14708
rect 47176 14640 47196 14674
rect 47230 14640 47250 14674
rect 47176 14606 47250 14640
rect 47176 14572 47196 14606
rect 47230 14572 47250 14606
rect 47176 14538 47250 14572
rect 47176 14504 47196 14538
rect 47230 14504 47250 14538
rect 47176 14470 47250 14504
rect 47176 14436 47196 14470
rect 47230 14436 47250 14470
rect 47176 14402 47250 14436
rect 47176 14368 47196 14402
rect 47230 14368 47250 14402
rect 47176 14334 47250 14368
rect 47176 14300 47196 14334
rect 47230 14300 47250 14334
rect 47176 14266 47250 14300
rect 47176 14232 47196 14266
rect 47230 14232 47250 14266
rect 47176 14198 47250 14232
rect 47176 14164 47196 14198
rect 47230 14164 47250 14198
rect 47176 14130 47250 14164
rect 47176 14096 47196 14130
rect 47230 14096 47250 14130
rect 47176 14062 47250 14096
rect 47176 14028 47196 14062
rect 47230 14028 47250 14062
rect 47176 13994 47250 14028
rect 47176 13960 47196 13994
rect 47230 13960 47250 13994
rect 47176 13926 47250 13960
rect 47176 13892 47196 13926
rect 47230 13892 47250 13926
rect 47176 13858 47250 13892
rect 47176 13824 47196 13858
rect 47230 13824 47250 13858
rect 47176 13790 47250 13824
rect 47176 13756 47196 13790
rect 47230 13756 47250 13790
rect 47176 13722 47250 13756
rect 47176 13688 47196 13722
rect 47230 13688 47250 13722
rect 47176 13654 47250 13688
rect 47176 13620 47196 13654
rect 47230 13620 47250 13654
rect 47176 13586 47250 13620
rect 47176 13552 47196 13586
rect 47230 13552 47250 13586
rect 47176 13518 47250 13552
rect 47176 13484 47196 13518
rect 47230 13484 47250 13518
rect 47176 13450 47250 13484
rect 47176 13416 47196 13450
rect 47230 13416 47250 13450
rect 47176 13382 47250 13416
rect 47176 13348 47196 13382
rect 47230 13348 47250 13382
rect 47176 13314 47250 13348
rect 47176 13280 47196 13314
rect 47230 13280 47250 13314
rect 47176 13246 47250 13280
rect 47176 13212 47196 13246
rect 47230 13212 47250 13246
rect 47176 13178 47250 13212
rect 47176 13144 47196 13178
rect 47230 13144 47250 13178
rect 47176 13110 47250 13144
rect 47176 13076 47196 13110
rect 47230 13076 47250 13110
rect 47176 13042 47250 13076
rect 47176 13008 47196 13042
rect 47230 13008 47250 13042
rect 47176 12974 47250 13008
rect 47176 12940 47196 12974
rect 47230 12940 47250 12974
rect 47176 12906 47250 12940
rect 47176 12872 47196 12906
rect 47230 12872 47250 12906
rect 47176 12838 47250 12872
rect 47176 12804 47196 12838
rect 47230 12804 47250 12838
rect 47176 12770 47250 12804
rect 47176 12736 47196 12770
rect 47230 12736 47250 12770
rect 47176 12702 47250 12736
rect 47176 12668 47196 12702
rect 47230 12668 47250 12702
rect 47176 12634 47250 12668
rect 47176 12600 47196 12634
rect 47230 12600 47250 12634
rect 47176 12566 47250 12600
rect 47176 12532 47196 12566
rect 47230 12532 47250 12566
rect 47176 12498 47250 12532
rect 47176 12464 47196 12498
rect 47230 12464 47250 12498
rect 47176 12430 47250 12464
rect 47176 12396 47196 12430
rect 47230 12396 47250 12430
rect 47176 12362 47250 12396
rect 47176 12328 47196 12362
rect 47230 12328 47250 12362
rect 47176 12294 47250 12328
rect 47176 12260 47196 12294
rect 47230 12260 47250 12294
rect 47176 12226 47250 12260
rect 47176 12192 47196 12226
rect 47230 12192 47250 12226
rect 47176 12158 47250 12192
rect 47176 12124 47196 12158
rect 47230 12124 47250 12158
rect 47176 12090 47250 12124
rect 47176 12056 47196 12090
rect 47230 12056 47250 12090
rect 47176 12022 47250 12056
rect 47176 11988 47196 12022
rect 47230 11988 47250 12022
rect 47176 11954 47250 11988
rect 47176 11920 47196 11954
rect 47230 11920 47250 11954
rect 47176 11886 47250 11920
rect 47176 11852 47196 11886
rect 47230 11852 47250 11886
rect 47176 11818 47250 11852
rect 47176 11784 47196 11818
rect 47230 11784 47250 11818
rect 47176 11750 47250 11784
rect 47176 11716 47196 11750
rect 47230 11716 47250 11750
rect 47176 11682 47250 11716
rect 47176 11648 47196 11682
rect 47230 11648 47250 11682
rect 47176 11614 47250 11648
rect 47176 11580 47196 11614
rect 47230 11580 47250 11614
rect 47176 11546 47250 11580
rect 47176 11512 47196 11546
rect 47230 11512 47250 11546
rect 47176 11478 47250 11512
rect 47176 11444 47196 11478
rect 47230 11444 47250 11478
rect 47176 11410 47250 11444
rect 47176 11376 47196 11410
rect 47230 11376 47250 11410
rect 47176 11342 47250 11376
rect 47176 11308 47196 11342
rect 47230 11308 47250 11342
rect 47176 11274 47250 11308
rect 47176 11240 47196 11274
rect 47230 11240 47250 11274
rect 47176 11206 47250 11240
rect 47176 11172 47196 11206
rect 47230 11172 47250 11206
rect 47176 11138 47250 11172
rect 47176 11104 47196 11138
rect 47230 11104 47250 11138
rect 47176 11070 47250 11104
rect 47176 11036 47196 11070
rect 47230 11036 47250 11070
rect 47176 11002 47250 11036
rect 47176 10968 47196 11002
rect 47230 10968 47250 11002
rect 47176 10934 47250 10968
rect 47176 10900 47196 10934
rect 47230 10900 47250 10934
rect 47176 10866 47250 10900
rect 47176 10832 47196 10866
rect 47230 10832 47250 10866
rect 47176 10798 47250 10832
rect 47176 10764 47196 10798
rect 47230 10764 47250 10798
rect 47176 10730 47250 10764
rect 47176 10696 47196 10730
rect 47230 10696 47250 10730
rect 47176 10662 47250 10696
rect 47176 10628 47196 10662
rect 47230 10628 47250 10662
rect 47176 10594 47250 10628
rect 47176 10560 47196 10594
rect 47230 10560 47250 10594
rect 47176 10526 47250 10560
rect 47176 10492 47196 10526
rect 47230 10492 47250 10526
rect 47176 10458 47250 10492
rect 47176 10424 47196 10458
rect 47230 10424 47250 10458
rect 47176 10390 47250 10424
rect 47176 10356 47196 10390
rect 47230 10356 47250 10390
rect 47176 10322 47250 10356
rect 47176 10288 47196 10322
rect 47230 10288 47250 10322
rect 47176 10254 47250 10288
rect 47176 10220 47196 10254
rect 47230 10220 47250 10254
rect 47176 10186 47250 10220
rect 47176 10152 47196 10186
rect 47230 10152 47250 10186
rect 47176 10118 47250 10152
rect 47176 10084 47196 10118
rect 47230 10084 47250 10118
rect 47176 10050 47250 10084
rect 47176 10016 47196 10050
rect 47230 10016 47250 10050
rect 47176 9982 47250 10016
rect 47176 9948 47196 9982
rect 47230 9948 47250 9982
rect 47176 9914 47250 9948
rect 47176 9880 47196 9914
rect 47230 9880 47250 9914
rect 47176 9846 47250 9880
rect 47176 9812 47196 9846
rect 47230 9812 47250 9846
rect 47176 9778 47250 9812
rect 47176 9744 47196 9778
rect 47230 9744 47250 9778
rect 47176 9710 47250 9744
rect 47176 9676 47196 9710
rect 47230 9676 47250 9710
rect 47176 9642 47250 9676
rect 47176 9608 47196 9642
rect 47230 9608 47250 9642
rect 47176 9574 47250 9608
rect 47176 9540 47196 9574
rect 47230 9540 47250 9574
rect 47176 9506 47250 9540
rect 47176 9472 47196 9506
rect 47230 9472 47250 9506
rect 47176 9438 47250 9472
rect 47176 9404 47196 9438
rect 47230 9404 47250 9438
rect 47176 9370 47250 9404
rect 47176 9336 47196 9370
rect 47230 9336 47250 9370
rect 47176 9302 47250 9336
rect 47176 9268 47196 9302
rect 47230 9268 47250 9302
rect 47176 9234 47250 9268
rect 47176 9200 47196 9234
rect 47230 9200 47250 9234
rect 47176 9166 47250 9200
rect 47176 9132 47196 9166
rect 47230 9132 47250 9166
rect 47176 9098 47250 9132
rect 47176 9064 47196 9098
rect 47230 9064 47250 9098
rect 47176 9030 47250 9064
rect 47176 8996 47196 9030
rect 47230 8996 47250 9030
rect 47176 8962 47250 8996
rect 47176 8928 47196 8962
rect 47230 8928 47250 8962
rect 47176 8894 47250 8928
rect 47176 8860 47196 8894
rect 47230 8860 47250 8894
rect 47176 8826 47250 8860
rect 47176 8792 47196 8826
rect 47230 8792 47250 8826
rect 47176 8758 47250 8792
rect 47176 8724 47196 8758
rect 47230 8724 47250 8758
rect 47176 8690 47250 8724
rect 47176 8656 47196 8690
rect 47230 8656 47250 8690
rect 47176 8622 47250 8656
rect 47176 8588 47196 8622
rect 47230 8588 47250 8622
rect 47176 8554 47250 8588
rect 47176 8520 47196 8554
rect 47230 8520 47250 8554
rect 47176 8486 47250 8520
rect 47176 8452 47196 8486
rect 47230 8452 47250 8486
rect 47176 8418 47250 8452
rect 47176 8384 47196 8418
rect 47230 8384 47250 8418
rect 47176 8350 47250 8384
rect 47176 8316 47196 8350
rect 47230 8316 47250 8350
rect 47176 8282 47250 8316
rect 47176 8248 47196 8282
rect 47230 8248 47250 8282
rect 47176 8214 47250 8248
rect 47176 8180 47196 8214
rect 47230 8180 47250 8214
rect 47176 8146 47250 8180
rect 47176 8112 47196 8146
rect 47230 8112 47250 8146
rect 47176 8078 47250 8112
rect 47176 8044 47196 8078
rect 47230 8044 47250 8078
rect 47176 8010 47250 8044
rect 47176 7976 47196 8010
rect 47230 7976 47250 8010
rect 47176 7942 47250 7976
rect 47176 7908 47196 7942
rect 47230 7908 47250 7942
rect 47176 7874 47250 7908
rect 47176 7840 47196 7874
rect 47230 7840 47250 7874
rect 47176 7806 47250 7840
rect 47176 7772 47196 7806
rect 47230 7772 47250 7806
rect 47176 7738 47250 7772
rect 47176 7704 47196 7738
rect 47230 7704 47250 7738
rect 47176 7670 47250 7704
rect 47176 7636 47196 7670
rect 47230 7636 47250 7670
rect 47176 7602 47250 7636
rect 47176 7568 47196 7602
rect 47230 7568 47250 7602
rect 47176 7534 47250 7568
rect 47176 7500 47196 7534
rect 47230 7500 47250 7534
rect 47176 7466 47250 7500
rect 47176 7432 47196 7466
rect 47230 7432 47250 7466
rect 47176 7398 47250 7432
rect 47176 7364 47196 7398
rect 47230 7364 47250 7398
rect 47176 7330 47250 7364
rect 47176 7296 47196 7330
rect 47230 7296 47250 7330
rect 47176 7262 47250 7296
rect 47176 7228 47196 7262
rect 47230 7228 47250 7262
rect 47176 7194 47250 7228
rect 47176 7160 47196 7194
rect 47230 7160 47250 7194
rect 47176 7126 47250 7160
rect 47176 7092 47196 7126
rect 47230 7092 47250 7126
rect 47176 7058 47250 7092
rect 47176 7024 47196 7058
rect 47230 7024 47250 7058
rect 47176 6990 47250 7024
rect 47176 6956 47196 6990
rect 47230 6956 47250 6990
rect 47176 6922 47250 6956
rect 47176 6888 47196 6922
rect 47230 6888 47250 6922
rect 47176 6854 47250 6888
rect 47176 6820 47196 6854
rect 47230 6820 47250 6854
rect 47176 6786 47250 6820
rect 47176 6752 47196 6786
rect 47230 6752 47250 6786
rect 47176 6718 47250 6752
rect 47176 6684 47196 6718
rect 47230 6684 47250 6718
rect 47176 6650 47250 6684
rect 47176 6616 47196 6650
rect 47230 6616 47250 6650
rect 47176 6582 47250 6616
rect 47176 6548 47196 6582
rect 47230 6548 47250 6582
rect 47176 6514 47250 6548
rect 47176 6480 47196 6514
rect 47230 6480 47250 6514
rect 47176 6446 47250 6480
rect 47176 6412 47196 6446
rect 47230 6412 47250 6446
rect 47176 6378 47250 6412
rect 47176 6344 47196 6378
rect 47230 6344 47250 6378
rect 47176 6310 47250 6344
rect 47176 6276 47196 6310
rect 47230 6276 47250 6310
rect 47176 6242 47250 6276
rect 47176 6208 47196 6242
rect 47230 6208 47250 6242
rect 47176 6174 47250 6208
rect 47176 6140 47196 6174
rect 47230 6140 47250 6174
rect 47176 6106 47250 6140
rect 47176 6072 47196 6106
rect 47230 6072 47250 6106
rect 47176 6038 47250 6072
rect 47176 6004 47196 6038
rect 47230 6004 47250 6038
rect 47176 5970 47250 6004
rect 47176 5936 47196 5970
rect 47230 5936 47250 5970
rect 47176 5902 47250 5936
rect 47176 5868 47196 5902
rect 47230 5868 47250 5902
rect 47176 5834 47250 5868
rect 47176 5800 47196 5834
rect 47230 5800 47250 5834
rect 47176 5766 47250 5800
rect 47176 5732 47196 5766
rect 47230 5732 47250 5766
rect 47176 5698 47250 5732
rect 47176 5664 47196 5698
rect 47230 5664 47250 5698
rect 47176 5630 47250 5664
rect 47176 5596 47196 5630
rect 47230 5596 47250 5630
rect 47176 5562 47250 5596
rect 47176 5528 47196 5562
rect 47230 5528 47250 5562
rect 47176 5494 47250 5528
rect 47176 5460 47196 5494
rect 47230 5460 47250 5494
rect 47176 5426 47250 5460
rect 47176 5392 47196 5426
rect 47230 5392 47250 5426
rect 47176 5358 47250 5392
rect 47176 5324 47196 5358
rect 47230 5324 47250 5358
rect 47176 5290 47250 5324
rect 47176 5256 47196 5290
rect 47230 5256 47250 5290
rect 47176 5222 47250 5256
rect 47176 5188 47196 5222
rect 47230 5188 47250 5222
rect 47176 5154 47250 5188
rect 47176 5120 47196 5154
rect 47230 5120 47250 5154
rect 47176 5086 47250 5120
rect 47176 5052 47196 5086
rect 47230 5052 47250 5086
rect 47176 5018 47250 5052
rect 47176 4984 47196 5018
rect 47230 4984 47250 5018
rect 47176 4950 47250 4984
rect 47176 4916 47196 4950
rect 47230 4916 47250 4950
rect 47176 4882 47250 4916
rect 47176 4848 47196 4882
rect 47230 4848 47250 4882
rect 47176 4814 47250 4848
rect 47176 4780 47196 4814
rect 47230 4780 47250 4814
rect 47176 4746 47250 4780
rect 47176 4712 47196 4746
rect 47230 4712 47250 4746
rect 47176 4678 47250 4712
rect 47176 4644 47196 4678
rect 47230 4644 47250 4678
rect 47176 4610 47250 4644
rect 47176 4576 47196 4610
rect 47230 4576 47250 4610
rect 47176 4542 47250 4576
rect 47176 4508 47196 4542
rect 47230 4508 47250 4542
rect 47176 4474 47250 4508
rect 47176 4440 47196 4474
rect 47230 4440 47250 4474
rect 47176 4406 47250 4440
rect 47176 4372 47196 4406
rect 47230 4372 47250 4406
rect 47176 4338 47250 4372
rect 47176 4304 47196 4338
rect 47230 4304 47250 4338
rect 47176 4270 47250 4304
rect 47176 4236 47196 4270
rect 47230 4236 47250 4270
rect 47176 4202 47250 4236
rect 47176 4168 47196 4202
rect 47230 4168 47250 4202
rect 47176 4134 47250 4168
rect 47176 4100 47196 4134
rect 47230 4100 47250 4134
rect 47176 4066 47250 4100
rect 47176 4032 47196 4066
rect 47230 4032 47250 4066
rect 47176 3998 47250 4032
rect 47176 3964 47196 3998
rect 47230 3964 47250 3998
rect 47176 3930 47250 3964
rect 47176 3896 47196 3930
rect 47230 3896 47250 3930
rect 47176 3862 47250 3896
rect 47176 3828 47196 3862
rect 47230 3828 47250 3862
rect 47176 3794 47250 3828
rect 47176 3760 47196 3794
rect 47230 3760 47250 3794
rect 47176 3726 47250 3760
rect 47176 3692 47196 3726
rect 47230 3692 47250 3726
rect 47176 3660 47250 3692
rect -2416 3640 47250 3660
rect -2416 3606 -2318 3640
rect -2284 3606 -2250 3640
rect -2216 3606 -2182 3640
rect -2148 3606 -2114 3640
rect -2080 3606 -2046 3640
rect -2012 3606 -1978 3640
rect -1944 3606 -1910 3640
rect -1876 3606 -1842 3640
rect -1808 3606 -1774 3640
rect -1740 3606 -1706 3640
rect -1672 3606 -1638 3640
rect -1604 3606 -1570 3640
rect -1536 3606 -1502 3640
rect -1468 3606 -1434 3640
rect -1400 3606 -1366 3640
rect -1332 3606 -1298 3640
rect -1264 3606 -1230 3640
rect -1196 3606 -1162 3640
rect -1128 3606 -1094 3640
rect -1060 3606 -1026 3640
rect -992 3606 -958 3640
rect -924 3606 -890 3640
rect -856 3606 -822 3640
rect -788 3606 -754 3640
rect -720 3606 -686 3640
rect -652 3606 -618 3640
rect -584 3606 -550 3640
rect -516 3606 -482 3640
rect -448 3606 -414 3640
rect -380 3606 -346 3640
rect -312 3606 -278 3640
rect -244 3606 -210 3640
rect -176 3606 -142 3640
rect -108 3606 -74 3640
rect -40 3606 -6 3640
rect 28 3606 62 3640
rect 96 3606 130 3640
rect 164 3606 198 3640
rect 232 3606 266 3640
rect 300 3606 334 3640
rect 368 3606 402 3640
rect 436 3606 470 3640
rect 504 3606 538 3640
rect 572 3606 606 3640
rect 640 3606 674 3640
rect 708 3606 742 3640
rect 776 3606 810 3640
rect 844 3606 878 3640
rect 912 3606 946 3640
rect 980 3606 1014 3640
rect 1048 3606 1082 3640
rect 1116 3606 1150 3640
rect 1184 3606 1218 3640
rect 1252 3606 1286 3640
rect 1320 3606 1354 3640
rect 1388 3606 1422 3640
rect 1456 3606 1490 3640
rect 1524 3606 1558 3640
rect 1592 3606 1626 3640
rect 1660 3606 1694 3640
rect 1728 3606 1762 3640
rect 1796 3606 1830 3640
rect 1864 3606 1898 3640
rect 1932 3606 1966 3640
rect 2000 3606 2034 3640
rect 2068 3606 2102 3640
rect 2136 3606 2170 3640
rect 2204 3606 2238 3640
rect 2272 3606 2306 3640
rect 2340 3606 2374 3640
rect 2408 3606 2442 3640
rect 2476 3606 2510 3640
rect 2544 3606 2578 3640
rect 2612 3606 2646 3640
rect 2680 3606 2714 3640
rect 2748 3606 2782 3640
rect 2816 3606 2850 3640
rect 2884 3606 2918 3640
rect 2952 3606 2986 3640
rect 3020 3606 3054 3640
rect 3088 3606 3122 3640
rect 3156 3606 3190 3640
rect 3224 3606 3258 3640
rect 3292 3606 3326 3640
rect 3360 3606 3394 3640
rect 3428 3606 3462 3640
rect 3496 3606 3530 3640
rect 3564 3606 3598 3640
rect 3632 3606 3666 3640
rect 3700 3606 3734 3640
rect 3768 3606 3802 3640
rect 3836 3606 3870 3640
rect 3904 3606 3938 3640
rect 3972 3606 4006 3640
rect 4040 3606 4074 3640
rect 4108 3606 4142 3640
rect 4176 3606 4210 3640
rect 4244 3606 4278 3640
rect 4312 3606 4346 3640
rect 4380 3606 4414 3640
rect 4448 3606 4482 3640
rect 4516 3606 4550 3640
rect 4584 3606 4618 3640
rect 4652 3606 4686 3640
rect 4720 3606 4754 3640
rect 4788 3606 4822 3640
rect 4856 3606 4890 3640
rect 4924 3606 4958 3640
rect 4992 3606 5026 3640
rect 5060 3606 5094 3640
rect 5128 3606 5162 3640
rect 5196 3606 5230 3640
rect 5264 3606 5298 3640
rect 5332 3606 5366 3640
rect 5400 3606 5434 3640
rect 5468 3606 5502 3640
rect 5536 3606 5570 3640
rect 5604 3606 5638 3640
rect 5672 3606 5706 3640
rect 5740 3606 5774 3640
rect 5808 3606 5842 3640
rect 5876 3606 5910 3640
rect 5944 3606 5978 3640
rect 6012 3606 6046 3640
rect 6080 3606 6114 3640
rect 6148 3606 6182 3640
rect 6216 3606 6250 3640
rect 6284 3606 6318 3640
rect 6352 3606 6386 3640
rect 6420 3606 6454 3640
rect 6488 3606 6522 3640
rect 6556 3606 6590 3640
rect 6624 3606 6658 3640
rect 6692 3606 6726 3640
rect 6760 3606 6794 3640
rect 6828 3606 6862 3640
rect 6896 3606 6930 3640
rect 6964 3606 6998 3640
rect 7032 3606 7066 3640
rect 7100 3606 7134 3640
rect 7168 3606 7202 3640
rect 7236 3606 7270 3640
rect 7304 3606 7338 3640
rect 7372 3606 7406 3640
rect 7440 3606 7474 3640
rect 7508 3606 7542 3640
rect 7576 3606 7610 3640
rect 7644 3606 7678 3640
rect 7712 3606 7746 3640
rect 7780 3606 7814 3640
rect 7848 3606 7882 3640
rect 7916 3606 7950 3640
rect 7984 3606 8018 3640
rect 8052 3606 8086 3640
rect 8120 3606 8154 3640
rect 8188 3606 8222 3640
rect 8256 3606 8290 3640
rect 8324 3606 8358 3640
rect 8392 3606 8426 3640
rect 8460 3606 8494 3640
rect 8528 3606 8562 3640
rect 8596 3606 8630 3640
rect 8664 3606 8698 3640
rect 8732 3606 8766 3640
rect 8800 3606 8834 3640
rect 8868 3606 8902 3640
rect 8936 3606 8970 3640
rect 9004 3606 9038 3640
rect 9072 3606 9106 3640
rect 9140 3606 9174 3640
rect 9208 3606 9242 3640
rect 9276 3606 9310 3640
rect 9344 3606 9378 3640
rect 9412 3606 9446 3640
rect 9480 3606 9514 3640
rect 9548 3606 9582 3640
rect 9616 3606 9650 3640
rect 9684 3606 9718 3640
rect 9752 3606 9786 3640
rect 9820 3606 9854 3640
rect 9888 3606 9922 3640
rect 9956 3606 9990 3640
rect 10024 3606 10058 3640
rect 10092 3606 10126 3640
rect 10160 3606 10194 3640
rect 10228 3606 10262 3640
rect 10296 3606 10330 3640
rect 10364 3606 10398 3640
rect 10432 3606 10466 3640
rect 10500 3606 10534 3640
rect 10568 3606 10602 3640
rect 10636 3606 10670 3640
rect 10704 3606 10738 3640
rect 10772 3606 10806 3640
rect 10840 3606 10874 3640
rect 10908 3606 10942 3640
rect 10976 3606 11010 3640
rect 11044 3606 11078 3640
rect 11112 3606 11146 3640
rect 11180 3606 11214 3640
rect 11248 3606 11282 3640
rect 11316 3606 11350 3640
rect 11384 3606 11418 3640
rect 11452 3606 11486 3640
rect 11520 3606 11554 3640
rect 11588 3606 11622 3640
rect 11656 3606 11690 3640
rect 11724 3606 11758 3640
rect 11792 3606 11826 3640
rect 11860 3606 11894 3640
rect 11928 3606 11962 3640
rect 11996 3606 12030 3640
rect 12064 3606 12098 3640
rect 12132 3606 12166 3640
rect 12200 3606 12234 3640
rect 12268 3606 12302 3640
rect 12336 3606 12370 3640
rect 12404 3606 12438 3640
rect 12472 3606 12506 3640
rect 12540 3606 12574 3640
rect 12608 3606 12642 3640
rect 12676 3606 12710 3640
rect 12744 3606 12778 3640
rect 12812 3606 12846 3640
rect 12880 3606 12914 3640
rect 12948 3606 12982 3640
rect 13016 3606 13050 3640
rect 13084 3606 13118 3640
rect 13152 3606 13186 3640
rect 13220 3606 13254 3640
rect 13288 3606 13322 3640
rect 13356 3606 13390 3640
rect 13424 3606 13458 3640
rect 13492 3606 13526 3640
rect 13560 3606 13594 3640
rect 13628 3606 13662 3640
rect 13696 3606 13730 3640
rect 13764 3606 13798 3640
rect 13832 3606 13866 3640
rect 13900 3606 13934 3640
rect 13968 3606 14002 3640
rect 14036 3606 14070 3640
rect 14104 3606 14138 3640
rect 14172 3606 14206 3640
rect 14240 3606 14274 3640
rect 14308 3606 14342 3640
rect 14376 3606 14410 3640
rect 14444 3606 14478 3640
rect 14512 3606 14546 3640
rect 14580 3606 14614 3640
rect 14648 3606 14682 3640
rect 14716 3606 14750 3640
rect 14784 3606 14818 3640
rect 14852 3606 14886 3640
rect 14920 3606 14954 3640
rect 14988 3606 15022 3640
rect 15056 3606 15090 3640
rect 15124 3606 15158 3640
rect 15192 3606 15226 3640
rect 15260 3606 15294 3640
rect 15328 3606 15362 3640
rect 15396 3606 15430 3640
rect 15464 3606 15498 3640
rect 15532 3606 15566 3640
rect 15600 3606 15634 3640
rect 15668 3606 15702 3640
rect 15736 3606 15770 3640
rect 15804 3606 15838 3640
rect 15872 3606 15906 3640
rect 15940 3606 15974 3640
rect 16008 3606 16042 3640
rect 16076 3606 16110 3640
rect 16144 3606 16178 3640
rect 16212 3606 16246 3640
rect 16280 3606 16314 3640
rect 16348 3606 16382 3640
rect 16416 3606 16450 3640
rect 16484 3606 16518 3640
rect 16552 3606 16586 3640
rect 16620 3606 16654 3640
rect 16688 3606 16722 3640
rect 16756 3606 16790 3640
rect 16824 3606 16858 3640
rect 16892 3606 16926 3640
rect 16960 3606 16994 3640
rect 17028 3606 17062 3640
rect 17096 3606 17130 3640
rect 17164 3606 17198 3640
rect 17232 3606 17266 3640
rect 17300 3606 17334 3640
rect 17368 3606 17402 3640
rect 17436 3606 17470 3640
rect 17504 3606 17538 3640
rect 17572 3606 17606 3640
rect 17640 3606 17674 3640
rect 17708 3606 17742 3640
rect 17776 3606 17810 3640
rect 17844 3606 17878 3640
rect 17912 3606 17946 3640
rect 17980 3606 18014 3640
rect 18048 3606 18082 3640
rect 18116 3606 18150 3640
rect 18184 3606 18218 3640
rect 18252 3606 18286 3640
rect 18320 3606 18354 3640
rect 18388 3606 18422 3640
rect 18456 3606 18490 3640
rect 18524 3606 18558 3640
rect 18592 3606 18626 3640
rect 18660 3606 18694 3640
rect 18728 3606 18762 3640
rect 18796 3606 18830 3640
rect 18864 3606 18898 3640
rect 18932 3606 18966 3640
rect 19000 3606 19034 3640
rect 19068 3606 19102 3640
rect 19136 3606 19170 3640
rect 19204 3606 19238 3640
rect 19272 3606 19306 3640
rect 19340 3606 19374 3640
rect 19408 3606 19442 3640
rect 19476 3606 19510 3640
rect 19544 3606 19578 3640
rect 19612 3606 19646 3640
rect 19680 3606 19714 3640
rect 19748 3606 19782 3640
rect 19816 3606 19850 3640
rect 19884 3606 19918 3640
rect 19952 3606 19986 3640
rect 20020 3606 20054 3640
rect 20088 3606 20122 3640
rect 20156 3606 20190 3640
rect 20224 3606 20258 3640
rect 20292 3606 20326 3640
rect 20360 3606 20394 3640
rect 20428 3606 20462 3640
rect 20496 3606 20530 3640
rect 20564 3606 20598 3640
rect 20632 3606 20666 3640
rect 20700 3606 20734 3640
rect 20768 3606 20802 3640
rect 20836 3606 20870 3640
rect 20904 3606 20938 3640
rect 20972 3606 21006 3640
rect 21040 3606 21074 3640
rect 21108 3606 21142 3640
rect 21176 3606 21210 3640
rect 21244 3606 21278 3640
rect 21312 3606 21346 3640
rect 21380 3606 21414 3640
rect 21448 3606 21482 3640
rect 21516 3606 21550 3640
rect 21584 3606 21618 3640
rect 21652 3606 21686 3640
rect 21720 3606 21754 3640
rect 21788 3606 21822 3640
rect 21856 3606 21890 3640
rect 21924 3606 21958 3640
rect 21992 3606 22026 3640
rect 22060 3606 22094 3640
rect 22128 3606 22162 3640
rect 22196 3606 22230 3640
rect 22264 3606 22298 3640
rect 22332 3606 22366 3640
rect 22400 3606 22434 3640
rect 22468 3606 22502 3640
rect 22536 3606 22570 3640
rect 22604 3606 22638 3640
rect 22672 3606 22706 3640
rect 22740 3606 22774 3640
rect 22808 3606 22842 3640
rect 22876 3606 22910 3640
rect 22944 3606 22978 3640
rect 23012 3606 23046 3640
rect 23080 3606 23114 3640
rect 23148 3606 23182 3640
rect 23216 3606 23250 3640
rect 23284 3606 23318 3640
rect 23352 3606 23386 3640
rect 23420 3606 23454 3640
rect 23488 3606 23522 3640
rect 23556 3606 23590 3640
rect 23624 3606 23658 3640
rect 23692 3606 23726 3640
rect 23760 3606 23794 3640
rect 23828 3606 23862 3640
rect 23896 3606 23930 3640
rect 23964 3606 23998 3640
rect 24032 3606 24066 3640
rect 24100 3606 24134 3640
rect 24168 3606 24202 3640
rect 24236 3606 24270 3640
rect 24304 3606 24338 3640
rect 24372 3606 24406 3640
rect 24440 3606 24474 3640
rect 24508 3606 24542 3640
rect 24576 3606 24610 3640
rect 24644 3606 24678 3640
rect 24712 3606 24746 3640
rect 24780 3606 24814 3640
rect 24848 3606 24882 3640
rect 24916 3606 24950 3640
rect 24984 3606 25018 3640
rect 25052 3606 25086 3640
rect 25120 3606 25154 3640
rect 25188 3606 25222 3640
rect 25256 3606 25290 3640
rect 25324 3606 25358 3640
rect 25392 3606 25426 3640
rect 25460 3606 25494 3640
rect 25528 3606 25562 3640
rect 25596 3606 25630 3640
rect 25664 3606 25698 3640
rect 25732 3606 25766 3640
rect 25800 3606 25834 3640
rect 25868 3606 25902 3640
rect 25936 3606 25970 3640
rect 26004 3606 26038 3640
rect 26072 3606 26106 3640
rect 26140 3606 26174 3640
rect 26208 3606 26242 3640
rect 26276 3606 26310 3640
rect 26344 3606 26378 3640
rect 26412 3606 26446 3640
rect 26480 3606 26514 3640
rect 26548 3606 26582 3640
rect 26616 3606 26650 3640
rect 26684 3606 26718 3640
rect 26752 3606 26786 3640
rect 26820 3606 26854 3640
rect 26888 3606 26922 3640
rect 26956 3606 26990 3640
rect 27024 3606 27058 3640
rect 27092 3606 27126 3640
rect 27160 3606 27194 3640
rect 27228 3606 27262 3640
rect 27296 3606 27330 3640
rect 27364 3606 27398 3640
rect 27432 3606 27466 3640
rect 27500 3606 27534 3640
rect 27568 3606 27602 3640
rect 27636 3606 27670 3640
rect 27704 3606 27738 3640
rect 27772 3606 27806 3640
rect 27840 3606 27874 3640
rect 27908 3606 27942 3640
rect 27976 3606 28010 3640
rect 28044 3606 28078 3640
rect 28112 3606 28146 3640
rect 28180 3606 28214 3640
rect 28248 3606 28282 3640
rect 28316 3606 28350 3640
rect 28384 3606 28418 3640
rect 28452 3606 28486 3640
rect 28520 3606 28554 3640
rect 28588 3606 28622 3640
rect 28656 3606 28690 3640
rect 28724 3606 28758 3640
rect 28792 3606 28826 3640
rect 28860 3606 28894 3640
rect 28928 3606 28962 3640
rect 28996 3606 29030 3640
rect 29064 3606 29098 3640
rect 29132 3606 29166 3640
rect 29200 3606 29234 3640
rect 29268 3606 29302 3640
rect 29336 3606 29370 3640
rect 29404 3606 29438 3640
rect 29472 3606 29506 3640
rect 29540 3606 29574 3640
rect 29608 3606 29642 3640
rect 29676 3606 29710 3640
rect 29744 3606 29778 3640
rect 29812 3606 29846 3640
rect 29880 3606 29914 3640
rect 29948 3606 29982 3640
rect 30016 3606 30050 3640
rect 30084 3606 30118 3640
rect 30152 3606 30186 3640
rect 30220 3606 30254 3640
rect 30288 3606 30322 3640
rect 30356 3606 30390 3640
rect 30424 3606 30458 3640
rect 30492 3606 30526 3640
rect 30560 3606 30594 3640
rect 30628 3606 30662 3640
rect 30696 3606 30730 3640
rect 30764 3606 30798 3640
rect 30832 3606 30866 3640
rect 30900 3606 30934 3640
rect 30968 3606 31002 3640
rect 31036 3606 31070 3640
rect 31104 3606 31138 3640
rect 31172 3606 31206 3640
rect 31240 3606 31274 3640
rect 31308 3606 31342 3640
rect 31376 3606 31410 3640
rect 31444 3606 31478 3640
rect 31512 3606 31546 3640
rect 31580 3606 31614 3640
rect 31648 3606 31682 3640
rect 31716 3606 31750 3640
rect 31784 3606 31818 3640
rect 31852 3606 31886 3640
rect 31920 3606 31954 3640
rect 31988 3606 32022 3640
rect 32056 3606 32090 3640
rect 32124 3606 32158 3640
rect 32192 3606 32226 3640
rect 32260 3606 32294 3640
rect 32328 3606 32362 3640
rect 32396 3606 32430 3640
rect 32464 3606 32498 3640
rect 32532 3606 32566 3640
rect 32600 3606 32634 3640
rect 32668 3606 32702 3640
rect 32736 3606 32770 3640
rect 32804 3606 32838 3640
rect 32872 3606 32906 3640
rect 32940 3606 32974 3640
rect 33008 3606 33042 3640
rect 33076 3606 33110 3640
rect 33144 3606 33178 3640
rect 33212 3606 33246 3640
rect 33280 3606 33314 3640
rect 33348 3606 33382 3640
rect 33416 3606 33450 3640
rect 33484 3606 33518 3640
rect 33552 3606 33586 3640
rect 33620 3606 33654 3640
rect 33688 3606 33722 3640
rect 33756 3606 33790 3640
rect 33824 3606 33858 3640
rect 33892 3606 33926 3640
rect 33960 3606 33994 3640
rect 34028 3606 34062 3640
rect 34096 3606 34130 3640
rect 34164 3606 34198 3640
rect 34232 3606 34266 3640
rect 34300 3606 34334 3640
rect 34368 3606 34402 3640
rect 34436 3606 34470 3640
rect 34504 3606 34538 3640
rect 34572 3606 34606 3640
rect 34640 3606 34674 3640
rect 34708 3606 34742 3640
rect 34776 3606 34810 3640
rect 34844 3606 34878 3640
rect 34912 3606 34946 3640
rect 34980 3606 35014 3640
rect 35048 3606 35082 3640
rect 35116 3606 35150 3640
rect 35184 3606 35218 3640
rect 35252 3606 35286 3640
rect 35320 3606 35354 3640
rect 35388 3606 35422 3640
rect 35456 3606 35490 3640
rect 35524 3606 35558 3640
rect 35592 3606 35626 3640
rect 35660 3606 35694 3640
rect 35728 3606 35762 3640
rect 35796 3606 35830 3640
rect 35864 3606 35898 3640
rect 35932 3606 35966 3640
rect 36000 3606 36034 3640
rect 36068 3606 36102 3640
rect 36136 3606 36170 3640
rect 36204 3606 36238 3640
rect 36272 3606 36306 3640
rect 36340 3606 36374 3640
rect 36408 3606 36442 3640
rect 36476 3606 36510 3640
rect 36544 3606 36578 3640
rect 36612 3606 36646 3640
rect 36680 3606 36714 3640
rect 36748 3606 36782 3640
rect 36816 3606 36850 3640
rect 36884 3606 36918 3640
rect 36952 3606 36986 3640
rect 37020 3606 37054 3640
rect 37088 3606 37122 3640
rect 37156 3606 37190 3640
rect 37224 3606 37258 3640
rect 37292 3606 37326 3640
rect 37360 3606 37394 3640
rect 37428 3606 37462 3640
rect 37496 3606 37530 3640
rect 37564 3606 37598 3640
rect 37632 3606 37666 3640
rect 37700 3606 37734 3640
rect 37768 3606 37802 3640
rect 37836 3606 37870 3640
rect 37904 3606 37938 3640
rect 37972 3606 38006 3640
rect 38040 3606 38074 3640
rect 38108 3606 38142 3640
rect 38176 3606 38210 3640
rect 38244 3606 38278 3640
rect 38312 3606 38346 3640
rect 38380 3606 38414 3640
rect 38448 3606 38482 3640
rect 38516 3606 38550 3640
rect 38584 3606 38618 3640
rect 38652 3606 38686 3640
rect 38720 3606 38754 3640
rect 38788 3606 38822 3640
rect 38856 3606 38890 3640
rect 38924 3606 38958 3640
rect 38992 3606 39026 3640
rect 39060 3606 39094 3640
rect 39128 3606 39162 3640
rect 39196 3606 39230 3640
rect 39264 3606 39298 3640
rect 39332 3606 39366 3640
rect 39400 3606 39434 3640
rect 39468 3606 39502 3640
rect 39536 3606 39570 3640
rect 39604 3606 39638 3640
rect 39672 3606 39706 3640
rect 39740 3606 39774 3640
rect 39808 3606 39842 3640
rect 39876 3606 39910 3640
rect 39944 3606 39978 3640
rect 40012 3606 40046 3640
rect 40080 3606 40114 3640
rect 40148 3606 40182 3640
rect 40216 3606 40250 3640
rect 40284 3606 40318 3640
rect 40352 3606 40386 3640
rect 40420 3606 40454 3640
rect 40488 3606 40522 3640
rect 40556 3606 40590 3640
rect 40624 3606 40658 3640
rect 40692 3606 40726 3640
rect 40760 3606 40794 3640
rect 40828 3606 40862 3640
rect 40896 3606 40930 3640
rect 40964 3606 40998 3640
rect 41032 3606 41066 3640
rect 41100 3606 41134 3640
rect 41168 3606 41202 3640
rect 41236 3606 41270 3640
rect 41304 3606 41338 3640
rect 41372 3606 41406 3640
rect 41440 3606 41474 3640
rect 41508 3606 41542 3640
rect 41576 3606 41610 3640
rect 41644 3606 41678 3640
rect 41712 3606 41746 3640
rect 41780 3606 41814 3640
rect 41848 3606 41882 3640
rect 41916 3606 41950 3640
rect 41984 3606 42018 3640
rect 42052 3606 42086 3640
rect 42120 3606 42154 3640
rect 42188 3606 42222 3640
rect 42256 3606 42290 3640
rect 42324 3606 42358 3640
rect 42392 3606 42426 3640
rect 42460 3606 42494 3640
rect 42528 3606 42562 3640
rect 42596 3606 42630 3640
rect 42664 3606 42698 3640
rect 42732 3606 42766 3640
rect 42800 3606 42834 3640
rect 42868 3606 42902 3640
rect 42936 3606 42970 3640
rect 43004 3606 43038 3640
rect 43072 3606 43106 3640
rect 43140 3606 43174 3640
rect 43208 3606 43242 3640
rect 43276 3606 43310 3640
rect 43344 3606 43378 3640
rect 43412 3606 43446 3640
rect 43480 3606 43514 3640
rect 43548 3606 43582 3640
rect 43616 3606 43650 3640
rect 43684 3606 43718 3640
rect 43752 3606 43786 3640
rect 43820 3606 43854 3640
rect 43888 3606 43922 3640
rect 43956 3606 43990 3640
rect 44024 3606 44058 3640
rect 44092 3606 44126 3640
rect 44160 3606 44194 3640
rect 44228 3606 44262 3640
rect 44296 3606 44330 3640
rect 44364 3606 44398 3640
rect 44432 3606 44466 3640
rect 44500 3606 44534 3640
rect 44568 3606 44602 3640
rect 44636 3606 44670 3640
rect 44704 3606 44738 3640
rect 44772 3606 44806 3640
rect 44840 3606 44874 3640
rect 44908 3606 44942 3640
rect 44976 3606 45010 3640
rect 45044 3606 45078 3640
rect 45112 3606 45146 3640
rect 45180 3606 45214 3640
rect 45248 3606 45282 3640
rect 45316 3606 45350 3640
rect 45384 3606 45418 3640
rect 45452 3606 45486 3640
rect 45520 3606 45554 3640
rect 45588 3606 45622 3640
rect 45656 3606 45690 3640
rect 45724 3606 45758 3640
rect 45792 3606 45826 3640
rect 45860 3606 45894 3640
rect 45928 3606 45962 3640
rect 45996 3606 46030 3640
rect 46064 3606 46098 3640
rect 46132 3606 46166 3640
rect 46200 3606 46234 3640
rect 46268 3606 46302 3640
rect 46336 3606 46370 3640
rect 46404 3606 46438 3640
rect 46472 3606 46506 3640
rect 46540 3606 46574 3640
rect 46608 3606 46642 3640
rect 46676 3606 46710 3640
rect 46744 3606 46778 3640
rect 46812 3606 46846 3640
rect 46880 3606 46914 3640
rect 46948 3606 46982 3640
rect 47016 3606 47050 3640
rect 47084 3606 47118 3640
rect 47152 3606 47250 3640
rect -2416 3586 47250 3606
<< nsubdiffcont >>
rect -2318 116750 -2284 116784
rect -2250 116750 -2216 116784
rect -2182 116750 -2148 116784
rect -2114 116750 -2080 116784
rect -2046 116750 -2012 116784
rect -1978 116750 -1944 116784
rect -1910 116750 -1876 116784
rect -1842 116750 -1808 116784
rect -1774 116750 -1740 116784
rect -1706 116750 -1672 116784
rect -1638 116750 -1604 116784
rect -1570 116750 -1536 116784
rect -1502 116750 -1468 116784
rect -1434 116750 -1400 116784
rect -1366 116750 -1332 116784
rect -1298 116750 -1264 116784
rect -1230 116750 -1196 116784
rect -1162 116750 -1128 116784
rect -1094 116750 -1060 116784
rect -1026 116750 -992 116784
rect -958 116750 -924 116784
rect -890 116750 -856 116784
rect -822 116750 -788 116784
rect -754 116750 -720 116784
rect -686 116750 -652 116784
rect -618 116750 -584 116784
rect -550 116750 -516 116784
rect -482 116750 -448 116784
rect -414 116750 -380 116784
rect -346 116750 -312 116784
rect -278 116750 -244 116784
rect -210 116750 -176 116784
rect -142 116750 -108 116784
rect -74 116750 -40 116784
rect -6 116750 28 116784
rect 62 116750 96 116784
rect 130 116750 164 116784
rect 198 116750 232 116784
rect 266 116750 300 116784
rect 334 116750 368 116784
rect 402 116750 436 116784
rect 470 116750 504 116784
rect 538 116750 572 116784
rect 606 116750 640 116784
rect 674 116750 708 116784
rect 742 116750 776 116784
rect 810 116750 844 116784
rect 878 116750 912 116784
rect 946 116750 980 116784
rect 1014 116750 1048 116784
rect 1082 116750 1116 116784
rect 1150 116750 1184 116784
rect 1218 116750 1252 116784
rect 1286 116750 1320 116784
rect 1354 116750 1388 116784
rect 1422 116750 1456 116784
rect 1490 116750 1524 116784
rect 1558 116750 1592 116784
rect 1626 116750 1660 116784
rect 1694 116750 1728 116784
rect 1762 116750 1796 116784
rect 1830 116750 1864 116784
rect 1898 116750 1932 116784
rect 1966 116750 2000 116784
rect 2034 116750 2068 116784
rect 2102 116750 2136 116784
rect 2170 116750 2204 116784
rect 2238 116750 2272 116784
rect 2306 116750 2340 116784
rect 2374 116750 2408 116784
rect 2442 116750 2476 116784
rect 2510 116750 2544 116784
rect 2578 116750 2612 116784
rect 2646 116750 2680 116784
rect 2714 116750 2748 116784
rect 2782 116750 2816 116784
rect 2850 116750 2884 116784
rect 2918 116750 2952 116784
rect 2986 116750 3020 116784
rect 3054 116750 3088 116784
rect 3122 116750 3156 116784
rect 3190 116750 3224 116784
rect 3258 116750 3292 116784
rect 3326 116750 3360 116784
rect 3394 116750 3428 116784
rect 3462 116750 3496 116784
rect 3530 116750 3564 116784
rect 3598 116750 3632 116784
rect 3666 116750 3700 116784
rect 3734 116750 3768 116784
rect 3802 116750 3836 116784
rect 3870 116750 3904 116784
rect 3938 116750 3972 116784
rect 4006 116750 4040 116784
rect 4074 116750 4108 116784
rect 4142 116750 4176 116784
rect 4210 116750 4244 116784
rect 4278 116750 4312 116784
rect 4346 116750 4380 116784
rect 4414 116750 4448 116784
rect 4482 116750 4516 116784
rect 4550 116750 4584 116784
rect 4618 116750 4652 116784
rect 4686 116750 4720 116784
rect 4754 116750 4788 116784
rect 4822 116750 4856 116784
rect 4890 116750 4924 116784
rect 4958 116750 4992 116784
rect 5026 116750 5060 116784
rect 5094 116750 5128 116784
rect 5162 116750 5196 116784
rect 5230 116750 5264 116784
rect 5298 116750 5332 116784
rect 5366 116750 5400 116784
rect 5434 116750 5468 116784
rect 5502 116750 5536 116784
rect 5570 116750 5604 116784
rect 5638 116750 5672 116784
rect 5706 116750 5740 116784
rect 5774 116750 5808 116784
rect 5842 116750 5876 116784
rect 5910 116750 5944 116784
rect 5978 116750 6012 116784
rect 6046 116750 6080 116784
rect 6114 116750 6148 116784
rect 6182 116750 6216 116784
rect 6250 116750 6284 116784
rect 6318 116750 6352 116784
rect 6386 116750 6420 116784
rect 6454 116750 6488 116784
rect 6522 116750 6556 116784
rect 6590 116750 6624 116784
rect 6658 116750 6692 116784
rect 6726 116750 6760 116784
rect 6794 116750 6828 116784
rect 6862 116750 6896 116784
rect 6930 116750 6964 116784
rect 6998 116750 7032 116784
rect 7066 116750 7100 116784
rect 7134 116750 7168 116784
rect 7202 116750 7236 116784
rect 7270 116750 7304 116784
rect 7338 116750 7372 116784
rect 7406 116750 7440 116784
rect 7474 116750 7508 116784
rect 7542 116750 7576 116784
rect 7610 116750 7644 116784
rect 7678 116750 7712 116784
rect 7746 116750 7780 116784
rect 7814 116750 7848 116784
rect 7882 116750 7916 116784
rect 7950 116750 7984 116784
rect 8018 116750 8052 116784
rect 8086 116750 8120 116784
rect 8154 116750 8188 116784
rect 8222 116750 8256 116784
rect 8290 116750 8324 116784
rect 8358 116750 8392 116784
rect 8426 116750 8460 116784
rect 8494 116750 8528 116784
rect 8562 116750 8596 116784
rect 8630 116750 8664 116784
rect 8698 116750 8732 116784
rect 8766 116750 8800 116784
rect 8834 116750 8868 116784
rect 8902 116750 8936 116784
rect 8970 116750 9004 116784
rect 9038 116750 9072 116784
rect 9106 116750 9140 116784
rect 9174 116750 9208 116784
rect 9242 116750 9276 116784
rect 9310 116750 9344 116784
rect 9378 116750 9412 116784
rect 9446 116750 9480 116784
rect 9514 116750 9548 116784
rect 9582 116750 9616 116784
rect 9650 116750 9684 116784
rect 9718 116750 9752 116784
rect 9786 116750 9820 116784
rect 9854 116750 9888 116784
rect 9922 116750 9956 116784
rect 9990 116750 10024 116784
rect 10058 116750 10092 116784
rect 10126 116750 10160 116784
rect 10194 116750 10228 116784
rect 10262 116750 10296 116784
rect 10330 116750 10364 116784
rect 10398 116750 10432 116784
rect 10466 116750 10500 116784
rect 10534 116750 10568 116784
rect 10602 116750 10636 116784
rect 10670 116750 10704 116784
rect 10738 116750 10772 116784
rect 10806 116750 10840 116784
rect 10874 116750 10908 116784
rect 10942 116750 10976 116784
rect 11010 116750 11044 116784
rect 11078 116750 11112 116784
rect 11146 116750 11180 116784
rect 11214 116750 11248 116784
rect 11282 116750 11316 116784
rect 11350 116750 11384 116784
rect 11418 116750 11452 116784
rect 11486 116750 11520 116784
rect 11554 116750 11588 116784
rect 11622 116750 11656 116784
rect 11690 116750 11724 116784
rect 11758 116750 11792 116784
rect 11826 116750 11860 116784
rect 11894 116750 11928 116784
rect 11962 116750 11996 116784
rect 12030 116750 12064 116784
rect 12098 116750 12132 116784
rect 12166 116750 12200 116784
rect 12234 116750 12268 116784
rect 12302 116750 12336 116784
rect 12370 116750 12404 116784
rect 12438 116750 12472 116784
rect 12506 116750 12540 116784
rect 12574 116750 12608 116784
rect 12642 116750 12676 116784
rect 12710 116750 12744 116784
rect 12778 116750 12812 116784
rect 12846 116750 12880 116784
rect 12914 116750 12948 116784
rect 12982 116750 13016 116784
rect 13050 116750 13084 116784
rect 13118 116750 13152 116784
rect 13186 116750 13220 116784
rect 13254 116750 13288 116784
rect 13322 116750 13356 116784
rect 13390 116750 13424 116784
rect 13458 116750 13492 116784
rect 13526 116750 13560 116784
rect 13594 116750 13628 116784
rect 13662 116750 13696 116784
rect 13730 116750 13764 116784
rect 13798 116750 13832 116784
rect 13866 116750 13900 116784
rect 13934 116750 13968 116784
rect 14002 116750 14036 116784
rect 14070 116750 14104 116784
rect 14138 116750 14172 116784
rect 14206 116750 14240 116784
rect 14274 116750 14308 116784
rect 14342 116750 14376 116784
rect 14410 116750 14444 116784
rect 14478 116750 14512 116784
rect 14546 116750 14580 116784
rect 14614 116750 14648 116784
rect 14682 116750 14716 116784
rect 14750 116750 14784 116784
rect 14818 116750 14852 116784
rect 14886 116750 14920 116784
rect 14954 116750 14988 116784
rect 15022 116750 15056 116784
rect 15090 116750 15124 116784
rect 15158 116750 15192 116784
rect 15226 116750 15260 116784
rect 15294 116750 15328 116784
rect 15362 116750 15396 116784
rect 15430 116750 15464 116784
rect 15498 116750 15532 116784
rect 15566 116750 15600 116784
rect 15634 116750 15668 116784
rect 15702 116750 15736 116784
rect 15770 116750 15804 116784
rect 15838 116750 15872 116784
rect 15906 116750 15940 116784
rect 15974 116750 16008 116784
rect 16042 116750 16076 116784
rect 16110 116750 16144 116784
rect 16178 116750 16212 116784
rect 16246 116750 16280 116784
rect 16314 116750 16348 116784
rect 16382 116750 16416 116784
rect 16450 116750 16484 116784
rect 16518 116750 16552 116784
rect 16586 116750 16620 116784
rect 16654 116750 16688 116784
rect 16722 116750 16756 116784
rect 16790 116750 16824 116784
rect 16858 116750 16892 116784
rect 16926 116750 16960 116784
rect 16994 116750 17028 116784
rect 17062 116750 17096 116784
rect 17130 116750 17164 116784
rect 17198 116750 17232 116784
rect 17266 116750 17300 116784
rect 17334 116750 17368 116784
rect 17402 116750 17436 116784
rect 17470 116750 17504 116784
rect 17538 116750 17572 116784
rect 17606 116750 17640 116784
rect 17674 116750 17708 116784
rect 17742 116750 17776 116784
rect 17810 116750 17844 116784
rect 17878 116750 17912 116784
rect 17946 116750 17980 116784
rect 18014 116750 18048 116784
rect 18082 116750 18116 116784
rect 18150 116750 18184 116784
rect 18218 116750 18252 116784
rect 18286 116750 18320 116784
rect 18354 116750 18388 116784
rect 18422 116750 18456 116784
rect 18490 116750 18524 116784
rect 18558 116750 18592 116784
rect 18626 116750 18660 116784
rect 18694 116750 18728 116784
rect 18762 116750 18796 116784
rect 18830 116750 18864 116784
rect 18898 116750 18932 116784
rect 18966 116750 19000 116784
rect 19034 116750 19068 116784
rect 19102 116750 19136 116784
rect 19170 116750 19204 116784
rect 19238 116750 19272 116784
rect 19306 116750 19340 116784
rect 19374 116750 19408 116784
rect 19442 116750 19476 116784
rect 19510 116750 19544 116784
rect 19578 116750 19612 116784
rect 19646 116750 19680 116784
rect 19714 116750 19748 116784
rect 19782 116750 19816 116784
rect 19850 116750 19884 116784
rect 19918 116750 19952 116784
rect 19986 116750 20020 116784
rect 20054 116750 20088 116784
rect 20122 116750 20156 116784
rect 20190 116750 20224 116784
rect 20258 116750 20292 116784
rect 20326 116750 20360 116784
rect 20394 116750 20428 116784
rect 20462 116750 20496 116784
rect 20530 116750 20564 116784
rect 20598 116750 20632 116784
rect 20666 116750 20700 116784
rect 20734 116750 20768 116784
rect 20802 116750 20836 116784
rect 20870 116750 20904 116784
rect 20938 116750 20972 116784
rect 21006 116750 21040 116784
rect 21074 116750 21108 116784
rect 21142 116750 21176 116784
rect 21210 116750 21244 116784
rect 21278 116750 21312 116784
rect 21346 116750 21380 116784
rect 21414 116750 21448 116784
rect 21482 116750 21516 116784
rect 21550 116750 21584 116784
rect 21618 116750 21652 116784
rect 21686 116750 21720 116784
rect 21754 116750 21788 116784
rect 21822 116750 21856 116784
rect 21890 116750 21924 116784
rect 21958 116750 21992 116784
rect 22026 116750 22060 116784
rect 22094 116750 22128 116784
rect 22162 116750 22196 116784
rect 22230 116750 22264 116784
rect 22298 116750 22332 116784
rect 22366 116750 22400 116784
rect 22434 116750 22468 116784
rect 22502 116750 22536 116784
rect 22570 116750 22604 116784
rect 22638 116750 22672 116784
rect 22706 116750 22740 116784
rect 22774 116750 22808 116784
rect 22842 116750 22876 116784
rect 22910 116750 22944 116784
rect 22978 116750 23012 116784
rect 23046 116750 23080 116784
rect 23114 116750 23148 116784
rect 23182 116750 23216 116784
rect 23250 116750 23284 116784
rect 23318 116750 23352 116784
rect 23386 116750 23420 116784
rect 23454 116750 23488 116784
rect 23522 116750 23556 116784
rect 23590 116750 23624 116784
rect 23658 116750 23692 116784
rect 23726 116750 23760 116784
rect 23794 116750 23828 116784
rect 23862 116750 23896 116784
rect 23930 116750 23964 116784
rect 23998 116750 24032 116784
rect 24066 116750 24100 116784
rect 24134 116750 24168 116784
rect 24202 116750 24236 116784
rect 24270 116750 24304 116784
rect 24338 116750 24372 116784
rect 24406 116750 24440 116784
rect 24474 116750 24508 116784
rect 24542 116750 24576 116784
rect 24610 116750 24644 116784
rect 24678 116750 24712 116784
rect 24746 116750 24780 116784
rect 24814 116750 24848 116784
rect 24882 116750 24916 116784
rect 24950 116750 24984 116784
rect 25018 116750 25052 116784
rect 25086 116750 25120 116784
rect 25154 116750 25188 116784
rect 25222 116750 25256 116784
rect 25290 116750 25324 116784
rect 25358 116750 25392 116784
rect 25426 116750 25460 116784
rect 25494 116750 25528 116784
rect 25562 116750 25596 116784
rect 25630 116750 25664 116784
rect 25698 116750 25732 116784
rect 25766 116750 25800 116784
rect 25834 116750 25868 116784
rect 25902 116750 25936 116784
rect 25970 116750 26004 116784
rect 26038 116750 26072 116784
rect 26106 116750 26140 116784
rect 26174 116750 26208 116784
rect 26242 116750 26276 116784
rect 26310 116750 26344 116784
rect 26378 116750 26412 116784
rect 26446 116750 26480 116784
rect 26514 116750 26548 116784
rect 26582 116750 26616 116784
rect 26650 116750 26684 116784
rect 26718 116750 26752 116784
rect 26786 116750 26820 116784
rect 26854 116750 26888 116784
rect 26922 116750 26956 116784
rect 26990 116750 27024 116784
rect 27058 116750 27092 116784
rect 27126 116750 27160 116784
rect 27194 116750 27228 116784
rect 27262 116750 27296 116784
rect 27330 116750 27364 116784
rect 27398 116750 27432 116784
rect 27466 116750 27500 116784
rect 27534 116750 27568 116784
rect 27602 116750 27636 116784
rect 27670 116750 27704 116784
rect 27738 116750 27772 116784
rect 27806 116750 27840 116784
rect 27874 116750 27908 116784
rect 27942 116750 27976 116784
rect 28010 116750 28044 116784
rect 28078 116750 28112 116784
rect 28146 116750 28180 116784
rect 28214 116750 28248 116784
rect 28282 116750 28316 116784
rect 28350 116750 28384 116784
rect 28418 116750 28452 116784
rect 28486 116750 28520 116784
rect 28554 116750 28588 116784
rect 28622 116750 28656 116784
rect 28690 116750 28724 116784
rect 28758 116750 28792 116784
rect 28826 116750 28860 116784
rect 28894 116750 28928 116784
rect 28962 116750 28996 116784
rect 29030 116750 29064 116784
rect 29098 116750 29132 116784
rect 29166 116750 29200 116784
rect 29234 116750 29268 116784
rect 29302 116750 29336 116784
rect 29370 116750 29404 116784
rect 29438 116750 29472 116784
rect 29506 116750 29540 116784
rect 29574 116750 29608 116784
rect 29642 116750 29676 116784
rect 29710 116750 29744 116784
rect 29778 116750 29812 116784
rect 29846 116750 29880 116784
rect 29914 116750 29948 116784
rect 29982 116750 30016 116784
rect 30050 116750 30084 116784
rect 30118 116750 30152 116784
rect 30186 116750 30220 116784
rect 30254 116750 30288 116784
rect 30322 116750 30356 116784
rect 30390 116750 30424 116784
rect 30458 116750 30492 116784
rect 30526 116750 30560 116784
rect 30594 116750 30628 116784
rect 30662 116750 30696 116784
rect 30730 116750 30764 116784
rect 30798 116750 30832 116784
rect 30866 116750 30900 116784
rect 30934 116750 30968 116784
rect 31002 116750 31036 116784
rect 31070 116750 31104 116784
rect 31138 116750 31172 116784
rect 31206 116750 31240 116784
rect 31274 116750 31308 116784
rect 31342 116750 31376 116784
rect 31410 116750 31444 116784
rect 31478 116750 31512 116784
rect 31546 116750 31580 116784
rect 31614 116750 31648 116784
rect 31682 116750 31716 116784
rect 31750 116750 31784 116784
rect 31818 116750 31852 116784
rect 31886 116750 31920 116784
rect 31954 116750 31988 116784
rect 32022 116750 32056 116784
rect 32090 116750 32124 116784
rect 32158 116750 32192 116784
rect 32226 116750 32260 116784
rect 32294 116750 32328 116784
rect 32362 116750 32396 116784
rect 32430 116750 32464 116784
rect 32498 116750 32532 116784
rect 32566 116750 32600 116784
rect 32634 116750 32668 116784
rect 32702 116750 32736 116784
rect 32770 116750 32804 116784
rect 32838 116750 32872 116784
rect 32906 116750 32940 116784
rect 32974 116750 33008 116784
rect 33042 116750 33076 116784
rect 33110 116750 33144 116784
rect 33178 116750 33212 116784
rect 33246 116750 33280 116784
rect 33314 116750 33348 116784
rect 33382 116750 33416 116784
rect 33450 116750 33484 116784
rect 33518 116750 33552 116784
rect 33586 116750 33620 116784
rect 33654 116750 33688 116784
rect 33722 116750 33756 116784
rect 33790 116750 33824 116784
rect 33858 116750 33892 116784
rect 33926 116750 33960 116784
rect 33994 116750 34028 116784
rect 34062 116750 34096 116784
rect 34130 116750 34164 116784
rect 34198 116750 34232 116784
rect 34266 116750 34300 116784
rect 34334 116750 34368 116784
rect 34402 116750 34436 116784
rect 34470 116750 34504 116784
rect 34538 116750 34572 116784
rect 34606 116750 34640 116784
rect 34674 116750 34708 116784
rect 34742 116750 34776 116784
rect 34810 116750 34844 116784
rect 34878 116750 34912 116784
rect 34946 116750 34980 116784
rect 35014 116750 35048 116784
rect 35082 116750 35116 116784
rect 35150 116750 35184 116784
rect 35218 116750 35252 116784
rect 35286 116750 35320 116784
rect 35354 116750 35388 116784
rect 35422 116750 35456 116784
rect 35490 116750 35524 116784
rect 35558 116750 35592 116784
rect 35626 116750 35660 116784
rect 35694 116750 35728 116784
rect 35762 116750 35796 116784
rect 35830 116750 35864 116784
rect 35898 116750 35932 116784
rect 35966 116750 36000 116784
rect 36034 116750 36068 116784
rect 36102 116750 36136 116784
rect 36170 116750 36204 116784
rect 36238 116750 36272 116784
rect 36306 116750 36340 116784
rect 36374 116750 36408 116784
rect 36442 116750 36476 116784
rect 36510 116750 36544 116784
rect 36578 116750 36612 116784
rect 36646 116750 36680 116784
rect 36714 116750 36748 116784
rect 36782 116750 36816 116784
rect 36850 116750 36884 116784
rect 36918 116750 36952 116784
rect 36986 116750 37020 116784
rect 37054 116750 37088 116784
rect 37122 116750 37156 116784
rect 37190 116750 37224 116784
rect 37258 116750 37292 116784
rect 37326 116750 37360 116784
rect 37394 116750 37428 116784
rect 37462 116750 37496 116784
rect 37530 116750 37564 116784
rect 37598 116750 37632 116784
rect 37666 116750 37700 116784
rect 37734 116750 37768 116784
rect 37802 116750 37836 116784
rect 37870 116750 37904 116784
rect 37938 116750 37972 116784
rect 38006 116750 38040 116784
rect 38074 116750 38108 116784
rect 38142 116750 38176 116784
rect 38210 116750 38244 116784
rect 38278 116750 38312 116784
rect 38346 116750 38380 116784
rect 38414 116750 38448 116784
rect 38482 116750 38516 116784
rect 38550 116750 38584 116784
rect 38618 116750 38652 116784
rect 38686 116750 38720 116784
rect 38754 116750 38788 116784
rect 38822 116750 38856 116784
rect 38890 116750 38924 116784
rect 38958 116750 38992 116784
rect 39026 116750 39060 116784
rect 39094 116750 39128 116784
rect 39162 116750 39196 116784
rect 39230 116750 39264 116784
rect 39298 116750 39332 116784
rect 39366 116750 39400 116784
rect 39434 116750 39468 116784
rect 39502 116750 39536 116784
rect 39570 116750 39604 116784
rect 39638 116750 39672 116784
rect 39706 116750 39740 116784
rect 39774 116750 39808 116784
rect 39842 116750 39876 116784
rect 39910 116750 39944 116784
rect 39978 116750 40012 116784
rect 40046 116750 40080 116784
rect 40114 116750 40148 116784
rect 40182 116750 40216 116784
rect 40250 116750 40284 116784
rect 40318 116750 40352 116784
rect 40386 116750 40420 116784
rect 40454 116750 40488 116784
rect 40522 116750 40556 116784
rect 40590 116750 40624 116784
rect 40658 116750 40692 116784
rect 40726 116750 40760 116784
rect 40794 116750 40828 116784
rect 40862 116750 40896 116784
rect 40930 116750 40964 116784
rect 40998 116750 41032 116784
rect 41066 116750 41100 116784
rect 41134 116750 41168 116784
rect 41202 116750 41236 116784
rect 41270 116750 41304 116784
rect 41338 116750 41372 116784
rect 41406 116750 41440 116784
rect 41474 116750 41508 116784
rect 41542 116750 41576 116784
rect 41610 116750 41644 116784
rect 41678 116750 41712 116784
rect 41746 116750 41780 116784
rect 41814 116750 41848 116784
rect 41882 116750 41916 116784
rect 41950 116750 41984 116784
rect 42018 116750 42052 116784
rect 42086 116750 42120 116784
rect 42154 116750 42188 116784
rect 42222 116750 42256 116784
rect 42290 116750 42324 116784
rect 42358 116750 42392 116784
rect 42426 116750 42460 116784
rect 42494 116750 42528 116784
rect 42562 116750 42596 116784
rect 42630 116750 42664 116784
rect 42698 116750 42732 116784
rect 42766 116750 42800 116784
rect 42834 116750 42868 116784
rect 42902 116750 42936 116784
rect 42970 116750 43004 116784
rect 43038 116750 43072 116784
rect 43106 116750 43140 116784
rect 43174 116750 43208 116784
rect 43242 116750 43276 116784
rect 43310 116750 43344 116784
rect 43378 116750 43412 116784
rect 43446 116750 43480 116784
rect 43514 116750 43548 116784
rect 43582 116750 43616 116784
rect 43650 116750 43684 116784
rect 43718 116750 43752 116784
rect 43786 116750 43820 116784
rect 43854 116750 43888 116784
rect 43922 116750 43956 116784
rect 43990 116750 44024 116784
rect 44058 116750 44092 116784
rect 44126 116750 44160 116784
rect 44194 116750 44228 116784
rect 44262 116750 44296 116784
rect 44330 116750 44364 116784
rect 44398 116750 44432 116784
rect 44466 116750 44500 116784
rect 44534 116750 44568 116784
rect 44602 116750 44636 116784
rect 44670 116750 44704 116784
rect 44738 116750 44772 116784
rect 44806 116750 44840 116784
rect 44874 116750 44908 116784
rect 44942 116750 44976 116784
rect 45010 116750 45044 116784
rect 45078 116750 45112 116784
rect 45146 116750 45180 116784
rect 45214 116750 45248 116784
rect 45282 116750 45316 116784
rect 45350 116750 45384 116784
rect 45418 116750 45452 116784
rect 45486 116750 45520 116784
rect 45554 116750 45588 116784
rect 45622 116750 45656 116784
rect 45690 116750 45724 116784
rect 45758 116750 45792 116784
rect 45826 116750 45860 116784
rect 45894 116750 45928 116784
rect 45962 116750 45996 116784
rect 46030 116750 46064 116784
rect 46098 116750 46132 116784
rect 46166 116750 46200 116784
rect 46234 116750 46268 116784
rect 46302 116750 46336 116784
rect 46370 116750 46404 116784
rect 46438 116750 46472 116784
rect 46506 116750 46540 116784
rect 46574 116750 46608 116784
rect 46642 116750 46676 116784
rect 46710 116750 46744 116784
rect 46778 116750 46812 116784
rect 46846 116750 46880 116784
rect 46914 116750 46948 116784
rect 46982 116750 47016 116784
rect 47050 116750 47084 116784
rect 47118 116750 47152 116784
rect -2396 116663 -2362 116697
rect -2396 116595 -2362 116629
rect -2396 116527 -2362 116561
rect -2396 116459 -2362 116493
rect -2396 116391 -2362 116425
rect -2396 116323 -2362 116357
rect -2396 116255 -2362 116289
rect -2396 116187 -2362 116221
rect -2396 116119 -2362 116153
rect -2396 116051 -2362 116085
rect -2396 115983 -2362 116017
rect -2396 115915 -2362 115949
rect -2396 115847 -2362 115881
rect -2396 115779 -2362 115813
rect -2396 115711 -2362 115745
rect -2396 115643 -2362 115677
rect -2396 115575 -2362 115609
rect -2396 115507 -2362 115541
rect -2396 115439 -2362 115473
rect -2396 115371 -2362 115405
rect -2396 115303 -2362 115337
rect -2396 115235 -2362 115269
rect -2396 115167 -2362 115201
rect -2396 115099 -2362 115133
rect -2396 115031 -2362 115065
rect -2396 114963 -2362 114997
rect -2396 114895 -2362 114929
rect -2396 114827 -2362 114861
rect -2396 114759 -2362 114793
rect -2396 114691 -2362 114725
rect -2396 114623 -2362 114657
rect -2396 114555 -2362 114589
rect -2396 114487 -2362 114521
rect -2396 114419 -2362 114453
rect -2396 114351 -2362 114385
rect -2396 114283 -2362 114317
rect -2396 114215 -2362 114249
rect -2396 114147 -2362 114181
rect -2396 114079 -2362 114113
rect -2396 114011 -2362 114045
rect -2396 113943 -2362 113977
rect -2396 113875 -2362 113909
rect -2396 113807 -2362 113841
rect -2396 113739 -2362 113773
rect -2396 113671 -2362 113705
rect -2396 113603 -2362 113637
rect -2396 113535 -2362 113569
rect -2396 113467 -2362 113501
rect -2396 113399 -2362 113433
rect -2396 113331 -2362 113365
rect -2396 113263 -2362 113297
rect -2396 113195 -2362 113229
rect -2396 113127 -2362 113161
rect -2396 113059 -2362 113093
rect -2396 112991 -2362 113025
rect -2396 112923 -2362 112957
rect -2396 112855 -2362 112889
rect -2396 112787 -2362 112821
rect -2396 112719 -2362 112753
rect -2396 112651 -2362 112685
rect -2396 112583 -2362 112617
rect -2396 112515 -2362 112549
rect -2396 112447 -2362 112481
rect -2396 112379 -2362 112413
rect -2396 112311 -2362 112345
rect -2396 112243 -2362 112277
rect -2396 112175 -2362 112209
rect -2396 112107 -2362 112141
rect -2396 112039 -2362 112073
rect -2396 111971 -2362 112005
rect -2396 111903 -2362 111937
rect -2396 111835 -2362 111869
rect -2396 111767 -2362 111801
rect -2396 111699 -2362 111733
rect -2396 111631 -2362 111665
rect -2396 111563 -2362 111597
rect -2396 111495 -2362 111529
rect -2396 111427 -2362 111461
rect -2396 111359 -2362 111393
rect -2396 111291 -2362 111325
rect -2396 111223 -2362 111257
rect -2396 111155 -2362 111189
rect -2396 111087 -2362 111121
rect -2396 111019 -2362 111053
rect -2396 110951 -2362 110985
rect -2396 110883 -2362 110917
rect -2396 110815 -2362 110849
rect -2396 110747 -2362 110781
rect -2396 110679 -2362 110713
rect -2396 110611 -2362 110645
rect -2396 110543 -2362 110577
rect -2396 110475 -2362 110509
rect -2396 110407 -2362 110441
rect -2396 110339 -2362 110373
rect -2396 110271 -2362 110305
rect -2396 110203 -2362 110237
rect -2396 110135 -2362 110169
rect -2396 110067 -2362 110101
rect -2396 109999 -2362 110033
rect -2396 109931 -2362 109965
rect -2396 109863 -2362 109897
rect -2396 109795 -2362 109829
rect -2396 109727 -2362 109761
rect -2396 109659 -2362 109693
rect -2396 109591 -2362 109625
rect -2396 109523 -2362 109557
rect -2396 109455 -2362 109489
rect -2396 109387 -2362 109421
rect -2396 109319 -2362 109353
rect -2396 109251 -2362 109285
rect -2396 109183 -2362 109217
rect -2396 109115 -2362 109149
rect -2396 109047 -2362 109081
rect -2396 108979 -2362 109013
rect -2396 108911 -2362 108945
rect -2396 108843 -2362 108877
rect -2396 108775 -2362 108809
rect -2396 108707 -2362 108741
rect -2396 108639 -2362 108673
rect -2396 108571 -2362 108605
rect -2396 108503 -2362 108537
rect -2396 108435 -2362 108469
rect -2396 108367 -2362 108401
rect -2396 108299 -2362 108333
rect -2396 108231 -2362 108265
rect -2396 108163 -2362 108197
rect -2396 108095 -2362 108129
rect -2396 108027 -2362 108061
rect -2396 107959 -2362 107993
rect -2396 107891 -2362 107925
rect -2396 107823 -2362 107857
rect -2396 107755 -2362 107789
rect -2396 107687 -2362 107721
rect -2396 107619 -2362 107653
rect -2396 107551 -2362 107585
rect -2396 107483 -2362 107517
rect -2396 107415 -2362 107449
rect -2396 107347 -2362 107381
rect -2396 107279 -2362 107313
rect -2396 107211 -2362 107245
rect -2396 107143 -2362 107177
rect -2396 107075 -2362 107109
rect -2396 107007 -2362 107041
rect -2396 106939 -2362 106973
rect -2396 106871 -2362 106905
rect -2396 106803 -2362 106837
rect -2396 106735 -2362 106769
rect -2396 106667 -2362 106701
rect -2396 106599 -2362 106633
rect -2396 106531 -2362 106565
rect -2396 106463 -2362 106497
rect -2396 106395 -2362 106429
rect -2396 106327 -2362 106361
rect -2396 106259 -2362 106293
rect -2396 106191 -2362 106225
rect -2396 106123 -2362 106157
rect -2396 106055 -2362 106089
rect -2396 105987 -2362 106021
rect -2396 105919 -2362 105953
rect -2396 105851 -2362 105885
rect -2396 105783 -2362 105817
rect -2396 105715 -2362 105749
rect -2396 105647 -2362 105681
rect -2396 105579 -2362 105613
rect -2396 105511 -2362 105545
rect -2396 105443 -2362 105477
rect -2396 105375 -2362 105409
rect -2396 105307 -2362 105341
rect -2396 105239 -2362 105273
rect -2396 105171 -2362 105205
rect -2396 105103 -2362 105137
rect -2396 105035 -2362 105069
rect -2396 104967 -2362 105001
rect -2396 104899 -2362 104933
rect -2396 104831 -2362 104865
rect -2396 104763 -2362 104797
rect -2396 104695 -2362 104729
rect -2396 104627 -2362 104661
rect -2396 104559 -2362 104593
rect -2396 104491 -2362 104525
rect -2396 104423 -2362 104457
rect -2396 104355 -2362 104389
rect -2396 104287 -2362 104321
rect -2396 104219 -2362 104253
rect -2396 104151 -2362 104185
rect -2396 104083 -2362 104117
rect -2396 104015 -2362 104049
rect -2396 103947 -2362 103981
rect -2396 103879 -2362 103913
rect -2396 103811 -2362 103845
rect -2396 103743 -2362 103777
rect -2396 103675 -2362 103709
rect -2396 103607 -2362 103641
rect -2396 103539 -2362 103573
rect -2396 103471 -2362 103505
rect -2396 103403 -2362 103437
rect -2396 103335 -2362 103369
rect -2396 103267 -2362 103301
rect -2396 103199 -2362 103233
rect -2396 103131 -2362 103165
rect -2396 103063 -2362 103097
rect -2396 102995 -2362 103029
rect -2396 102927 -2362 102961
rect -2396 102859 -2362 102893
rect -2396 102791 -2362 102825
rect -2396 102723 -2362 102757
rect -2396 102655 -2362 102689
rect -2396 102587 -2362 102621
rect -2396 102519 -2362 102553
rect -2396 102451 -2362 102485
rect -2396 102383 -2362 102417
rect -2396 102315 -2362 102349
rect -2396 102247 -2362 102281
rect -2396 102179 -2362 102213
rect -2396 102111 -2362 102145
rect -2396 102043 -2362 102077
rect -2396 101975 -2362 102009
rect -2396 101907 -2362 101941
rect -2396 101839 -2362 101873
rect -2396 101771 -2362 101805
rect -2396 101703 -2362 101737
rect -2396 101635 -2362 101669
rect -2396 101567 -2362 101601
rect -2396 101499 -2362 101533
rect -2396 101431 -2362 101465
rect -2396 101363 -2362 101397
rect -2396 101295 -2362 101329
rect -2396 101227 -2362 101261
rect -2396 101159 -2362 101193
rect -2396 101091 -2362 101125
rect -2396 101023 -2362 101057
rect -2396 100955 -2362 100989
rect 47196 116663 47230 116697
rect 47196 116595 47230 116629
rect 47196 116527 47230 116561
rect 47196 116459 47230 116493
rect 47196 116391 47230 116425
rect 47196 116323 47230 116357
rect 47196 116255 47230 116289
rect 47196 116187 47230 116221
rect 47196 116119 47230 116153
rect 47196 116051 47230 116085
rect 47196 115983 47230 116017
rect 47196 115915 47230 115949
rect 47196 115847 47230 115881
rect 47196 115779 47230 115813
rect 47196 115711 47230 115745
rect 47196 115643 47230 115677
rect 47196 115575 47230 115609
rect 47196 115507 47230 115541
rect 47196 115439 47230 115473
rect 47196 115371 47230 115405
rect 47196 115303 47230 115337
rect 47196 115235 47230 115269
rect 47196 115167 47230 115201
rect 47196 115099 47230 115133
rect 47196 115031 47230 115065
rect 47196 114963 47230 114997
rect 47196 114895 47230 114929
rect 47196 114827 47230 114861
rect 47196 114759 47230 114793
rect 47196 114691 47230 114725
rect 47196 114623 47230 114657
rect 47196 114555 47230 114589
rect 47196 114487 47230 114521
rect 47196 114419 47230 114453
rect 47196 114351 47230 114385
rect 47196 114283 47230 114317
rect 47196 114215 47230 114249
rect 47196 114147 47230 114181
rect 47196 114079 47230 114113
rect 47196 114011 47230 114045
rect 47196 113943 47230 113977
rect 47196 113875 47230 113909
rect 47196 113807 47230 113841
rect 47196 113739 47230 113773
rect 47196 113671 47230 113705
rect 47196 113603 47230 113637
rect 47196 113535 47230 113569
rect 47196 113467 47230 113501
rect 47196 113399 47230 113433
rect 47196 113331 47230 113365
rect 47196 113263 47230 113297
rect 47196 113195 47230 113229
rect 47196 113127 47230 113161
rect 47196 113059 47230 113093
rect 47196 112991 47230 113025
rect 47196 112923 47230 112957
rect 47196 112855 47230 112889
rect 47196 112787 47230 112821
rect 47196 112719 47230 112753
rect 47196 112651 47230 112685
rect 47196 112583 47230 112617
rect 47196 112515 47230 112549
rect 47196 112447 47230 112481
rect 47196 112379 47230 112413
rect 47196 112311 47230 112345
rect 47196 112243 47230 112277
rect 47196 112175 47230 112209
rect 47196 112107 47230 112141
rect 47196 112039 47230 112073
rect 47196 111971 47230 112005
rect 47196 111903 47230 111937
rect 47196 111835 47230 111869
rect 47196 111767 47230 111801
rect 47196 111699 47230 111733
rect 47196 111631 47230 111665
rect 47196 111563 47230 111597
rect 47196 111495 47230 111529
rect 47196 111427 47230 111461
rect 47196 111359 47230 111393
rect 47196 111291 47230 111325
rect 47196 111223 47230 111257
rect 47196 111155 47230 111189
rect 47196 111087 47230 111121
rect 47196 111019 47230 111053
rect 47196 110951 47230 110985
rect 47196 110883 47230 110917
rect 47196 110815 47230 110849
rect 47196 110747 47230 110781
rect 47196 110679 47230 110713
rect 47196 110611 47230 110645
rect 47196 110543 47230 110577
rect 47196 110475 47230 110509
rect 47196 110407 47230 110441
rect 47196 110339 47230 110373
rect 47196 110271 47230 110305
rect 47196 110203 47230 110237
rect 47196 110135 47230 110169
rect 47196 110067 47230 110101
rect 47196 109999 47230 110033
rect 47196 109931 47230 109965
rect 47196 109863 47230 109897
rect 47196 109795 47230 109829
rect 47196 109727 47230 109761
rect 47196 109659 47230 109693
rect 47196 109591 47230 109625
rect 47196 109523 47230 109557
rect 47196 109455 47230 109489
rect 47196 109387 47230 109421
rect 47196 109319 47230 109353
rect 47196 109251 47230 109285
rect 47196 109183 47230 109217
rect 47196 109115 47230 109149
rect 47196 109047 47230 109081
rect 47196 108979 47230 109013
rect 47196 108911 47230 108945
rect 47196 108843 47230 108877
rect 47196 108775 47230 108809
rect 47196 108707 47230 108741
rect 47196 108639 47230 108673
rect 47196 108571 47230 108605
rect 47196 108503 47230 108537
rect 47196 108435 47230 108469
rect 47196 108367 47230 108401
rect 47196 108299 47230 108333
rect 47196 108231 47230 108265
rect 47196 108163 47230 108197
rect 47196 108095 47230 108129
rect 47196 108027 47230 108061
rect 47196 107959 47230 107993
rect 47196 107891 47230 107925
rect 47196 107823 47230 107857
rect 47196 107755 47230 107789
rect 47196 107687 47230 107721
rect 47196 107619 47230 107653
rect 47196 107551 47230 107585
rect 47196 107483 47230 107517
rect 47196 107415 47230 107449
rect 47196 107347 47230 107381
rect 47196 107279 47230 107313
rect 47196 107211 47230 107245
rect 47196 107143 47230 107177
rect 47196 107075 47230 107109
rect 47196 107007 47230 107041
rect 47196 106939 47230 106973
rect 47196 106871 47230 106905
rect 47196 106803 47230 106837
rect 47196 106735 47230 106769
rect 47196 106667 47230 106701
rect 47196 106599 47230 106633
rect 47196 106531 47230 106565
rect 47196 106463 47230 106497
rect 47196 106395 47230 106429
rect 47196 106327 47230 106361
rect 47196 106259 47230 106293
rect 47196 106191 47230 106225
rect 47196 106123 47230 106157
rect 47196 106055 47230 106089
rect 47196 105987 47230 106021
rect 47196 105919 47230 105953
rect 47196 105851 47230 105885
rect 47196 105783 47230 105817
rect 47196 105715 47230 105749
rect 47196 105647 47230 105681
rect 47196 105579 47230 105613
rect 47196 105511 47230 105545
rect 47196 105443 47230 105477
rect 47196 105375 47230 105409
rect 47196 105307 47230 105341
rect 47196 105239 47230 105273
rect 47196 105171 47230 105205
rect 47196 105103 47230 105137
rect 47196 105035 47230 105069
rect 47196 104967 47230 105001
rect 47196 104899 47230 104933
rect 47196 104831 47230 104865
rect 47196 104763 47230 104797
rect 47196 104695 47230 104729
rect 47196 104627 47230 104661
rect 47196 104559 47230 104593
rect 47196 104491 47230 104525
rect 47196 104423 47230 104457
rect 47196 104355 47230 104389
rect 47196 104287 47230 104321
rect 47196 104219 47230 104253
rect 47196 104151 47230 104185
rect 47196 104083 47230 104117
rect 47196 104015 47230 104049
rect 47196 103947 47230 103981
rect 47196 103879 47230 103913
rect 47196 103811 47230 103845
rect 47196 103743 47230 103777
rect 47196 103675 47230 103709
rect 47196 103607 47230 103641
rect 47196 103539 47230 103573
rect 47196 103471 47230 103505
rect 47196 103403 47230 103437
rect 47196 103335 47230 103369
rect 47196 103267 47230 103301
rect 47196 103199 47230 103233
rect 47196 103131 47230 103165
rect 47196 103063 47230 103097
rect 47196 102995 47230 103029
rect 47196 102927 47230 102961
rect 47196 102859 47230 102893
rect 47196 102791 47230 102825
rect 47196 102723 47230 102757
rect 47196 102655 47230 102689
rect 47196 102587 47230 102621
rect 47196 102519 47230 102553
rect 47196 102451 47230 102485
rect 47196 102383 47230 102417
rect 47196 102315 47230 102349
rect 47196 102247 47230 102281
rect 47196 102179 47230 102213
rect 47196 102111 47230 102145
rect 47196 102043 47230 102077
rect 47196 101975 47230 102009
rect 47196 101907 47230 101941
rect 47196 101839 47230 101873
rect 47196 101771 47230 101805
rect 47196 101703 47230 101737
rect 47196 101635 47230 101669
rect 47196 101567 47230 101601
rect 47196 101499 47230 101533
rect 47196 101431 47230 101465
rect 47196 101363 47230 101397
rect 47196 101295 47230 101329
rect 47196 101227 47230 101261
rect 47196 101159 47230 101193
rect 47196 101091 47230 101125
rect 47196 101023 47230 101057
rect 47196 100955 47230 100989
rect -2318 100869 -2284 100903
rect -2250 100869 -2216 100903
rect -2182 100869 -2148 100903
rect -2114 100869 -2080 100903
rect -2046 100869 -2012 100903
rect -1978 100869 -1944 100903
rect -1910 100869 -1876 100903
rect -1842 100869 -1808 100903
rect -1774 100869 -1740 100903
rect -1706 100869 -1672 100903
rect -1638 100869 -1604 100903
rect -1570 100869 -1536 100903
rect -1502 100869 -1468 100903
rect -1434 100869 -1400 100903
rect -1366 100869 -1332 100903
rect -1298 100869 -1264 100903
rect -1230 100869 -1196 100903
rect -1162 100869 -1128 100903
rect -1094 100869 -1060 100903
rect -1026 100869 -992 100903
rect -958 100869 -924 100903
rect -890 100869 -856 100903
rect -822 100869 -788 100903
rect -754 100869 -720 100903
rect -686 100869 -652 100903
rect -618 100869 -584 100903
rect -550 100869 -516 100903
rect -482 100869 -448 100903
rect -414 100869 -380 100903
rect -346 100869 -312 100903
rect -278 100869 -244 100903
rect -210 100869 -176 100903
rect -142 100869 -108 100903
rect -74 100869 -40 100903
rect -6 100869 28 100903
rect 62 100869 96 100903
rect 130 100869 164 100903
rect 198 100869 232 100903
rect 266 100869 300 100903
rect 334 100869 368 100903
rect 402 100869 436 100903
rect 470 100869 504 100903
rect 538 100869 572 100903
rect 606 100869 640 100903
rect 674 100869 708 100903
rect 742 100869 776 100903
rect 810 100869 844 100903
rect 878 100869 912 100903
rect 946 100869 980 100903
rect 1014 100869 1048 100903
rect 1082 100869 1116 100903
rect 1150 100869 1184 100903
rect 1218 100869 1252 100903
rect 1286 100869 1320 100903
rect 1354 100869 1388 100903
rect 1422 100869 1456 100903
rect 1490 100869 1524 100903
rect 1558 100869 1592 100903
rect 1626 100869 1660 100903
rect 1694 100869 1728 100903
rect 1762 100869 1796 100903
rect 1830 100869 1864 100903
rect 1898 100869 1932 100903
rect 1966 100869 2000 100903
rect 2034 100869 2068 100903
rect 2102 100869 2136 100903
rect 2170 100869 2204 100903
rect 2238 100869 2272 100903
rect 2306 100869 2340 100903
rect 2374 100869 2408 100903
rect 2442 100869 2476 100903
rect 2510 100869 2544 100903
rect 2578 100869 2612 100903
rect 2646 100869 2680 100903
rect 2714 100869 2748 100903
rect 2782 100869 2816 100903
rect 2850 100869 2884 100903
rect 2918 100869 2952 100903
rect 2986 100869 3020 100903
rect 3054 100869 3088 100903
rect 3122 100869 3156 100903
rect 3190 100869 3224 100903
rect 3258 100869 3292 100903
rect 3326 100869 3360 100903
rect 3394 100869 3428 100903
rect 3462 100869 3496 100903
rect 3530 100869 3564 100903
rect 3598 100869 3632 100903
rect 3666 100869 3700 100903
rect 3734 100869 3768 100903
rect 3802 100869 3836 100903
rect 3870 100869 3904 100903
rect 3938 100869 3972 100903
rect 4006 100869 4040 100903
rect 4074 100869 4108 100903
rect 4142 100869 4176 100903
rect 4210 100869 4244 100903
rect 4278 100869 4312 100903
rect 4346 100869 4380 100903
rect 4414 100869 4448 100903
rect 4482 100869 4516 100903
rect 4550 100869 4584 100903
rect 4618 100869 4652 100903
rect 4686 100869 4720 100903
rect 4754 100869 4788 100903
rect 4822 100869 4856 100903
rect 4890 100869 4924 100903
rect 4958 100869 4992 100903
rect 5026 100869 5060 100903
rect 5094 100869 5128 100903
rect 5162 100869 5196 100903
rect 5230 100869 5264 100903
rect 5298 100869 5332 100903
rect 5366 100869 5400 100903
rect 5434 100869 5468 100903
rect 5502 100869 5536 100903
rect 5570 100869 5604 100903
rect 5638 100869 5672 100903
rect 5706 100869 5740 100903
rect 5774 100869 5808 100903
rect 5842 100869 5876 100903
rect 5910 100869 5944 100903
rect 5978 100869 6012 100903
rect 6046 100869 6080 100903
rect 6114 100869 6148 100903
rect 6182 100869 6216 100903
rect 6250 100869 6284 100903
rect 6318 100869 6352 100903
rect 6386 100869 6420 100903
rect 6454 100869 6488 100903
rect 6522 100869 6556 100903
rect 6590 100869 6624 100903
rect 6658 100869 6692 100903
rect 6726 100869 6760 100903
rect 6794 100869 6828 100903
rect 6862 100869 6896 100903
rect 6930 100869 6964 100903
rect 6998 100869 7032 100903
rect 7066 100869 7100 100903
rect 7134 100869 7168 100903
rect 7202 100869 7236 100903
rect 7270 100869 7304 100903
rect 7338 100869 7372 100903
rect 7406 100869 7440 100903
rect 7474 100869 7508 100903
rect 7542 100869 7576 100903
rect 7610 100869 7644 100903
rect 7678 100869 7712 100903
rect 7746 100869 7780 100903
rect 7814 100869 7848 100903
rect 7882 100869 7916 100903
rect 7950 100869 7984 100903
rect 8018 100869 8052 100903
rect 8086 100869 8120 100903
rect 8154 100869 8188 100903
rect 8222 100869 8256 100903
rect 8290 100869 8324 100903
rect 8358 100869 8392 100903
rect 8426 100869 8460 100903
rect 8494 100869 8528 100903
rect 8562 100869 8596 100903
rect 8630 100869 8664 100903
rect 8698 100869 8732 100903
rect 8766 100869 8800 100903
rect 8834 100869 8868 100903
rect 8902 100869 8936 100903
rect 8970 100869 9004 100903
rect 9038 100869 9072 100903
rect 9106 100869 9140 100903
rect 9174 100869 9208 100903
rect 9242 100869 9276 100903
rect 9310 100869 9344 100903
rect 9378 100869 9412 100903
rect 9446 100869 9480 100903
rect 9514 100869 9548 100903
rect 9582 100869 9616 100903
rect 9650 100869 9684 100903
rect 9718 100869 9752 100903
rect 9786 100869 9820 100903
rect 9854 100869 9888 100903
rect 9922 100869 9956 100903
rect 9990 100869 10024 100903
rect 10058 100869 10092 100903
rect 10126 100869 10160 100903
rect 10194 100869 10228 100903
rect 10262 100869 10296 100903
rect 10330 100869 10364 100903
rect 10398 100869 10432 100903
rect 10466 100869 10500 100903
rect 10534 100869 10568 100903
rect 10602 100869 10636 100903
rect 10670 100869 10704 100903
rect 10738 100869 10772 100903
rect 10806 100869 10840 100903
rect 10874 100869 10908 100903
rect 10942 100869 10976 100903
rect 11010 100869 11044 100903
rect 11078 100869 11112 100903
rect 11146 100869 11180 100903
rect 11214 100869 11248 100903
rect 11282 100869 11316 100903
rect 11350 100869 11384 100903
rect 11418 100869 11452 100903
rect 11486 100869 11520 100903
rect 11554 100869 11588 100903
rect 11622 100869 11656 100903
rect 11690 100869 11724 100903
rect 11758 100869 11792 100903
rect 11826 100869 11860 100903
rect 11894 100869 11928 100903
rect 11962 100869 11996 100903
rect 12030 100869 12064 100903
rect 12098 100869 12132 100903
rect 12166 100869 12200 100903
rect 12234 100869 12268 100903
rect 12302 100869 12336 100903
rect 12370 100869 12404 100903
rect 12438 100869 12472 100903
rect 12506 100869 12540 100903
rect 12574 100869 12608 100903
rect 12642 100869 12676 100903
rect 12710 100869 12744 100903
rect 12778 100869 12812 100903
rect 12846 100869 12880 100903
rect 12914 100869 12948 100903
rect 12982 100869 13016 100903
rect 13050 100869 13084 100903
rect 13118 100869 13152 100903
rect 13186 100869 13220 100903
rect 13254 100869 13288 100903
rect 13322 100869 13356 100903
rect 13390 100869 13424 100903
rect 13458 100869 13492 100903
rect 13526 100869 13560 100903
rect 13594 100869 13628 100903
rect 13662 100869 13696 100903
rect 13730 100869 13764 100903
rect 13798 100869 13832 100903
rect 13866 100869 13900 100903
rect 13934 100869 13968 100903
rect 14002 100869 14036 100903
rect 14070 100869 14104 100903
rect 14138 100869 14172 100903
rect 14206 100869 14240 100903
rect 14274 100869 14308 100903
rect 14342 100869 14376 100903
rect 14410 100869 14444 100903
rect 14478 100869 14512 100903
rect 14546 100869 14580 100903
rect 14614 100869 14648 100903
rect 14682 100869 14716 100903
rect 14750 100869 14784 100903
rect 14818 100869 14852 100903
rect 14886 100869 14920 100903
rect 14954 100869 14988 100903
rect 15022 100869 15056 100903
rect 15090 100869 15124 100903
rect 15158 100869 15192 100903
rect 15226 100869 15260 100903
rect 15294 100869 15328 100903
rect 15362 100869 15396 100903
rect 15430 100869 15464 100903
rect 15498 100869 15532 100903
rect 15566 100869 15600 100903
rect 15634 100869 15668 100903
rect 15702 100869 15736 100903
rect 15770 100869 15804 100903
rect 15838 100869 15872 100903
rect 15906 100869 15940 100903
rect 15974 100869 16008 100903
rect 16042 100869 16076 100903
rect 16110 100869 16144 100903
rect 16178 100869 16212 100903
rect 16246 100869 16280 100903
rect 16314 100869 16348 100903
rect 16382 100869 16416 100903
rect 16450 100869 16484 100903
rect 16518 100869 16552 100903
rect 16586 100869 16620 100903
rect 16654 100869 16688 100903
rect 16722 100869 16756 100903
rect 16790 100869 16824 100903
rect 16858 100869 16892 100903
rect 16926 100869 16960 100903
rect 16994 100869 17028 100903
rect 17062 100869 17096 100903
rect 17130 100869 17164 100903
rect 17198 100869 17232 100903
rect 17266 100869 17300 100903
rect 17334 100869 17368 100903
rect 17402 100869 17436 100903
rect 17470 100869 17504 100903
rect 17538 100869 17572 100903
rect 17606 100869 17640 100903
rect 17674 100869 17708 100903
rect 17742 100869 17776 100903
rect 17810 100869 17844 100903
rect 17878 100869 17912 100903
rect 17946 100869 17980 100903
rect 18014 100869 18048 100903
rect 18082 100869 18116 100903
rect 18150 100869 18184 100903
rect 18218 100869 18252 100903
rect 18286 100869 18320 100903
rect 18354 100869 18388 100903
rect 18422 100869 18456 100903
rect 18490 100869 18524 100903
rect 18558 100869 18592 100903
rect 18626 100869 18660 100903
rect 18694 100869 18728 100903
rect 18762 100869 18796 100903
rect 18830 100869 18864 100903
rect 18898 100869 18932 100903
rect 18966 100869 19000 100903
rect 19034 100869 19068 100903
rect 19102 100869 19136 100903
rect 19170 100869 19204 100903
rect 19238 100869 19272 100903
rect 19306 100869 19340 100903
rect 19374 100869 19408 100903
rect 19442 100869 19476 100903
rect 19510 100869 19544 100903
rect 19578 100869 19612 100903
rect 19646 100869 19680 100903
rect 19714 100869 19748 100903
rect 19782 100869 19816 100903
rect 19850 100869 19884 100903
rect 19918 100869 19952 100903
rect 19986 100869 20020 100903
rect 20054 100869 20088 100903
rect 20122 100869 20156 100903
rect 20190 100869 20224 100903
rect 20258 100869 20292 100903
rect 20326 100869 20360 100903
rect 20394 100869 20428 100903
rect 20462 100869 20496 100903
rect 20530 100869 20564 100903
rect 20598 100869 20632 100903
rect 20666 100869 20700 100903
rect 20734 100869 20768 100903
rect 20802 100869 20836 100903
rect 20870 100869 20904 100903
rect 20938 100869 20972 100903
rect 21006 100869 21040 100903
rect 21074 100869 21108 100903
rect 21142 100869 21176 100903
rect 21210 100869 21244 100903
rect 21278 100869 21312 100903
rect 21346 100869 21380 100903
rect 21414 100869 21448 100903
rect 21482 100869 21516 100903
rect 21550 100869 21584 100903
rect 21618 100869 21652 100903
rect 21686 100869 21720 100903
rect 21754 100869 21788 100903
rect 21822 100869 21856 100903
rect 21890 100869 21924 100903
rect 21958 100869 21992 100903
rect 22026 100869 22060 100903
rect 22094 100869 22128 100903
rect 22162 100869 22196 100903
rect 22230 100869 22264 100903
rect 22298 100869 22332 100903
rect 22366 100869 22400 100903
rect 22434 100869 22468 100903
rect 22502 100869 22536 100903
rect 22570 100869 22604 100903
rect 22638 100869 22672 100903
rect 22706 100869 22740 100903
rect 22774 100869 22808 100903
rect 22842 100869 22876 100903
rect 22910 100869 22944 100903
rect 22978 100869 23012 100903
rect 23046 100869 23080 100903
rect 23114 100869 23148 100903
rect 23182 100869 23216 100903
rect 23250 100869 23284 100903
rect 23318 100869 23352 100903
rect 23386 100869 23420 100903
rect 23454 100869 23488 100903
rect 23522 100869 23556 100903
rect 23590 100869 23624 100903
rect 23658 100869 23692 100903
rect 23726 100869 23760 100903
rect 23794 100869 23828 100903
rect 23862 100869 23896 100903
rect 23930 100869 23964 100903
rect 23998 100869 24032 100903
rect 24066 100869 24100 100903
rect 24134 100869 24168 100903
rect 24202 100869 24236 100903
rect 24270 100869 24304 100903
rect 24338 100869 24372 100903
rect 24406 100869 24440 100903
rect 24474 100869 24508 100903
rect 24542 100869 24576 100903
rect 24610 100869 24644 100903
rect 24678 100869 24712 100903
rect 24746 100869 24780 100903
rect 24814 100869 24848 100903
rect 24882 100869 24916 100903
rect 24950 100869 24984 100903
rect 25018 100869 25052 100903
rect 25086 100869 25120 100903
rect 25154 100869 25188 100903
rect 25222 100869 25256 100903
rect 25290 100869 25324 100903
rect 25358 100869 25392 100903
rect 25426 100869 25460 100903
rect 25494 100869 25528 100903
rect 25562 100869 25596 100903
rect 25630 100869 25664 100903
rect 25698 100869 25732 100903
rect 25766 100869 25800 100903
rect 25834 100869 25868 100903
rect 25902 100869 25936 100903
rect 25970 100869 26004 100903
rect 26038 100869 26072 100903
rect 26106 100869 26140 100903
rect 26174 100869 26208 100903
rect 26242 100869 26276 100903
rect 26310 100869 26344 100903
rect 26378 100869 26412 100903
rect 26446 100869 26480 100903
rect 26514 100869 26548 100903
rect 26582 100869 26616 100903
rect 26650 100869 26684 100903
rect 26718 100869 26752 100903
rect 26786 100869 26820 100903
rect 26854 100869 26888 100903
rect 26922 100869 26956 100903
rect 26990 100869 27024 100903
rect 27058 100869 27092 100903
rect 27126 100869 27160 100903
rect 27194 100869 27228 100903
rect 27262 100869 27296 100903
rect 27330 100869 27364 100903
rect 27398 100869 27432 100903
rect 27466 100869 27500 100903
rect 27534 100869 27568 100903
rect 27602 100869 27636 100903
rect 27670 100869 27704 100903
rect 27738 100869 27772 100903
rect 27806 100869 27840 100903
rect 27874 100869 27908 100903
rect 27942 100869 27976 100903
rect 28010 100869 28044 100903
rect 28078 100869 28112 100903
rect 28146 100869 28180 100903
rect 28214 100869 28248 100903
rect 28282 100869 28316 100903
rect 28350 100869 28384 100903
rect 28418 100869 28452 100903
rect 28486 100869 28520 100903
rect 28554 100869 28588 100903
rect 28622 100869 28656 100903
rect 28690 100869 28724 100903
rect 28758 100869 28792 100903
rect 28826 100869 28860 100903
rect 28894 100869 28928 100903
rect 28962 100869 28996 100903
rect 29030 100869 29064 100903
rect 29098 100869 29132 100903
rect 29166 100869 29200 100903
rect 29234 100869 29268 100903
rect 29302 100869 29336 100903
rect 29370 100869 29404 100903
rect 29438 100869 29472 100903
rect 29506 100869 29540 100903
rect 29574 100869 29608 100903
rect 29642 100869 29676 100903
rect 29710 100869 29744 100903
rect 29778 100869 29812 100903
rect 29846 100869 29880 100903
rect 29914 100869 29948 100903
rect 29982 100869 30016 100903
rect 30050 100869 30084 100903
rect 30118 100869 30152 100903
rect 30186 100869 30220 100903
rect 30254 100869 30288 100903
rect 30322 100869 30356 100903
rect 30390 100869 30424 100903
rect 30458 100869 30492 100903
rect 30526 100869 30560 100903
rect 30594 100869 30628 100903
rect 30662 100869 30696 100903
rect 30730 100869 30764 100903
rect 30798 100869 30832 100903
rect 30866 100869 30900 100903
rect 30934 100869 30968 100903
rect 31002 100869 31036 100903
rect 31070 100869 31104 100903
rect 31138 100869 31172 100903
rect 31206 100869 31240 100903
rect 31274 100869 31308 100903
rect 31342 100869 31376 100903
rect 31410 100869 31444 100903
rect 31478 100869 31512 100903
rect 31546 100869 31580 100903
rect 31614 100869 31648 100903
rect 31682 100869 31716 100903
rect 31750 100869 31784 100903
rect 31818 100869 31852 100903
rect 31886 100869 31920 100903
rect 31954 100869 31988 100903
rect 32022 100869 32056 100903
rect 32090 100869 32124 100903
rect 32158 100869 32192 100903
rect 32226 100869 32260 100903
rect 32294 100869 32328 100903
rect 32362 100869 32396 100903
rect 32430 100869 32464 100903
rect 32498 100869 32532 100903
rect 32566 100869 32600 100903
rect 32634 100869 32668 100903
rect 32702 100869 32736 100903
rect 32770 100869 32804 100903
rect 32838 100869 32872 100903
rect 32906 100869 32940 100903
rect 32974 100869 33008 100903
rect 33042 100869 33076 100903
rect 33110 100869 33144 100903
rect 33178 100869 33212 100903
rect 33246 100869 33280 100903
rect 33314 100869 33348 100903
rect 33382 100869 33416 100903
rect 33450 100869 33484 100903
rect 33518 100869 33552 100903
rect 33586 100869 33620 100903
rect 33654 100869 33688 100903
rect 33722 100869 33756 100903
rect 33790 100869 33824 100903
rect 33858 100869 33892 100903
rect 33926 100869 33960 100903
rect 33994 100869 34028 100903
rect 34062 100869 34096 100903
rect 34130 100869 34164 100903
rect 34198 100869 34232 100903
rect 34266 100869 34300 100903
rect 34334 100869 34368 100903
rect 34402 100869 34436 100903
rect 34470 100869 34504 100903
rect 34538 100869 34572 100903
rect 34606 100869 34640 100903
rect 34674 100869 34708 100903
rect 34742 100869 34776 100903
rect 34810 100869 34844 100903
rect 34878 100869 34912 100903
rect 34946 100869 34980 100903
rect 35014 100869 35048 100903
rect 35082 100869 35116 100903
rect 35150 100869 35184 100903
rect 35218 100869 35252 100903
rect 35286 100869 35320 100903
rect 35354 100869 35388 100903
rect 35422 100869 35456 100903
rect 35490 100869 35524 100903
rect 35558 100869 35592 100903
rect 35626 100869 35660 100903
rect 35694 100869 35728 100903
rect 35762 100869 35796 100903
rect 35830 100869 35864 100903
rect 35898 100869 35932 100903
rect 35966 100869 36000 100903
rect 36034 100869 36068 100903
rect 36102 100869 36136 100903
rect 36170 100869 36204 100903
rect 36238 100869 36272 100903
rect 36306 100869 36340 100903
rect 36374 100869 36408 100903
rect 36442 100869 36476 100903
rect 36510 100869 36544 100903
rect 36578 100869 36612 100903
rect 36646 100869 36680 100903
rect 36714 100869 36748 100903
rect 36782 100869 36816 100903
rect 36850 100869 36884 100903
rect 36918 100869 36952 100903
rect 36986 100869 37020 100903
rect 37054 100869 37088 100903
rect 37122 100869 37156 100903
rect 37190 100869 37224 100903
rect 37258 100869 37292 100903
rect 37326 100869 37360 100903
rect 37394 100869 37428 100903
rect 37462 100869 37496 100903
rect 37530 100869 37564 100903
rect 37598 100869 37632 100903
rect 37666 100869 37700 100903
rect 37734 100869 37768 100903
rect 37802 100869 37836 100903
rect 37870 100869 37904 100903
rect 37938 100869 37972 100903
rect 38006 100869 38040 100903
rect 38074 100869 38108 100903
rect 38142 100869 38176 100903
rect 38210 100869 38244 100903
rect 38278 100869 38312 100903
rect 38346 100869 38380 100903
rect 38414 100869 38448 100903
rect 38482 100869 38516 100903
rect 38550 100869 38584 100903
rect 38618 100869 38652 100903
rect 38686 100869 38720 100903
rect 38754 100869 38788 100903
rect 38822 100869 38856 100903
rect 38890 100869 38924 100903
rect 38958 100869 38992 100903
rect 39026 100869 39060 100903
rect 39094 100869 39128 100903
rect 39162 100869 39196 100903
rect 39230 100869 39264 100903
rect 39298 100869 39332 100903
rect 39366 100869 39400 100903
rect 39434 100869 39468 100903
rect 39502 100869 39536 100903
rect 39570 100869 39604 100903
rect 39638 100869 39672 100903
rect 39706 100869 39740 100903
rect 39774 100869 39808 100903
rect 39842 100869 39876 100903
rect 39910 100869 39944 100903
rect 39978 100869 40012 100903
rect 40046 100869 40080 100903
rect 40114 100869 40148 100903
rect 40182 100869 40216 100903
rect 40250 100869 40284 100903
rect 40318 100869 40352 100903
rect 40386 100869 40420 100903
rect 40454 100869 40488 100903
rect 40522 100869 40556 100903
rect 40590 100869 40624 100903
rect 40658 100869 40692 100903
rect 40726 100869 40760 100903
rect 40794 100869 40828 100903
rect 40862 100869 40896 100903
rect 40930 100869 40964 100903
rect 40998 100869 41032 100903
rect 41066 100869 41100 100903
rect 41134 100869 41168 100903
rect 41202 100869 41236 100903
rect 41270 100869 41304 100903
rect 41338 100869 41372 100903
rect 41406 100869 41440 100903
rect 41474 100869 41508 100903
rect 41542 100869 41576 100903
rect 41610 100869 41644 100903
rect 41678 100869 41712 100903
rect 41746 100869 41780 100903
rect 41814 100869 41848 100903
rect 41882 100869 41916 100903
rect 41950 100869 41984 100903
rect 42018 100869 42052 100903
rect 42086 100869 42120 100903
rect 42154 100869 42188 100903
rect 42222 100869 42256 100903
rect 42290 100869 42324 100903
rect 42358 100869 42392 100903
rect 42426 100869 42460 100903
rect 42494 100869 42528 100903
rect 42562 100869 42596 100903
rect 42630 100869 42664 100903
rect 42698 100869 42732 100903
rect 42766 100869 42800 100903
rect 42834 100869 42868 100903
rect 42902 100869 42936 100903
rect 42970 100869 43004 100903
rect 43038 100869 43072 100903
rect 43106 100869 43140 100903
rect 43174 100869 43208 100903
rect 43242 100869 43276 100903
rect 43310 100869 43344 100903
rect 43378 100869 43412 100903
rect 43446 100869 43480 100903
rect 43514 100869 43548 100903
rect 43582 100869 43616 100903
rect 43650 100869 43684 100903
rect 43718 100869 43752 100903
rect 43786 100869 43820 100903
rect 43854 100869 43888 100903
rect 43922 100869 43956 100903
rect 43990 100869 44024 100903
rect 44058 100869 44092 100903
rect 44126 100869 44160 100903
rect 44194 100869 44228 100903
rect 44262 100869 44296 100903
rect 44330 100869 44364 100903
rect 44398 100869 44432 100903
rect 44466 100869 44500 100903
rect 44534 100869 44568 100903
rect 44602 100869 44636 100903
rect 44670 100869 44704 100903
rect 44738 100869 44772 100903
rect 44806 100869 44840 100903
rect 44874 100869 44908 100903
rect 44942 100869 44976 100903
rect 45010 100869 45044 100903
rect 45078 100869 45112 100903
rect 45146 100869 45180 100903
rect 45214 100869 45248 100903
rect 45282 100869 45316 100903
rect 45350 100869 45384 100903
rect 45418 100869 45452 100903
rect 45486 100869 45520 100903
rect 45554 100869 45588 100903
rect 45622 100869 45656 100903
rect 45690 100869 45724 100903
rect 45758 100869 45792 100903
rect 45826 100869 45860 100903
rect 45894 100869 45928 100903
rect 45962 100869 45996 100903
rect 46030 100869 46064 100903
rect 46098 100869 46132 100903
rect 46166 100869 46200 100903
rect 46234 100869 46268 100903
rect 46302 100869 46336 100903
rect 46370 100869 46404 100903
rect 46438 100869 46472 100903
rect 46506 100869 46540 100903
rect 46574 100869 46608 100903
rect 46642 100869 46676 100903
rect 46710 100869 46744 100903
rect 46778 100869 46812 100903
rect 46846 100869 46880 100903
rect 46914 100869 46948 100903
rect 46982 100869 47016 100903
rect 47050 100869 47084 100903
rect 47118 100869 47152 100903
rect -10609 76110 -10575 76144
rect -10541 76110 -10507 76144
rect -10473 76110 -10439 76144
rect -10405 76110 -10371 76144
rect -10337 76110 -10303 76144
rect -10269 76110 -10235 76144
rect -10201 76110 -10167 76144
rect -10133 76110 -10099 76144
rect -10065 76110 -10031 76144
rect -9997 76110 -9963 76144
rect -9929 76110 -9895 76144
rect -9861 76110 -9827 76144
rect -9793 76110 -9759 76144
rect -9725 76110 -9691 76144
rect -9657 76110 -9623 76144
rect -9589 76110 -9555 76144
rect -9521 76110 -9487 76144
rect -9453 76110 -9419 76144
rect -9385 76110 -9351 76144
rect -9317 76110 -9283 76144
rect -9249 76110 -9215 76144
rect -9181 76110 -9147 76144
rect -9113 76110 -9079 76144
rect -9045 76110 -9011 76144
rect -8977 76110 -8943 76144
rect -8909 76110 -8875 76144
rect -8841 76110 -8807 76144
rect -8773 76110 -8739 76144
rect -8705 76110 -8671 76144
rect -8637 76110 -8603 76144
rect -8569 76110 -8535 76144
rect -8501 76110 -8467 76144
rect -8433 76110 -8399 76144
rect -8365 76110 -8331 76144
rect -8297 76110 -8263 76144
rect -8229 76110 -8195 76144
rect -8161 76110 -8127 76144
rect -8093 76110 -8059 76144
rect -8025 76110 -7991 76144
rect -7957 76110 -7923 76144
rect -7889 76110 -7855 76144
rect -7821 76110 -7787 76144
rect -7753 76110 -7719 76144
rect -7685 76110 -7651 76144
rect -7617 76110 -7583 76144
rect -7549 76110 -7515 76144
rect -7481 76110 -7447 76144
rect -7413 76110 -7379 76144
rect -7345 76110 -7311 76144
rect -7277 76110 -7243 76144
rect -7209 76110 -7175 76144
rect -7141 76110 -7107 76144
rect -7073 76110 -7039 76144
rect -7005 76110 -6971 76144
rect -6937 76110 -6903 76144
rect -6869 76110 -6835 76144
rect -6801 76110 -6767 76144
rect -6733 76110 -6699 76144
rect -6665 76110 -6631 76144
rect -6597 76110 -6563 76144
rect -6529 76110 -6495 76144
rect -6461 76110 -6427 76144
rect -6393 76110 -6359 76144
rect -6325 76110 -6291 76144
rect -6257 76110 -6223 76144
rect -6189 76110 -6155 76144
rect -6121 76110 -6087 76144
rect -6053 76110 -6019 76144
rect -5985 76110 -5951 76144
rect -5917 76110 -5883 76144
rect -5849 76110 -5815 76144
rect -5781 76110 -5747 76144
rect -5713 76110 -5679 76144
rect -5645 76110 -5611 76144
rect -5577 76110 -5543 76144
rect -5509 76110 -5475 76144
rect -5441 76110 -5407 76144
rect -5373 76110 -5339 76144
rect -5305 76110 -5271 76144
rect -5237 76110 -5203 76144
rect -5169 76110 -5135 76144
rect -5101 76110 -5067 76144
rect -5033 76110 -4999 76144
rect -4965 76110 -4931 76144
rect -4897 76110 -4863 76144
rect -4829 76110 -4795 76144
rect -4761 76110 -4727 76144
rect -4693 76110 -4659 76144
rect -4625 76110 -4591 76144
rect -4557 76110 -4523 76144
rect -4489 76110 -4455 76144
rect -4421 76110 -4387 76144
rect -4353 76110 -4319 76144
rect -4285 76110 -4251 76144
rect -4217 76110 -4183 76144
rect -4149 76110 -4115 76144
rect -4081 76110 -4047 76144
rect -4013 76110 -3979 76144
rect -3945 76110 -3911 76144
rect -3877 76110 -3843 76144
rect -3809 76110 -3775 76144
rect -10699 76050 -10665 76084
rect -10699 75982 -10665 76016
rect -10699 75914 -10665 75948
rect -10699 75846 -10665 75880
rect -10699 75778 -10665 75812
rect -10699 75710 -10665 75744
rect -10699 75642 -10665 75676
rect -10699 75574 -10665 75608
rect -10699 75506 -10665 75540
rect -10699 75438 -10665 75472
rect -10699 75370 -10665 75404
rect -10699 75302 -10665 75336
rect -10699 75234 -10665 75268
rect -10699 75166 -10665 75200
rect -10699 75098 -10665 75132
rect -10699 75030 -10665 75064
rect -10699 74962 -10665 74996
rect -10699 74894 -10665 74928
rect -10699 74826 -10665 74860
rect -10699 74758 -10665 74792
rect -10699 74690 -10665 74724
rect -10699 74622 -10665 74656
rect -10699 74554 -10665 74588
rect -10699 74486 -10665 74520
rect -10699 74418 -10665 74452
rect -10699 74350 -10665 74384
rect -10699 74282 -10665 74316
rect -10699 74214 -10665 74248
rect -10699 74146 -10665 74180
rect -10699 74078 -10665 74112
rect -10699 74010 -10665 74044
rect -10699 73942 -10665 73976
rect -10699 73874 -10665 73908
rect -10699 73806 -10665 73840
rect -10699 73738 -10665 73772
rect -10699 73670 -10665 73704
rect -10699 73602 -10665 73636
rect -10699 73534 -10665 73568
rect -10699 73466 -10665 73500
rect -10699 73398 -10665 73432
rect -10699 73330 -10665 73364
rect -10699 73262 -10665 73296
rect -10699 73194 -10665 73228
rect -10699 73126 -10665 73160
rect -10699 73058 -10665 73092
rect -10699 72990 -10665 73024
rect -10699 72922 -10665 72956
rect -10699 72854 -10665 72888
rect -10699 72786 -10665 72820
rect -10699 72718 -10665 72752
rect -10699 72650 -10665 72684
rect -10699 72582 -10665 72616
rect -10699 72514 -10665 72548
rect -10699 72446 -10665 72480
rect -10699 72378 -10665 72412
rect -10699 72310 -10665 72344
rect -10699 72242 -10665 72276
rect -10699 72174 -10665 72208
rect -10699 72106 -10665 72140
rect -10699 72038 -10665 72072
rect -10699 71970 -10665 72004
rect -10699 71902 -10665 71936
rect -10699 71834 -10665 71868
rect -10699 71766 -10665 71800
rect -10699 71698 -10665 71732
rect -10699 71630 -10665 71664
rect -10699 71562 -10665 71596
rect -10699 71494 -10665 71528
rect -10699 71426 -10665 71460
rect -10699 71358 -10665 71392
rect -10699 71290 -10665 71324
rect -10699 71222 -10665 71256
rect -10699 71154 -10665 71188
rect -10699 71086 -10665 71120
rect -10699 71018 -10665 71052
rect -10699 70950 -10665 70984
rect -10699 70882 -10665 70916
rect -10699 70814 -10665 70848
rect -10699 70746 -10665 70780
rect -10699 70678 -10665 70712
rect -10699 70610 -10665 70644
rect -10699 70542 -10665 70576
rect -10699 70474 -10665 70508
rect -10699 70406 -10665 70440
rect -10699 70338 -10665 70372
rect -10699 70270 -10665 70304
rect -10699 70202 -10665 70236
rect -10699 70134 -10665 70168
rect -10699 70066 -10665 70100
rect -10699 69998 -10665 70032
rect -10699 69930 -10665 69964
rect -10699 69862 -10665 69896
rect -10699 69794 -10665 69828
rect -10699 69726 -10665 69760
rect -10699 69658 -10665 69692
rect -10699 69590 -10665 69624
rect -10699 69522 -10665 69556
rect -10699 69454 -10665 69488
rect -10699 69386 -10665 69420
rect -10699 69318 -10665 69352
rect -10699 69250 -10665 69284
rect -10699 69182 -10665 69216
rect -10699 69114 -10665 69148
rect -10699 69046 -10665 69080
rect -10699 68978 -10665 69012
rect -10699 68910 -10665 68944
rect -10699 68842 -10665 68876
rect -10699 68774 -10665 68808
rect -10699 68706 -10665 68740
rect -10699 68638 -10665 68672
rect -10699 68570 -10665 68604
rect -10699 68502 -10665 68536
rect -10699 68434 -10665 68468
rect -10699 68366 -10665 68400
rect -10699 68298 -10665 68332
rect -10699 68230 -10665 68264
rect -10699 68162 -10665 68196
rect -10699 68094 -10665 68128
rect -10699 68026 -10665 68060
rect -10699 67958 -10665 67992
rect -10699 67890 -10665 67924
rect -10699 67822 -10665 67856
rect -10699 67754 -10665 67788
rect -10699 67686 -10665 67720
rect -10699 67618 -10665 67652
rect -10699 67550 -10665 67584
rect -10699 67482 -10665 67516
rect -10699 67414 -10665 67448
rect -10699 67346 -10665 67380
rect -10699 67278 -10665 67312
rect -10699 67210 -10665 67244
rect -10699 67142 -10665 67176
rect -10699 67074 -10665 67108
rect -10699 67006 -10665 67040
rect -10699 66938 -10665 66972
rect -10699 66870 -10665 66904
rect -10699 66802 -10665 66836
rect -10699 66734 -10665 66768
rect -10699 66666 -10665 66700
rect -10699 66598 -10665 66632
rect -10699 66530 -10665 66564
rect -10699 66462 -10665 66496
rect -10699 66394 -10665 66428
rect -10699 66326 -10665 66360
rect -10699 66258 -10665 66292
rect -10699 66190 -10665 66224
rect -10699 66122 -10665 66156
rect -10699 66054 -10665 66088
rect -10699 65986 -10665 66020
rect -10699 65918 -10665 65952
rect -10699 65850 -10665 65884
rect -10699 65782 -10665 65816
rect -10699 65714 -10665 65748
rect -10699 65646 -10665 65680
rect -10699 65578 -10665 65612
rect -10699 65510 -10665 65544
rect -10699 65442 -10665 65476
rect -10699 65374 -10665 65408
rect -10699 65306 -10665 65340
rect -10699 65238 -10665 65272
rect -10699 65170 -10665 65204
rect -10699 65102 -10665 65136
rect -10699 65034 -10665 65068
rect -10699 64966 -10665 65000
rect -10699 64898 -10665 64932
rect -10699 64830 -10665 64864
rect -10699 64762 -10665 64796
rect -10699 64694 -10665 64728
rect -10699 64626 -10665 64660
rect -10699 64558 -10665 64592
rect -10699 64490 -10665 64524
rect -10699 64422 -10665 64456
rect -10699 64354 -10665 64388
rect -10699 64286 -10665 64320
rect -10699 64218 -10665 64252
rect -10699 64150 -10665 64184
rect -3718 76022 -3684 76056
rect -3718 75954 -3684 75988
rect -3718 75886 -3684 75920
rect -3718 75818 -3684 75852
rect -3718 75750 -3684 75784
rect -3718 75682 -3684 75716
rect -3718 75614 -3684 75648
rect -3718 75546 -3684 75580
rect -3718 75478 -3684 75512
rect -3718 75410 -3684 75444
rect -3718 75342 -3684 75376
rect -3718 75274 -3684 75308
rect -3718 75206 -3684 75240
rect -3718 75138 -3684 75172
rect -3718 75070 -3684 75104
rect -3718 75002 -3684 75036
rect -3718 74934 -3684 74968
rect -3718 74866 -3684 74900
rect -3718 74798 -3684 74832
rect -3718 74730 -3684 74764
rect -3718 74662 -3684 74696
rect -3718 74594 -3684 74628
rect -3718 74526 -3684 74560
rect -3718 74458 -3684 74492
rect -3718 74390 -3684 74424
rect -3718 74322 -3684 74356
rect -3718 74254 -3684 74288
rect -3718 74186 -3684 74220
rect -3718 74118 -3684 74152
rect -3718 74050 -3684 74084
rect -3718 73982 -3684 74016
rect -3718 73914 -3684 73948
rect -3718 73846 -3684 73880
rect -3718 73778 -3684 73812
rect -3718 73710 -3684 73744
rect -3718 73642 -3684 73676
rect -3718 73574 -3684 73608
rect -3718 73506 -3684 73540
rect -3718 73438 -3684 73472
rect -3718 73370 -3684 73404
rect -3718 73302 -3684 73336
rect -3718 73234 -3684 73268
rect -3718 73166 -3684 73200
rect -3718 73098 -3684 73132
rect -3718 73030 -3684 73064
rect -3718 72962 -3684 72996
rect -3718 72894 -3684 72928
rect -3718 72826 -3684 72860
rect -3718 72758 -3684 72792
rect -3718 72690 -3684 72724
rect -3718 72622 -3684 72656
rect -3718 72554 -3684 72588
rect -3718 72486 -3684 72520
rect -3718 72418 -3684 72452
rect -3718 72350 -3684 72384
rect -3718 72282 -3684 72316
rect -3718 72214 -3684 72248
rect -3718 72146 -3684 72180
rect -3718 72078 -3684 72112
rect -3718 72010 -3684 72044
rect -3718 71942 -3684 71976
rect -3718 71874 -3684 71908
rect -3718 71806 -3684 71840
rect -3718 71738 -3684 71772
rect -3718 71670 -3684 71704
rect -3718 71602 -3684 71636
rect -3718 71534 -3684 71568
rect -3718 71466 -3684 71500
rect -3718 71398 -3684 71432
rect -3718 71330 -3684 71364
rect -3718 71262 -3684 71296
rect -3718 71194 -3684 71228
rect -3718 71126 -3684 71160
rect -3718 71058 -3684 71092
rect -3718 70990 -3684 71024
rect -3718 70922 -3684 70956
rect -3718 70854 -3684 70888
rect -3718 70786 -3684 70820
rect -3718 70718 -3684 70752
rect -3718 70650 -3684 70684
rect -3718 70582 -3684 70616
rect -3718 70514 -3684 70548
rect -3718 70446 -3684 70480
rect -3718 70378 -3684 70412
rect -3718 70310 -3684 70344
rect -3718 70242 -3684 70276
rect -3718 70174 -3684 70208
rect -3718 70106 -3684 70140
rect -3718 70038 -3684 70072
rect -3718 69970 -3684 70004
rect -3718 69902 -3684 69936
rect -3718 69834 -3684 69868
rect -3718 69766 -3684 69800
rect -3718 69698 -3684 69732
rect -3718 69630 -3684 69664
rect -3718 69562 -3684 69596
rect -3718 69494 -3684 69528
rect -3718 69426 -3684 69460
rect -3718 69358 -3684 69392
rect -3718 69290 -3684 69324
rect -3718 69222 -3684 69256
rect -3718 69154 -3684 69188
rect -3718 69086 -3684 69120
rect -3718 69018 -3684 69052
rect -3718 68950 -3684 68984
rect -3718 68882 -3684 68916
rect -3718 68814 -3684 68848
rect -3718 68746 -3684 68780
rect -3718 68678 -3684 68712
rect -3718 68610 -3684 68644
rect -3718 68542 -3684 68576
rect -3718 68474 -3684 68508
rect -3718 68406 -3684 68440
rect -3718 68338 -3684 68372
rect -3718 68270 -3684 68304
rect -3718 68202 -3684 68236
rect -3718 68134 -3684 68168
rect -3718 68066 -3684 68100
rect -3718 67998 -3684 68032
rect -3718 67930 -3684 67964
rect -3718 67862 -3684 67896
rect -3718 67794 -3684 67828
rect -3718 67726 -3684 67760
rect -3718 67658 -3684 67692
rect -3718 67590 -3684 67624
rect -3718 67522 -3684 67556
rect -3718 67454 -3684 67488
rect -3718 67386 -3684 67420
rect -3718 67318 -3684 67352
rect -3718 67250 -3684 67284
rect -3718 67182 -3684 67216
rect -3718 67114 -3684 67148
rect -3718 67046 -3684 67080
rect -3718 66978 -3684 67012
rect -3718 66910 -3684 66944
rect -3718 66842 -3684 66876
rect -3718 66774 -3684 66808
rect -3718 66706 -3684 66740
rect -3718 66638 -3684 66672
rect -3718 66570 -3684 66604
rect -3718 66502 -3684 66536
rect -3718 66434 -3684 66468
rect -3718 66366 -3684 66400
rect -3718 66298 -3684 66332
rect -3718 66230 -3684 66264
rect -3718 66162 -3684 66196
rect -3718 66094 -3684 66128
rect -3718 66026 -3684 66060
rect -3718 65958 -3684 65992
rect -3718 65890 -3684 65924
rect -3718 65822 -3684 65856
rect -3718 65754 -3684 65788
rect -3718 65686 -3684 65720
rect -3718 65618 -3684 65652
rect -3718 65550 -3684 65584
rect -3718 65482 -3684 65516
rect -3718 65414 -3684 65448
rect -3718 65346 -3684 65380
rect -3718 65278 -3684 65312
rect -3718 65210 -3684 65244
rect -3718 65142 -3684 65176
rect -3718 65074 -3684 65108
rect -3718 65006 -3684 65040
rect -3718 64938 -3684 64972
rect -3718 64870 -3684 64904
rect -3718 64802 -3684 64836
rect -3718 64734 -3684 64768
rect -3718 64666 -3684 64700
rect -3718 64598 -3684 64632
rect -3718 64530 -3684 64564
rect -3718 64462 -3684 64496
rect -3718 64394 -3684 64428
rect -3718 64326 -3684 64360
rect -3718 64258 -3684 64292
rect -3718 64190 -3684 64224
rect -10624 64086 -10590 64120
rect -10556 64086 -10522 64120
rect -10488 64086 -10454 64120
rect -10420 64086 -10386 64120
rect -10352 64086 -10318 64120
rect -10284 64086 -10250 64120
rect -10216 64086 -10182 64120
rect -10148 64086 -10114 64120
rect -10080 64086 -10046 64120
rect -10012 64086 -9978 64120
rect -9944 64086 -9910 64120
rect -9876 64086 -9842 64120
rect -9808 64086 -9774 64120
rect -9740 64086 -9706 64120
rect -9672 64086 -9638 64120
rect -9604 64086 -9570 64120
rect -9536 64086 -9502 64120
rect -9468 64086 -9434 64120
rect -9400 64086 -9366 64120
rect -9332 64086 -9298 64120
rect -9264 64086 -9230 64120
rect -9196 64086 -9162 64120
rect -9128 64086 -9094 64120
rect -9060 64086 -9026 64120
rect -8992 64086 -8958 64120
rect -8924 64086 -8890 64120
rect -8856 64086 -8822 64120
rect -8788 64086 -8754 64120
rect -8720 64086 -8686 64120
rect -8652 64086 -8618 64120
rect -8584 64086 -8550 64120
rect -8516 64086 -8482 64120
rect -8448 64086 -8414 64120
rect -8380 64086 -8346 64120
rect -8312 64086 -8278 64120
rect -8244 64086 -8210 64120
rect -8176 64086 -8142 64120
rect -8108 64086 -8074 64120
rect -8040 64086 -8006 64120
rect -7972 64086 -7938 64120
rect -7904 64086 -7870 64120
rect -7836 64086 -7802 64120
rect -7768 64086 -7734 64120
rect -7700 64086 -7666 64120
rect -7632 64086 -7598 64120
rect -7564 64086 -7530 64120
rect -7496 64086 -7462 64120
rect -7428 64086 -7394 64120
rect -7360 64086 -7326 64120
rect -7292 64086 -7258 64120
rect -7207 64025 -7173 64059
rect -7207 63957 -7173 63991
rect -7207 63889 -7173 63923
rect -7207 63821 -7173 63855
rect -7207 63753 -7173 63787
rect -7207 63685 -7173 63719
rect -7207 63617 -7173 63651
rect -7207 63549 -7173 63583
rect -7207 63481 -7173 63515
rect -7207 63413 -7173 63447
rect -7207 63345 -7173 63379
rect -7207 63277 -7173 63311
rect -7207 63209 -7173 63243
rect -7207 63141 -7173 63175
rect -7207 63073 -7173 63107
rect -7207 63005 -7173 63039
rect -7207 62937 -7173 62971
rect -7207 62869 -7173 62903
rect -7207 62801 -7173 62835
rect -7207 62733 -7173 62767
rect -7207 62665 -7173 62699
rect -7207 62597 -7173 62631
rect -7207 62529 -7173 62563
rect -7207 62461 -7173 62495
rect -7207 62393 -7173 62427
rect -7207 62325 -7173 62359
rect -7207 62257 -7173 62291
rect -7207 62189 -7173 62223
rect -7207 62121 -7173 62155
rect -7207 62053 -7173 62087
rect -7207 61985 -7173 62019
rect -7207 61917 -7173 61951
rect -7207 61849 -7173 61883
rect -7207 61781 -7173 61815
rect -7207 61713 -7173 61747
rect -7207 61645 -7173 61679
rect -7207 61577 -7173 61611
rect -7207 61509 -7173 61543
rect -7207 61441 -7173 61475
rect -7207 61373 -7173 61407
rect -7207 61305 -7173 61339
rect -7207 61237 -7173 61271
rect -7207 61169 -7173 61203
rect -7207 61101 -7173 61135
rect -7207 61033 -7173 61067
rect -7207 60965 -7173 60999
rect -7207 60897 -7173 60931
rect -7207 60829 -7173 60863
rect -7207 60761 -7173 60795
rect -7207 60693 -7173 60727
rect -7207 60625 -7173 60659
rect -7207 60557 -7173 60591
rect -7207 60489 -7173 60523
rect -7207 60421 -7173 60455
rect -7207 60353 -7173 60387
rect -7207 60285 -7173 60319
rect -7207 60217 -7173 60251
rect -7207 60149 -7173 60183
rect -7207 60081 -7173 60115
rect -7207 60013 -7173 60047
rect -7207 59945 -7173 59979
rect -7207 59877 -7173 59911
rect -7207 59809 -7173 59843
rect -7207 59741 -7173 59775
rect -7207 59673 -7173 59707
rect -7207 59605 -7173 59639
rect -7207 59537 -7173 59571
rect -7207 59469 -7173 59503
rect -7207 59401 -7173 59435
rect -7207 59333 -7173 59367
rect -7207 59265 -7173 59299
rect -7207 59197 -7173 59231
rect -7207 59129 -7173 59163
rect -7207 59061 -7173 59095
rect -7207 58993 -7173 59027
rect -7207 58925 -7173 58959
rect -7207 58857 -7173 58891
rect -7207 58789 -7173 58823
rect -7207 58721 -7173 58755
rect -7207 58653 -7173 58687
rect -7207 58585 -7173 58619
rect -7207 58517 -7173 58551
rect -7207 58449 -7173 58483
rect -7207 58381 -7173 58415
rect -7207 58313 -7173 58347
rect -7207 58245 -7173 58279
rect -7207 58177 -7173 58211
rect -7207 58109 -7173 58143
rect -7207 58041 -7173 58075
rect -7207 57973 -7173 58007
rect -7207 57905 -7173 57939
rect -7207 57837 -7173 57871
rect -7207 57769 -7173 57803
rect -7207 57701 -7173 57735
rect -7207 57633 -7173 57667
rect -7207 57565 -7173 57599
rect -7207 57497 -7173 57531
rect -7207 57429 -7173 57463
rect -7207 57361 -7173 57395
rect -7207 57293 -7173 57327
rect -7207 57225 -7173 57259
rect -7207 57157 -7173 57191
rect -7207 57089 -7173 57123
rect -7207 57021 -7173 57055
rect -7207 56953 -7173 56987
rect -7207 56885 -7173 56919
rect -7207 56817 -7173 56851
rect -7207 56749 -7173 56783
rect -7207 56681 -7173 56715
rect -7207 56613 -7173 56647
rect -7207 56545 -7173 56579
rect -7207 56477 -7173 56511
rect -7207 56409 -7173 56443
rect -7207 56341 -7173 56375
rect -10614 56270 -10580 56304
rect -10546 56270 -10512 56304
rect -10478 56270 -10444 56304
rect -10410 56270 -10376 56304
rect -10342 56270 -10308 56304
rect -10274 56270 -10240 56304
rect -10206 56270 -10172 56304
rect -10138 56270 -10104 56304
rect -10070 56270 -10036 56304
rect -10002 56270 -9968 56304
rect -9934 56270 -9900 56304
rect -9866 56270 -9832 56304
rect -9798 56270 -9764 56304
rect -9730 56270 -9696 56304
rect -9662 56270 -9628 56304
rect -9594 56270 -9560 56304
rect -9526 56270 -9492 56304
rect -9458 56270 -9424 56304
rect -9390 56270 -9356 56304
rect -9322 56270 -9288 56304
rect -9254 56270 -9220 56304
rect -9186 56270 -9152 56304
rect -9118 56270 -9084 56304
rect -9050 56270 -9016 56304
rect -8982 56270 -8948 56304
rect -8914 56270 -8880 56304
rect -8846 56270 -8812 56304
rect -8778 56270 -8744 56304
rect -8710 56270 -8676 56304
rect -8642 56270 -8608 56304
rect -8574 56270 -8540 56304
rect -8506 56270 -8472 56304
rect -8438 56270 -8404 56304
rect -8370 56270 -8336 56304
rect -8302 56270 -8268 56304
rect -8234 56270 -8200 56304
rect -8166 56270 -8132 56304
rect -8098 56270 -8064 56304
rect -8030 56270 -7996 56304
rect -7962 56270 -7928 56304
rect -7894 56270 -7860 56304
rect -7826 56270 -7792 56304
rect -7758 56270 -7724 56304
rect -7690 56270 -7656 56304
rect -7622 56270 -7588 56304
rect -7554 56270 -7520 56304
rect -7486 56270 -7452 56304
rect -7418 56270 -7384 56304
rect -7350 56270 -7316 56304
rect -7282 56270 -7248 56304
rect -3718 64122 -3684 64156
rect -3718 64054 -3684 64088
rect -3718 63986 -3684 64020
rect -3718 63918 -3684 63952
rect -3718 63850 -3684 63884
rect -3718 63782 -3684 63816
rect -3718 63714 -3684 63748
rect -3718 63646 -3684 63680
rect -3718 63578 -3684 63612
rect -3718 63510 -3684 63544
rect -3718 63442 -3684 63476
rect -3718 63374 -3684 63408
rect -3718 63306 -3684 63340
rect -3718 63238 -3684 63272
rect -3718 63170 -3684 63204
rect -3718 63102 -3684 63136
rect -3718 63034 -3684 63068
rect -3718 62966 -3684 63000
rect -3718 62898 -3684 62932
rect -3718 62830 -3684 62864
rect -3718 62762 -3684 62796
rect -3718 62694 -3684 62728
rect -3718 62626 -3684 62660
rect -3718 62558 -3684 62592
rect -3718 62490 -3684 62524
rect -3718 62422 -3684 62456
rect -3718 62354 -3684 62388
rect -3718 62286 -3684 62320
rect -3718 62218 -3684 62252
rect -3718 62150 -3684 62184
rect -3718 62082 -3684 62116
rect 59191 74772 59225 74806
rect 59259 74772 59293 74806
rect 59327 74772 59361 74806
rect 59395 74772 59429 74806
rect 59463 74772 59497 74806
rect 59531 74772 59565 74806
rect 59599 74772 59633 74806
rect 59667 74772 59701 74806
rect 59735 74772 59769 74806
rect 59803 74772 59837 74806
rect 59871 74772 59905 74806
rect 59939 74772 59973 74806
rect 60007 74772 60041 74806
rect 60075 74772 60109 74806
rect 60143 74772 60177 74806
rect 60211 74772 60245 74806
rect 60279 74772 60313 74806
rect 60347 74772 60381 74806
rect 60415 74772 60449 74806
rect 60483 74772 60517 74806
rect 60551 74772 60585 74806
rect 60619 74772 60653 74806
rect 60687 74772 60721 74806
rect 60755 74772 60789 74806
rect 60823 74772 60857 74806
rect 60891 74772 60925 74806
rect 60959 74772 60993 74806
rect 61027 74772 61061 74806
rect 61095 74772 61129 74806
rect 61163 74772 61197 74806
rect 61231 74772 61265 74806
rect 61299 74772 61333 74806
rect 61367 74772 61401 74806
rect 61435 74772 61469 74806
rect 61503 74772 61537 74806
rect 61571 74772 61605 74806
rect 61639 74772 61673 74806
rect 61707 74772 61741 74806
rect 61775 74772 61809 74806
rect 61843 74772 61877 74806
rect 61911 74772 61945 74806
rect 61979 74772 62013 74806
rect 62047 74772 62081 74806
rect 62115 74772 62149 74806
rect 62183 74772 62217 74806
rect 62251 74772 62285 74806
rect 62319 74772 62353 74806
rect 62387 74772 62421 74806
rect 62455 74772 62489 74806
rect 62523 74772 62557 74806
rect 62591 74772 62625 74806
rect 62659 74772 62693 74806
rect 62727 74772 62761 74806
rect 62795 74772 62829 74806
rect 62863 74772 62897 74806
rect 62931 74772 62965 74806
rect 62999 74772 63033 74806
rect 63067 74772 63101 74806
rect 63135 74772 63169 74806
rect 63203 74772 63237 74806
rect 63271 74772 63305 74806
rect 63339 74772 63373 74806
rect 63407 74772 63441 74806
rect 63475 74772 63509 74806
rect 63543 74772 63577 74806
rect 63611 74772 63645 74806
rect 63679 74772 63713 74806
rect 63747 74772 63781 74806
rect 63815 74772 63849 74806
rect 63883 74772 63917 74806
rect 63951 74772 63985 74806
rect 64019 74772 64053 74806
rect 64087 74772 64121 74806
rect 64155 74772 64189 74806
rect 64223 74772 64257 74806
rect 64291 74772 64325 74806
rect 64359 74772 64393 74806
rect 64427 74772 64461 74806
rect 64495 74772 64529 74806
rect 64563 74772 64597 74806
rect 64631 74772 64665 74806
rect 64699 74772 64733 74806
rect 64767 74772 64801 74806
rect 64835 74772 64869 74806
rect 64903 74772 64937 74806
rect 64971 74772 65005 74806
rect 65039 74772 65073 74806
rect 65107 74772 65141 74806
rect 65175 74772 65209 74806
rect 65243 74772 65277 74806
rect 65311 74772 65345 74806
rect 65379 74772 65413 74806
rect 65447 74772 65481 74806
rect 65515 74772 65549 74806
rect 65583 74772 65617 74806
rect 65651 74772 65685 74806
rect 65719 74772 65753 74806
rect 65787 74772 65821 74806
rect 65855 74772 65889 74806
rect 65923 74772 65957 74806
rect 65991 74772 66025 74806
rect 66059 74772 66093 74806
rect 66127 74772 66161 74806
rect 66195 74772 66229 74806
rect 66263 74772 66297 74806
rect 66331 74772 66365 74806
rect 66399 74772 66433 74806
rect 66467 74772 66501 74806
rect 66535 74772 66569 74806
rect 66603 74772 66637 74806
rect 66671 74772 66705 74806
rect 66739 74772 66773 74806
rect 66807 74772 66841 74806
rect 66875 74772 66909 74806
rect 66943 74772 66977 74806
rect 67011 74772 67045 74806
rect 67079 74772 67113 74806
rect 67147 74772 67181 74806
rect 67215 74772 67249 74806
rect 67283 74772 67317 74806
rect 67351 74772 67385 74806
rect 67419 74772 67453 74806
rect 67487 74772 67521 74806
rect 67555 74772 67589 74806
rect 67623 74772 67657 74806
rect 67691 74772 67725 74806
rect 67759 74772 67793 74806
rect 67827 74772 67861 74806
rect 67895 74772 67929 74806
rect 67963 74772 67997 74806
rect 68031 74772 68065 74806
rect 68099 74772 68133 74806
rect 68167 74772 68201 74806
rect 68235 74772 68269 74806
rect 68303 74772 68337 74806
rect 68371 74772 68405 74806
rect 68439 74772 68473 74806
rect 68507 74772 68541 74806
rect 68575 74772 68609 74806
rect 68643 74772 68677 74806
rect 68711 74772 68745 74806
rect 68779 74772 68813 74806
rect 68847 74772 68881 74806
rect 68915 74772 68949 74806
rect 68983 74772 69017 74806
rect 69051 74772 69085 74806
rect 69119 74772 69153 74806
rect 69187 74772 69221 74806
rect 69255 74772 69289 74806
rect 69323 74772 69357 74806
rect 69391 74772 69425 74806
rect 69459 74772 69493 74806
rect 69527 74772 69561 74806
rect 69595 74772 69629 74806
rect 69663 74772 69697 74806
rect 69731 74772 69765 74806
rect 69799 74772 69833 74806
rect 69867 74772 69901 74806
rect 69935 74772 69969 74806
rect 70003 74772 70037 74806
rect 70071 74772 70105 74806
rect 70139 74772 70173 74806
rect 70207 74772 70241 74806
rect 70275 74772 70309 74806
rect 70343 74772 70377 74806
rect 70411 74772 70445 74806
rect 70479 74772 70513 74806
rect 70547 74772 70581 74806
rect 70615 74772 70649 74806
rect 70683 74772 70717 74806
rect 70751 74772 70785 74806
rect 59104 74711 59138 74745
rect 59104 74643 59138 74677
rect 59104 74575 59138 74609
rect 59104 74507 59138 74541
rect 59104 74439 59138 74473
rect 59104 74371 59138 74405
rect 59104 74303 59138 74337
rect 59104 74235 59138 74269
rect 59104 74167 59138 74201
rect 59104 74099 59138 74133
rect 59104 74031 59138 74065
rect 59104 73963 59138 73997
rect 59104 73895 59138 73929
rect 59104 73827 59138 73861
rect 59104 73759 59138 73793
rect 59104 73691 59138 73725
rect 59104 73623 59138 73657
rect 59104 73555 59138 73589
rect 59104 73487 59138 73521
rect 59104 73419 59138 73453
rect 59104 73351 59138 73385
rect 59104 73283 59138 73317
rect 59104 73215 59138 73249
rect 59104 73147 59138 73181
rect 59104 73079 59138 73113
rect 59104 73011 59138 73045
rect 59104 72943 59138 72977
rect 59104 72875 59138 72909
rect 59104 72807 59138 72841
rect 59104 72739 59138 72773
rect 59104 72671 59138 72705
rect 59104 72603 59138 72637
rect 59104 72535 59138 72569
rect 59104 72467 59138 72501
rect 59104 72399 59138 72433
rect 59104 72331 59138 72365
rect 59104 72263 59138 72297
rect 59104 72195 59138 72229
rect 59104 72127 59138 72161
rect 59104 72059 59138 72093
rect 59104 71991 59138 72025
rect 59104 71923 59138 71957
rect 59104 71855 59138 71889
rect 59104 71787 59138 71821
rect 59104 71719 59138 71753
rect 59104 71651 59138 71685
rect 59104 71583 59138 71617
rect 59104 71515 59138 71549
rect 59104 71447 59138 71481
rect 59104 71379 59138 71413
rect 59104 71311 59138 71345
rect 59104 71243 59138 71277
rect 59104 71175 59138 71209
rect 59104 71107 59138 71141
rect 59104 71039 59138 71073
rect 59104 70971 59138 71005
rect 59104 70903 59138 70937
rect 59104 70835 59138 70869
rect 59104 70767 59138 70801
rect 59104 70699 59138 70733
rect 59104 70631 59138 70665
rect 59104 70563 59138 70597
rect 59104 70495 59138 70529
rect 59104 70427 59138 70461
rect 59104 70359 59138 70393
rect 59104 70291 59138 70325
rect 59104 70223 59138 70257
rect 59104 70155 59138 70189
rect 59104 70087 59138 70121
rect 59104 70019 59138 70053
rect 59104 69951 59138 69985
rect 59104 69883 59138 69917
rect 59104 69815 59138 69849
rect 59104 69747 59138 69781
rect 59104 69679 59138 69713
rect 59104 69611 59138 69645
rect 59104 69543 59138 69577
rect 59104 69475 59138 69509
rect 59104 69407 59138 69441
rect 59104 69339 59138 69373
rect 59104 69271 59138 69305
rect 59104 69203 59138 69237
rect 59104 69135 59138 69169
rect 59104 69067 59138 69101
rect 59104 68999 59138 69033
rect 59104 68931 59138 68965
rect 59104 68863 59138 68897
rect 59104 68795 59138 68829
rect 59104 68727 59138 68761
rect 59104 68659 59138 68693
rect 59104 68591 59138 68625
rect 59104 68523 59138 68557
rect 59104 68455 59138 68489
rect 59104 68387 59138 68421
rect 59104 68319 59138 68353
rect 59104 68251 59138 68285
rect 59104 68183 59138 68217
rect 59104 68115 59138 68149
rect 59104 68047 59138 68081
rect 59104 67979 59138 68013
rect 59104 67911 59138 67945
rect 59104 67843 59138 67877
rect 59104 67775 59138 67809
rect 59104 67707 59138 67741
rect 59104 67639 59138 67673
rect 59104 67571 59138 67605
rect 59104 67503 59138 67537
rect 59104 67435 59138 67469
rect 59104 67367 59138 67401
rect 59104 67299 59138 67333
rect 59104 67231 59138 67265
rect 59104 67163 59138 67197
rect 59104 67095 59138 67129
rect 59104 67027 59138 67061
rect 59104 66959 59138 66993
rect 59104 66891 59138 66925
rect 59104 66823 59138 66857
rect 59104 66755 59138 66789
rect 59104 66687 59138 66721
rect 59104 66619 59138 66653
rect 59104 66551 59138 66585
rect 59104 66483 59138 66517
rect 59104 66415 59138 66449
rect 59104 66347 59138 66381
rect 59104 66279 59138 66313
rect 59104 66211 59138 66245
rect 59104 66143 59138 66177
rect 59104 66075 59138 66109
rect 59104 66007 59138 66041
rect 59104 65939 59138 65973
rect 59104 65871 59138 65905
rect 59104 65803 59138 65837
rect 59104 65735 59138 65769
rect 59104 65667 59138 65701
rect 59104 65599 59138 65633
rect 59104 65531 59138 65565
rect 59104 65463 59138 65497
rect 59104 65395 59138 65429
rect 59104 65327 59138 65361
rect 59104 65259 59138 65293
rect 59104 65191 59138 65225
rect 59104 65123 59138 65157
rect 59104 65055 59138 65089
rect 59104 64987 59138 65021
rect 59104 64919 59138 64953
rect 59104 64851 59138 64885
rect 59104 64783 59138 64817
rect 59104 64715 59138 64749
rect 59104 64647 59138 64681
rect 59104 64579 59138 64613
rect 59104 64511 59138 64545
rect 59104 64443 59138 64477
rect 59104 64375 59138 64409
rect 59104 64307 59138 64341
rect 59104 64239 59138 64273
rect 59104 64171 59138 64205
rect 59104 64103 59138 64137
rect 59104 64035 59138 64069
rect 59104 63967 59138 64001
rect 59104 63899 59138 63933
rect 59104 63831 59138 63865
rect 59104 63763 59138 63797
rect 59104 63695 59138 63729
rect 59104 63627 59138 63661
rect 59104 63559 59138 63593
rect 59104 63491 59138 63525
rect 59104 63423 59138 63457
rect 59104 63355 59138 63389
rect 59104 63287 59138 63321
rect 59104 63219 59138 63253
rect 59104 63151 59138 63185
rect 59104 63083 59138 63117
rect 59104 63015 59138 63049
rect 59104 62947 59138 62981
rect 59104 62879 59138 62913
rect 59104 62811 59138 62845
rect 59104 62743 59138 62777
rect 59104 62675 59138 62709
rect 59104 62607 59138 62641
rect 59104 62539 59138 62573
rect 59104 62471 59138 62505
rect 59104 62403 59138 62437
rect 59104 62335 59138 62369
rect 59104 62267 59138 62301
rect 59104 62199 59138 62233
rect 59104 62131 59138 62165
rect 59104 62063 59138 62097
rect -3718 62014 -3684 62048
rect -3718 61946 -3684 61980
rect -3718 61878 -3684 61912
rect -3718 61810 -3684 61844
rect -3718 61742 -3684 61776
rect -3718 61674 -3684 61708
rect -3718 61606 -3684 61640
rect -3718 61538 -3684 61572
rect -3718 61470 -3684 61504
rect -3718 61402 -3684 61436
rect -3718 61334 -3684 61368
rect -3718 61266 -3684 61300
rect -3718 61198 -3684 61232
rect -3718 61130 -3684 61164
rect -3718 61062 -3684 61096
rect -3718 60994 -3684 61028
rect -3718 60926 -3684 60960
rect -3718 60858 -3684 60892
rect -3718 60790 -3684 60824
rect -3718 60722 -3684 60756
rect -3718 60654 -3684 60688
rect -3718 60586 -3684 60620
rect -3718 60518 -3684 60552
rect -3718 60450 -3684 60484
rect -3718 60382 -3684 60416
rect -3718 60314 -3684 60348
rect -3718 60246 -3684 60280
rect -3718 60178 -3684 60212
rect -3718 60110 -3684 60144
rect -3718 60042 -3684 60076
rect -3718 59974 -3684 60008
rect -3718 59906 -3684 59940
rect -3718 59838 -3684 59872
rect -3718 59770 -3684 59804
rect -3718 59702 -3684 59736
rect -3718 59634 -3684 59668
rect -3718 59566 -3684 59600
rect -3718 59498 -3684 59532
rect -3718 59430 -3684 59464
rect -3718 59362 -3684 59396
rect -3718 59294 -3684 59328
rect -3718 59226 -3684 59260
rect -3718 59158 -3684 59192
rect -3718 59090 -3684 59124
rect -3718 59022 -3684 59056
rect -3718 58954 -3684 58988
rect -3718 58886 -3684 58920
rect -3718 58818 -3684 58852
rect -3718 58750 -3684 58784
rect -3718 58682 -3684 58716
rect -3718 58614 -3684 58648
rect -3718 58546 -3684 58580
rect -3718 58478 -3684 58512
rect -3718 58410 -3684 58444
rect -3718 58342 -3684 58376
rect 50530 62006 50564 62040
rect 50598 62006 50632 62040
rect 50666 62006 50700 62040
rect 50734 62006 50768 62040
rect 50802 62006 50836 62040
rect 50870 62006 50904 62040
rect 50938 62006 50972 62040
rect 51006 62006 51040 62040
rect 51074 62006 51108 62040
rect 51142 62006 51176 62040
rect 51210 62006 51244 62040
rect 51278 62006 51312 62040
rect 51346 62006 51380 62040
rect 51414 62006 51448 62040
rect 51482 62006 51516 62040
rect 51550 62006 51584 62040
rect 51618 62006 51652 62040
rect 51686 62006 51720 62040
rect 51754 62006 51788 62040
rect 51822 62006 51856 62040
rect 51890 62006 51924 62040
rect 51958 62006 51992 62040
rect 52026 62006 52060 62040
rect 52094 62006 52128 62040
rect 52162 62006 52196 62040
rect 52230 62006 52264 62040
rect 52298 62006 52332 62040
rect 52366 62006 52400 62040
rect 52434 62006 52468 62040
rect 52502 62006 52536 62040
rect 52570 62006 52604 62040
rect 52638 62006 52672 62040
rect 52706 62006 52740 62040
rect 52774 62006 52808 62040
rect 52842 62006 52876 62040
rect 52910 62006 52944 62040
rect 52978 62006 53012 62040
rect 53046 62006 53080 62040
rect 53114 62006 53148 62040
rect 53182 62006 53216 62040
rect 53250 62006 53284 62040
rect 53318 62006 53352 62040
rect 53386 62006 53420 62040
rect 53454 62006 53488 62040
rect 53522 62006 53556 62040
rect 53590 62006 53624 62040
rect 53658 62006 53692 62040
rect 53726 62006 53760 62040
rect 53794 62006 53828 62040
rect 53862 62006 53896 62040
rect 53930 62006 53964 62040
rect 53998 62006 54032 62040
rect 54066 62006 54100 62040
rect 54134 62006 54168 62040
rect 54202 62006 54236 62040
rect 54270 62006 54304 62040
rect 54338 62006 54372 62040
rect 54406 62006 54440 62040
rect 54474 62006 54508 62040
rect 54542 62006 54576 62040
rect 54610 62006 54644 62040
rect 54678 62006 54712 62040
rect 54746 62006 54780 62040
rect 54814 62006 54848 62040
rect 54882 62006 54916 62040
rect 54950 62006 54984 62040
rect 55018 62006 55052 62040
rect 55086 62006 55120 62040
rect 55154 62006 55188 62040
rect 55222 62006 55256 62040
rect 55290 62006 55324 62040
rect 55358 62006 55392 62040
rect 55426 62006 55460 62040
rect 55494 62006 55528 62040
rect 55562 62006 55596 62040
rect 55630 62006 55664 62040
rect 55698 62006 55732 62040
rect 55766 62006 55800 62040
rect 55834 62006 55868 62040
rect 55902 62006 55936 62040
rect 55970 62006 56004 62040
rect 56038 62006 56072 62040
rect 56106 62006 56140 62040
rect 56174 62006 56208 62040
rect 56242 62006 56276 62040
rect 50456 61942 50490 61976
rect 50456 61874 50490 61908
rect 50456 61806 50490 61840
rect 50456 61738 50490 61772
rect 50456 61670 50490 61704
rect 50456 61602 50490 61636
rect 50456 61534 50490 61568
rect 50456 61466 50490 61500
rect 50456 61398 50490 61432
rect 50456 61330 50490 61364
rect 50456 61262 50490 61296
rect 50456 61194 50490 61228
rect 50456 61126 50490 61160
rect 50456 61058 50490 61092
rect 50456 60990 50490 61024
rect 50456 60922 50490 60956
rect 50456 60854 50490 60888
rect 50456 60786 50490 60820
rect 50456 60718 50490 60752
rect 50456 60650 50490 60684
rect 50456 60582 50490 60616
rect 50456 60514 50490 60548
rect 50456 60446 50490 60480
rect 50456 60378 50490 60412
rect 50456 60310 50490 60344
rect 50456 60242 50490 60276
rect 50456 60174 50490 60208
rect 50456 60106 50490 60140
rect 50456 60038 50490 60072
rect 50456 59970 50490 60004
rect 50456 59902 50490 59936
rect 50456 59834 50490 59868
rect 50456 59766 50490 59800
rect 50456 59698 50490 59732
rect 50456 59630 50490 59664
rect 50456 59562 50490 59596
rect 50456 59494 50490 59528
rect 50456 59426 50490 59460
rect 50456 59358 50490 59392
rect 50456 59290 50490 59324
rect 50456 59222 50490 59256
rect 50456 59154 50490 59188
rect 50456 59086 50490 59120
rect 50456 59018 50490 59052
rect 50456 58950 50490 58984
rect 50456 58882 50490 58916
rect 50456 58814 50490 58848
rect 50456 58746 50490 58780
rect 50456 58678 50490 58712
rect 50456 58610 50490 58644
rect 50456 58542 50490 58576
rect 50456 58474 50490 58508
rect 50456 58406 50490 58440
rect 56316 61942 56350 61976
rect 56316 61874 56350 61908
rect 56316 61806 56350 61840
rect 56316 61738 56350 61772
rect 56316 61670 56350 61704
rect 56316 61602 56350 61636
rect 56316 61534 56350 61568
rect 56316 61466 56350 61500
rect 56316 61398 56350 61432
rect 56316 61330 56350 61364
rect 56316 61262 56350 61296
rect 56316 61194 56350 61228
rect 56316 61126 56350 61160
rect 56316 61058 56350 61092
rect 56316 60990 56350 61024
rect 56316 60922 56350 60956
rect 56316 60854 56350 60888
rect 56316 60786 56350 60820
rect 56316 60718 56350 60752
rect 56316 60650 56350 60684
rect 56316 60582 56350 60616
rect 56316 60514 56350 60548
rect 56316 60446 56350 60480
rect 56316 60378 56350 60412
rect 56316 60310 56350 60344
rect 56316 60242 56350 60276
rect 56316 60174 56350 60208
rect 56316 60106 56350 60140
rect 56316 60038 56350 60072
rect 56316 59970 56350 60004
rect 56316 59902 56350 59936
rect 56316 59834 56350 59868
rect 56316 59766 56350 59800
rect 56316 59698 56350 59732
rect 56316 59630 56350 59664
rect 56316 59562 56350 59596
rect 56316 59494 56350 59528
rect 56316 59426 56350 59460
rect 56316 59358 56350 59392
rect 56316 59290 56350 59324
rect 56316 59222 56350 59256
rect 56316 59154 56350 59188
rect 56316 59086 56350 59120
rect 56316 59018 56350 59052
rect 56316 58950 56350 58984
rect 56316 58882 56350 58916
rect 56316 58814 56350 58848
rect 56316 58746 56350 58780
rect 56316 58678 56350 58712
rect 56316 58610 56350 58644
rect 56316 58542 56350 58576
rect 56316 58474 56350 58508
rect 56316 58406 56350 58440
rect 50530 58342 50564 58376
rect 50598 58342 50632 58376
rect 50666 58342 50700 58376
rect 50734 58342 50768 58376
rect 50802 58342 50836 58376
rect 50870 58342 50904 58376
rect 50938 58342 50972 58376
rect 51006 58342 51040 58376
rect 51074 58342 51108 58376
rect 51142 58342 51176 58376
rect 51210 58342 51244 58376
rect 51278 58342 51312 58376
rect 51346 58342 51380 58376
rect 51414 58342 51448 58376
rect 51482 58342 51516 58376
rect 51550 58342 51584 58376
rect 51618 58342 51652 58376
rect 51686 58342 51720 58376
rect 51754 58342 51788 58376
rect 51822 58342 51856 58376
rect 51890 58342 51924 58376
rect 51958 58342 51992 58376
rect 52026 58342 52060 58376
rect 52094 58342 52128 58376
rect 52162 58342 52196 58376
rect 52230 58342 52264 58376
rect 52298 58342 52332 58376
rect 52366 58342 52400 58376
rect 52434 58342 52468 58376
rect 52502 58342 52536 58376
rect 52570 58342 52604 58376
rect 52638 58342 52672 58376
rect 52706 58342 52740 58376
rect 52774 58342 52808 58376
rect 52842 58342 52876 58376
rect 52910 58342 52944 58376
rect 52978 58342 53012 58376
rect 53046 58342 53080 58376
rect 53114 58342 53148 58376
rect 53182 58342 53216 58376
rect 53250 58342 53284 58376
rect 53318 58342 53352 58376
rect 53386 58342 53420 58376
rect 53454 58342 53488 58376
rect 53522 58342 53556 58376
rect 53590 58342 53624 58376
rect 53658 58342 53692 58376
rect 53726 58342 53760 58376
rect 53794 58342 53828 58376
rect 53862 58342 53896 58376
rect 53930 58342 53964 58376
rect 53998 58342 54032 58376
rect 54066 58342 54100 58376
rect 54134 58342 54168 58376
rect 54202 58342 54236 58376
rect 54270 58342 54304 58376
rect 54338 58342 54372 58376
rect 54406 58342 54440 58376
rect 54474 58342 54508 58376
rect 54542 58342 54576 58376
rect 54610 58342 54644 58376
rect 54678 58342 54712 58376
rect 54746 58342 54780 58376
rect 54814 58342 54848 58376
rect 54882 58342 54916 58376
rect 54950 58342 54984 58376
rect 55018 58342 55052 58376
rect 55086 58342 55120 58376
rect 55154 58342 55188 58376
rect 55222 58342 55256 58376
rect 55290 58342 55324 58376
rect 55358 58342 55392 58376
rect 55426 58342 55460 58376
rect 55494 58342 55528 58376
rect 55562 58342 55596 58376
rect 55630 58342 55664 58376
rect 55698 58342 55732 58376
rect 55766 58342 55800 58376
rect 55834 58342 55868 58376
rect 55902 58342 55936 58376
rect 55970 58342 56004 58376
rect 56038 58342 56072 58376
rect 56106 58342 56140 58376
rect 56174 58342 56208 58376
rect 56242 58342 56276 58376
rect 59104 61995 59138 62029
rect 59104 61927 59138 61961
rect 59104 61859 59138 61893
rect 59104 61791 59138 61825
rect 59104 61723 59138 61757
rect 59104 61655 59138 61689
rect 59104 61587 59138 61621
rect 59104 61519 59138 61553
rect 59104 61451 59138 61485
rect 59104 61383 59138 61417
rect 59104 61315 59138 61349
rect 59104 61247 59138 61281
rect 59104 61179 59138 61213
rect 59104 61111 59138 61145
rect 59104 61043 59138 61077
rect 59104 60975 59138 61009
rect 59104 60907 59138 60941
rect 59104 60839 59138 60873
rect 59104 60771 59138 60805
rect 59104 60703 59138 60737
rect 59104 60635 59138 60669
rect 59104 60567 59138 60601
rect 59104 60499 59138 60533
rect 59104 60431 59138 60465
rect 59104 60363 59138 60397
rect 59104 60295 59138 60329
rect 59104 60227 59138 60261
rect 59104 60159 59138 60193
rect 59104 60091 59138 60125
rect 59104 60023 59138 60057
rect 59104 59955 59138 59989
rect 59104 59887 59138 59921
rect 59104 59819 59138 59853
rect 59104 59751 59138 59785
rect 59104 59683 59138 59717
rect 59104 59615 59138 59649
rect 59104 59547 59138 59581
rect 59104 59479 59138 59513
rect 59104 59411 59138 59445
rect 59104 59343 59138 59377
rect 59104 59275 59138 59309
rect 59104 59207 59138 59241
rect 59104 59139 59138 59173
rect 59104 59071 59138 59105
rect 59104 59003 59138 59037
rect 59104 58935 59138 58969
rect 59104 58867 59138 58901
rect 59104 58799 59138 58833
rect 59104 58731 59138 58765
rect 59104 58663 59138 58697
rect 59104 58595 59138 58629
rect 59104 58527 59138 58561
rect 59104 58459 59138 58493
rect 59104 58391 59138 58425
rect 59104 58323 59138 58357
rect -3718 58274 -3684 58308
rect -3718 58206 -3684 58240
rect -3718 58138 -3684 58172
rect -3718 58070 -3684 58104
rect -3718 58002 -3684 58036
rect -3718 57934 -3684 57968
rect -3718 57866 -3684 57900
rect -3718 57798 -3684 57832
rect -3718 57730 -3684 57764
rect -3718 57662 -3684 57696
rect -3718 57594 -3684 57628
rect -3718 57526 -3684 57560
rect -3718 57458 -3684 57492
rect -3718 57390 -3684 57424
rect -3718 57322 -3684 57356
rect -3718 57254 -3684 57288
rect -3718 57186 -3684 57220
rect -3718 57118 -3684 57152
rect -3718 57050 -3684 57084
rect -3718 56982 -3684 57016
rect -3718 56914 -3684 56948
rect -3718 56846 -3684 56880
rect -3718 56778 -3684 56812
rect -3718 56710 -3684 56744
rect -3718 56642 -3684 56676
rect -3718 56574 -3684 56608
rect -3718 56506 -3684 56540
rect -3718 56438 -3684 56472
rect -3718 56370 -3684 56404
rect -3718 56302 -3684 56336
rect -10699 56211 -10665 56245
rect -10699 56143 -10665 56177
rect -10699 56075 -10665 56109
rect -10699 56007 -10665 56041
rect -10699 55939 -10665 55973
rect -10699 55871 -10665 55905
rect -10699 55803 -10665 55837
rect -10699 55735 -10665 55769
rect -10699 55667 -10665 55701
rect -10699 55599 -10665 55633
rect -10699 55531 -10665 55565
rect -10699 55463 -10665 55497
rect -10699 55395 -10665 55429
rect -10699 55327 -10665 55361
rect -10699 55259 -10665 55293
rect -10699 55191 -10665 55225
rect -10699 55123 -10665 55157
rect -10699 55055 -10665 55089
rect -10699 54987 -10665 55021
rect -10699 54919 -10665 54953
rect -10699 54851 -10665 54885
rect -10699 54783 -10665 54817
rect -10699 54715 -10665 54749
rect -10699 54647 -10665 54681
rect -10699 54579 -10665 54613
rect -10699 54511 -10665 54545
rect -10699 54443 -10665 54477
rect -10699 54375 -10665 54409
rect -10699 54307 -10665 54341
rect -10699 54239 -10665 54273
rect -10699 54171 -10665 54205
rect -10699 54103 -10665 54137
rect -10699 54035 -10665 54069
rect -10699 53967 -10665 54001
rect -10699 53899 -10665 53933
rect -10699 53831 -10665 53865
rect -10699 53763 -10665 53797
rect -10699 53695 -10665 53729
rect -10699 53627 -10665 53661
rect -10699 53559 -10665 53593
rect -10699 53491 -10665 53525
rect -10699 53423 -10665 53457
rect -10699 53355 -10665 53389
rect -10699 53287 -10665 53321
rect -10699 53219 -10665 53253
rect -10699 53151 -10665 53185
rect -10699 53083 -10665 53117
rect -10699 53015 -10665 53049
rect -10699 52947 -10665 52981
rect -10699 52879 -10665 52913
rect -10699 52811 -10665 52845
rect -10699 52743 -10665 52777
rect -10699 52675 -10665 52709
rect -10699 52607 -10665 52641
rect -10699 52539 -10665 52573
rect -10699 52471 -10665 52505
rect -10699 52403 -10665 52437
rect -10699 52335 -10665 52369
rect -10699 52267 -10665 52301
rect -10699 52199 -10665 52233
rect -10699 52131 -10665 52165
rect -10699 52063 -10665 52097
rect -10699 51995 -10665 52029
rect -10699 51927 -10665 51961
rect -10699 51859 -10665 51893
rect -10699 51791 -10665 51825
rect -10699 51723 -10665 51757
rect -10699 51655 -10665 51689
rect -10699 51587 -10665 51621
rect -10699 51519 -10665 51553
rect -10699 51451 -10665 51485
rect -10699 51383 -10665 51417
rect -10699 51315 -10665 51349
rect -10699 51247 -10665 51281
rect -10699 51179 -10665 51213
rect -10699 51111 -10665 51145
rect -10699 51043 -10665 51077
rect -10699 50975 -10665 51009
rect -10699 50907 -10665 50941
rect -10699 50839 -10665 50873
rect -10699 50771 -10665 50805
rect -10699 50703 -10665 50737
rect -10699 50635 -10665 50669
rect -10699 50567 -10665 50601
rect -10699 50499 -10665 50533
rect -10699 50431 -10665 50465
rect -10699 50363 -10665 50397
rect -10699 50295 -10665 50329
rect -10699 50227 -10665 50261
rect -10699 50159 -10665 50193
rect -10699 50091 -10665 50125
rect -10699 50023 -10665 50057
rect -10699 49955 -10665 49989
rect -10699 49887 -10665 49921
rect -10699 49819 -10665 49853
rect -10699 49751 -10665 49785
rect -10699 49683 -10665 49717
rect -10699 49615 -10665 49649
rect -10699 49547 -10665 49581
rect -10699 49479 -10665 49513
rect -10699 49411 -10665 49445
rect -10699 49343 -10665 49377
rect -10699 49275 -10665 49309
rect -10699 49207 -10665 49241
rect -10699 49139 -10665 49173
rect -10699 49071 -10665 49105
rect -10699 49003 -10665 49037
rect -10699 48935 -10665 48969
rect -10699 48867 -10665 48901
rect -10699 48799 -10665 48833
rect -10699 48731 -10665 48765
rect -10699 48663 -10665 48697
rect -10699 48595 -10665 48629
rect -10699 48527 -10665 48561
rect -10699 48459 -10665 48493
rect -10699 48391 -10665 48425
rect -10699 48323 -10665 48357
rect -10699 48255 -10665 48289
rect -10699 48187 -10665 48221
rect -10699 48119 -10665 48153
rect -10699 48051 -10665 48085
rect -10699 47983 -10665 48017
rect -10699 47915 -10665 47949
rect -10699 47847 -10665 47881
rect -10699 47779 -10665 47813
rect -10699 47711 -10665 47745
rect -10699 47643 -10665 47677
rect -10699 47575 -10665 47609
rect -10699 47507 -10665 47541
rect -10699 47439 -10665 47473
rect -10699 47371 -10665 47405
rect -10699 47303 -10665 47337
rect -10699 47235 -10665 47269
rect -10699 47167 -10665 47201
rect -10699 47099 -10665 47133
rect -10699 47031 -10665 47065
rect -10699 46963 -10665 46997
rect -10699 46895 -10665 46929
rect -10699 46827 -10665 46861
rect -10699 46759 -10665 46793
rect -10699 46691 -10665 46725
rect -10699 46623 -10665 46657
rect -10699 46555 -10665 46589
rect -10699 46487 -10665 46521
rect -10699 46419 -10665 46453
rect -10699 46351 -10665 46385
rect -10699 46283 -10665 46317
rect -10699 46215 -10665 46249
rect -10699 46147 -10665 46181
rect -10699 46079 -10665 46113
rect -10699 46011 -10665 46045
rect -10699 45943 -10665 45977
rect -10699 45875 -10665 45909
rect -10699 45807 -10665 45841
rect -10699 45739 -10665 45773
rect -10699 45671 -10665 45705
rect -10699 45603 -10665 45637
rect -10699 45535 -10665 45569
rect -10699 45467 -10665 45501
rect -10699 45399 -10665 45433
rect -10699 45331 -10665 45365
rect -10699 45263 -10665 45297
rect -10699 45195 -10665 45229
rect -10699 45127 -10665 45161
rect -10699 45059 -10665 45093
rect -10699 44991 -10665 45025
rect -10699 44923 -10665 44957
rect -10699 44855 -10665 44889
rect -10699 44787 -10665 44821
rect -10699 44719 -10665 44753
rect -10699 44651 -10665 44685
rect -10699 44583 -10665 44617
rect -10699 44515 -10665 44549
rect -10699 44447 -10665 44481
rect -10699 44379 -10665 44413
rect -10699 44311 -10665 44345
rect -3718 56234 -3684 56268
rect -3718 56166 -3684 56200
rect -3718 56098 -3684 56132
rect -3718 56030 -3684 56064
rect -3718 55962 -3684 55996
rect -3718 55894 -3684 55928
rect -3718 55826 -3684 55860
rect -3718 55758 -3684 55792
rect -3718 55690 -3684 55724
rect -3718 55622 -3684 55656
rect -3718 55554 -3684 55588
rect -3718 55486 -3684 55520
rect -3718 55418 -3684 55452
rect -3718 55350 -3684 55384
rect -3718 55282 -3684 55316
rect -3718 55214 -3684 55248
rect -3718 55146 -3684 55180
rect -3718 55078 -3684 55112
rect -3718 55010 -3684 55044
rect -3718 54942 -3684 54976
rect -3718 54874 -3684 54908
rect -3718 54806 -3684 54840
rect -3718 54738 -3684 54772
rect -3718 54670 -3684 54704
rect -3718 54602 -3684 54636
rect -3718 54534 -3684 54568
rect -3718 54466 -3684 54500
rect -3718 54398 -3684 54432
rect -3718 54330 -3684 54364
rect -3718 54262 -3684 54296
rect -3718 54194 -3684 54228
rect -3718 54126 -3684 54160
rect -3718 54058 -3684 54092
rect -3718 53990 -3684 54024
rect -3718 53922 -3684 53956
rect -3718 53854 -3684 53888
rect -3718 53786 -3684 53820
rect -3718 53718 -3684 53752
rect -3718 53650 -3684 53684
rect -3718 53582 -3684 53616
rect -3718 53514 -3684 53548
rect -3718 53446 -3684 53480
rect -3718 53378 -3684 53412
rect -3718 53310 -3684 53344
rect -3718 53242 -3684 53276
rect -3718 53174 -3684 53208
rect -3718 53106 -3684 53140
rect -3718 53038 -3684 53072
rect -3718 52970 -3684 53004
rect -3718 52902 -3684 52936
rect -3718 52834 -3684 52868
rect -3718 52766 -3684 52800
rect -3718 52698 -3684 52732
rect -3718 52630 -3684 52664
rect -3718 52562 -3684 52596
rect -3718 52494 -3684 52528
rect -3718 52426 -3684 52460
rect -3718 52358 -3684 52392
rect -3718 52290 -3684 52324
rect -3718 52222 -3684 52256
rect -3718 52154 -3684 52188
rect -3718 52086 -3684 52120
rect -3718 52018 -3684 52052
rect -3718 51950 -3684 51984
rect -3718 51882 -3684 51916
rect -3718 51814 -3684 51848
rect -3718 51746 -3684 51780
rect -3718 51678 -3684 51712
rect -3718 51610 -3684 51644
rect -3718 51542 -3684 51576
rect -3718 51474 -3684 51508
rect -3718 51406 -3684 51440
rect -3718 51338 -3684 51372
rect -3718 51270 -3684 51304
rect -3718 51202 -3684 51236
rect -3718 51134 -3684 51168
rect -3718 51066 -3684 51100
rect -3718 50998 -3684 51032
rect -3718 50930 -3684 50964
rect -3718 50862 -3684 50896
rect -3718 50794 -3684 50828
rect -3718 50726 -3684 50760
rect -3718 50658 -3684 50692
rect -3718 50590 -3684 50624
rect -3718 50522 -3684 50556
rect -3718 50454 -3684 50488
rect -3718 50386 -3684 50420
rect -3718 50318 -3684 50352
rect -3718 50250 -3684 50284
rect -3718 50182 -3684 50216
rect -3718 50114 -3684 50148
rect -3718 50046 -3684 50080
rect -3718 49978 -3684 50012
rect -3718 49910 -3684 49944
rect -3718 49842 -3684 49876
rect -3718 49774 -3684 49808
rect -3718 49706 -3684 49740
rect -3718 49638 -3684 49672
rect -3718 49570 -3684 49604
rect -3718 49502 -3684 49536
rect -3718 49434 -3684 49468
rect -3718 49366 -3684 49400
rect -3718 49298 -3684 49332
rect -3718 49230 -3684 49264
rect -3718 49162 -3684 49196
rect -3718 49094 -3684 49128
rect -3718 49026 -3684 49060
rect -3718 48958 -3684 48992
rect -3718 48890 -3684 48924
rect -3718 48822 -3684 48856
rect -3718 48754 -3684 48788
rect -3718 48686 -3684 48720
rect -3718 48618 -3684 48652
rect -3718 48550 -3684 48584
rect -3718 48482 -3684 48516
rect -3718 48414 -3684 48448
rect -3718 48346 -3684 48380
rect -3718 48278 -3684 48312
rect -3718 48210 -3684 48244
rect -3718 48142 -3684 48176
rect -3718 48074 -3684 48108
rect -3718 48006 -3684 48040
rect -3718 47938 -3684 47972
rect -3718 47870 -3684 47904
rect -3718 47802 -3684 47836
rect -3718 47734 -3684 47768
rect -3718 47666 -3684 47700
rect -3718 47598 -3684 47632
rect -3718 47530 -3684 47564
rect -3718 47462 -3684 47496
rect -3718 47394 -3684 47428
rect -3718 47326 -3684 47360
rect -3718 47258 -3684 47292
rect -3718 47190 -3684 47224
rect -3718 47122 -3684 47156
rect -3718 47054 -3684 47088
rect -3718 46986 -3684 47020
rect -3718 46918 -3684 46952
rect -3718 46850 -3684 46884
rect -3718 46782 -3684 46816
rect -3718 46714 -3684 46748
rect -3718 46646 -3684 46680
rect -3718 46578 -3684 46612
rect -3718 46510 -3684 46544
rect -3718 46442 -3684 46476
rect -3718 46374 -3684 46408
rect -3718 46306 -3684 46340
rect -3718 46238 -3684 46272
rect -3718 46170 -3684 46204
rect -3718 46102 -3684 46136
rect -3718 46034 -3684 46068
rect -3718 45966 -3684 46000
rect -3718 45898 -3684 45932
rect 59104 58255 59138 58289
rect 59104 58187 59138 58221
rect 59104 58119 59138 58153
rect 59104 58051 59138 58085
rect 59104 57983 59138 58017
rect 59104 57915 59138 57949
rect 59104 57847 59138 57881
rect 59104 57779 59138 57813
rect 59104 57711 59138 57745
rect 59104 57643 59138 57677
rect 59104 57575 59138 57609
rect 59104 57507 59138 57541
rect 59104 57439 59138 57473
rect 59104 57371 59138 57405
rect 59104 57303 59138 57337
rect 59104 57235 59138 57269
rect 59104 57167 59138 57201
rect 59104 57099 59138 57133
rect 59104 57031 59138 57065
rect 59104 56963 59138 56997
rect 59104 56895 59138 56929
rect 59104 56827 59138 56861
rect 59104 56759 59138 56793
rect 59104 56691 59138 56725
rect 59104 56623 59138 56657
rect 59104 56555 59138 56589
rect 59104 56487 59138 56521
rect 59104 56419 59138 56453
rect 59104 56351 59138 56385
rect 59104 56283 59138 56317
rect 59104 56215 59138 56249
rect 59104 56147 59138 56181
rect 59104 56079 59138 56113
rect 59104 56011 59138 56045
rect 59104 55943 59138 55977
rect 59104 55875 59138 55909
rect 59104 55807 59138 55841
rect 59104 55739 59138 55773
rect 59104 55671 59138 55705
rect 59104 55603 59138 55637
rect 59104 55535 59138 55569
rect 59104 55467 59138 55501
rect 59104 55399 59138 55433
rect 59104 55331 59138 55365
rect 59104 55263 59138 55297
rect 59104 55195 59138 55229
rect 59104 55127 59138 55161
rect 59104 55059 59138 55093
rect 59104 54991 59138 55025
rect 59104 54923 59138 54957
rect 59104 54855 59138 54889
rect 59104 54787 59138 54821
rect 59104 54719 59138 54753
rect 59104 54651 59138 54685
rect 59104 54583 59138 54617
rect 59104 54515 59138 54549
rect 59104 54447 59138 54481
rect 59104 54379 59138 54413
rect 59104 54311 59138 54345
rect 59104 54243 59138 54277
rect 59104 54175 59138 54209
rect 59104 54107 59138 54141
rect 59104 54039 59138 54073
rect 59104 53971 59138 54005
rect 59104 53903 59138 53937
rect 59104 53835 59138 53869
rect 59104 53767 59138 53801
rect 59104 53699 59138 53733
rect 59104 53631 59138 53665
rect 59104 53563 59138 53597
rect 59104 53495 59138 53529
rect 59104 53427 59138 53461
rect 59104 53359 59138 53393
rect 59104 53291 59138 53325
rect 59104 53223 59138 53257
rect 59104 53155 59138 53189
rect 59104 53087 59138 53121
rect 59104 53019 59138 53053
rect 59104 52951 59138 52985
rect 59104 52883 59138 52917
rect 59104 52815 59138 52849
rect 59104 52747 59138 52781
rect 59104 52679 59138 52713
rect 59104 52611 59138 52645
rect 59104 52543 59138 52577
rect 59104 52475 59138 52509
rect 59104 52407 59138 52441
rect 59104 52339 59138 52373
rect 59104 52271 59138 52305
rect 59104 52203 59138 52237
rect 59104 52135 59138 52169
rect 59104 52067 59138 52101
rect 59104 51999 59138 52033
rect 59104 51931 59138 51965
rect 59104 51863 59138 51897
rect 59104 51795 59138 51829
rect 59104 51727 59138 51761
rect 59104 51659 59138 51693
rect 59104 51591 59138 51625
rect 59104 51523 59138 51557
rect 59104 51455 59138 51489
rect 59104 51387 59138 51421
rect 59104 51319 59138 51353
rect 59104 51251 59138 51285
rect 59104 51183 59138 51217
rect 59104 51115 59138 51149
rect 59104 51047 59138 51081
rect 59104 50979 59138 51013
rect 59104 50911 59138 50945
rect 59104 50843 59138 50877
rect 59104 50775 59138 50809
rect 59104 50707 59138 50741
rect 59104 50639 59138 50673
rect 59104 50571 59138 50605
rect 59104 50503 59138 50537
rect 59104 50435 59138 50469
rect 59104 50367 59138 50401
rect 59104 50299 59138 50333
rect 59104 50231 59138 50265
rect 59104 50163 59138 50197
rect 59104 50095 59138 50129
rect 59104 50027 59138 50061
rect 59104 49959 59138 49993
rect 59104 49891 59138 49925
rect 59104 49823 59138 49857
rect 59104 49755 59138 49789
rect 59104 49687 59138 49721
rect 59104 49619 59138 49653
rect 59104 49551 59138 49585
rect 59104 49483 59138 49517
rect 59104 49415 59138 49449
rect 59104 49347 59138 49381
rect 59104 49279 59138 49313
rect 59104 49211 59138 49245
rect 59104 49143 59138 49177
rect 59104 49075 59138 49109
rect 59104 49007 59138 49041
rect 59104 48939 59138 48973
rect 59104 48871 59138 48905
rect 59104 48803 59138 48837
rect 59104 48735 59138 48769
rect 59104 48667 59138 48701
rect 59104 48599 59138 48633
rect 59104 48531 59138 48565
rect 59104 48463 59138 48497
rect 59104 48395 59138 48429
rect 59104 48327 59138 48361
rect 59104 48259 59138 48293
rect 59104 48191 59138 48225
rect 59104 48123 59138 48157
rect 59104 48055 59138 48089
rect 59104 47987 59138 48021
rect 59104 47919 59138 47953
rect 59104 47851 59138 47885
rect 59104 47783 59138 47817
rect 59104 47715 59138 47749
rect 59104 47647 59138 47681
rect 59104 47579 59138 47613
rect 59104 47511 59138 47545
rect 59104 47443 59138 47477
rect 59104 47375 59138 47409
rect 59104 47307 59138 47341
rect 59104 47239 59138 47273
rect 59104 47171 59138 47205
rect 59104 47103 59138 47137
rect 59104 47035 59138 47069
rect 59104 46967 59138 47001
rect 59104 46899 59138 46933
rect 59104 46831 59138 46865
rect 59104 46763 59138 46797
rect 59104 46695 59138 46729
rect 59104 46627 59138 46661
rect 59104 46559 59138 46593
rect 59104 46491 59138 46525
rect 59104 46423 59138 46457
rect 59104 46355 59138 46389
rect 59104 46287 59138 46321
rect 59104 46219 59138 46253
rect 59104 46151 59138 46185
rect 59104 46083 59138 46117
rect 59104 46015 59138 46049
rect 59104 45947 59138 45981
rect 70838 74711 70872 74745
rect 70838 74643 70872 74677
rect 70838 74575 70872 74609
rect 70838 74507 70872 74541
rect 70838 74439 70872 74473
rect 70838 74371 70872 74405
rect 70838 74303 70872 74337
rect 70838 74235 70872 74269
rect 70838 74167 70872 74201
rect 70838 74099 70872 74133
rect 70838 74031 70872 74065
rect 70838 73963 70872 73997
rect 70838 73895 70872 73929
rect 70838 73827 70872 73861
rect 70838 73759 70872 73793
rect 70838 73691 70872 73725
rect 70838 73623 70872 73657
rect 70838 73555 70872 73589
rect 70838 73487 70872 73521
rect 70838 73419 70872 73453
rect 70838 73351 70872 73385
rect 70838 73283 70872 73317
rect 70838 73215 70872 73249
rect 70838 73147 70872 73181
rect 70838 73079 70872 73113
rect 70838 73011 70872 73045
rect 70838 72943 70872 72977
rect 70838 72875 70872 72909
rect 70838 72807 70872 72841
rect 70838 72739 70872 72773
rect 70838 72671 70872 72705
rect 70838 72603 70872 72637
rect 70838 72535 70872 72569
rect 70838 72467 70872 72501
rect 70838 72399 70872 72433
rect 70838 72331 70872 72365
rect 70838 72263 70872 72297
rect 70838 72195 70872 72229
rect 70838 72127 70872 72161
rect 70838 72059 70872 72093
rect 70838 71991 70872 72025
rect 70838 71923 70872 71957
rect 70838 71855 70872 71889
rect 70838 71787 70872 71821
rect 70838 71719 70872 71753
rect 70838 71651 70872 71685
rect 70838 71583 70872 71617
rect 70838 71515 70872 71549
rect 70838 71447 70872 71481
rect 70838 71379 70872 71413
rect 70838 71311 70872 71345
rect 70838 71243 70872 71277
rect 70838 71175 70872 71209
rect 70838 71107 70872 71141
rect 70838 71039 70872 71073
rect 70838 70971 70872 71005
rect 70838 70903 70872 70937
rect 70838 70835 70872 70869
rect 70838 70767 70872 70801
rect 70838 70699 70872 70733
rect 70838 70631 70872 70665
rect 70838 70563 70872 70597
rect 70838 70495 70872 70529
rect 70838 70427 70872 70461
rect 70838 70359 70872 70393
rect 70838 70291 70872 70325
rect 70838 70223 70872 70257
rect 70838 70155 70872 70189
rect 70838 70087 70872 70121
rect 70838 70019 70872 70053
rect 70838 69951 70872 69985
rect 70838 69883 70872 69917
rect 70838 69815 70872 69849
rect 70838 69747 70872 69781
rect 70838 69679 70872 69713
rect 70838 69611 70872 69645
rect 70838 69543 70872 69577
rect 70838 69475 70872 69509
rect 70838 69407 70872 69441
rect 70838 69339 70872 69373
rect 70838 69271 70872 69305
rect 70838 69203 70872 69237
rect 70838 69135 70872 69169
rect 70838 69067 70872 69101
rect 70838 68999 70872 69033
rect 70838 68931 70872 68965
rect 70838 68863 70872 68897
rect 70838 68795 70872 68829
rect 70838 68727 70872 68761
rect 70838 68659 70872 68693
rect 70838 68591 70872 68625
rect 70838 68523 70872 68557
rect 70838 68455 70872 68489
rect 70838 68387 70872 68421
rect 70838 68319 70872 68353
rect 70838 68251 70872 68285
rect 70838 68183 70872 68217
rect 70838 68115 70872 68149
rect 70838 68047 70872 68081
rect 70838 67979 70872 68013
rect 70838 67911 70872 67945
rect 70838 67843 70872 67877
rect 70838 67775 70872 67809
rect 70838 67707 70872 67741
rect 70838 67639 70872 67673
rect 70838 67571 70872 67605
rect 70838 67503 70872 67537
rect 70838 67435 70872 67469
rect 70838 67367 70872 67401
rect 70838 67299 70872 67333
rect 70838 67231 70872 67265
rect 70838 67163 70872 67197
rect 70838 67095 70872 67129
rect 70838 67027 70872 67061
rect 70838 66959 70872 66993
rect 70838 66891 70872 66925
rect 70838 66823 70872 66857
rect 70838 66755 70872 66789
rect 70838 66687 70872 66721
rect 70838 66619 70872 66653
rect 70838 66551 70872 66585
rect 70838 66483 70872 66517
rect 70838 66415 70872 66449
rect 70838 66347 70872 66381
rect 70838 66279 70872 66313
rect 70838 66211 70872 66245
rect 70838 66143 70872 66177
rect 70838 66075 70872 66109
rect 70838 66007 70872 66041
rect 70838 65939 70872 65973
rect 70838 65871 70872 65905
rect 70838 65803 70872 65837
rect 70838 65735 70872 65769
rect 70838 65667 70872 65701
rect 70838 65599 70872 65633
rect 70838 65531 70872 65565
rect 70838 65463 70872 65497
rect 70838 65395 70872 65429
rect 70838 65327 70872 65361
rect 70838 65259 70872 65293
rect 70838 65191 70872 65225
rect 70838 65123 70872 65157
rect 70838 65055 70872 65089
rect 70838 64987 70872 65021
rect 70838 64919 70872 64953
rect 70838 64851 70872 64885
rect 70838 64783 70872 64817
rect 70838 64715 70872 64749
rect 70838 64647 70872 64681
rect 70838 64579 70872 64613
rect 70838 64511 70872 64545
rect 70838 64443 70872 64477
rect 70838 64375 70872 64409
rect 70838 64307 70872 64341
rect 70838 64239 70872 64273
rect 70838 64171 70872 64205
rect 70838 64103 70872 64137
rect 70838 64035 70872 64069
rect 70838 63967 70872 64001
rect 70838 63899 70872 63933
rect 70838 63831 70872 63865
rect 70838 63763 70872 63797
rect 70838 63695 70872 63729
rect 70838 63627 70872 63661
rect 70838 63559 70872 63593
rect 70838 63491 70872 63525
rect 70838 63423 70872 63457
rect 70838 63355 70872 63389
rect 70838 63287 70872 63321
rect 70838 63219 70872 63253
rect 70838 63151 70872 63185
rect 70838 63083 70872 63117
rect 70838 63015 70872 63049
rect 70838 62947 70872 62981
rect 70838 62879 70872 62913
rect 70838 62811 70872 62845
rect 70838 62743 70872 62777
rect 70838 62675 70872 62709
rect 70838 62607 70872 62641
rect 70838 62539 70872 62573
rect 70838 62471 70872 62505
rect 70838 62403 70872 62437
rect 70838 62335 70872 62369
rect 70838 62267 70872 62301
rect 70838 62199 70872 62233
rect 70838 62131 70872 62165
rect 70838 62063 70872 62097
rect 70838 61995 70872 62029
rect 70838 61927 70872 61961
rect 70838 61859 70872 61893
rect 70838 61791 70872 61825
rect 70838 61723 70872 61757
rect 70838 61655 70872 61689
rect 70838 61587 70872 61621
rect 70838 61519 70872 61553
rect 70838 61451 70872 61485
rect 70838 61383 70872 61417
rect 70838 61315 70872 61349
rect 70838 61247 70872 61281
rect 70838 61179 70872 61213
rect 70838 61111 70872 61145
rect 70838 61043 70872 61077
rect 70838 60975 70872 61009
rect 70838 60907 70872 60941
rect 70838 60839 70872 60873
rect 70838 60771 70872 60805
rect 70838 60703 70872 60737
rect 70838 60635 70872 60669
rect 70838 60567 70872 60601
rect 70838 60499 70872 60533
rect 70838 60431 70872 60465
rect 70838 60363 70872 60397
rect 70838 60295 70872 60329
rect 70838 60227 70872 60261
rect 70838 60159 70872 60193
rect 70838 60091 70872 60125
rect 70838 60023 70872 60057
rect 70838 59955 70872 59989
rect 70838 59887 70872 59921
rect 70838 59819 70872 59853
rect 70838 59751 70872 59785
rect 70838 59683 70872 59717
rect 70838 59615 70872 59649
rect 70838 59547 70872 59581
rect 70838 59479 70872 59513
rect 70838 59411 70872 59445
rect 70838 59343 70872 59377
rect 70838 59275 70872 59309
rect 70838 59207 70872 59241
rect 70838 59139 70872 59173
rect 70838 59071 70872 59105
rect 70838 59003 70872 59037
rect 70838 58935 70872 58969
rect 70838 58867 70872 58901
rect 70838 58799 70872 58833
rect 70838 58731 70872 58765
rect 70838 58663 70872 58697
rect 70838 58595 70872 58629
rect 70838 58527 70872 58561
rect 70838 58459 70872 58493
rect 70838 58391 70872 58425
rect 70838 58323 70872 58357
rect 70838 58255 70872 58289
rect 70838 58187 70872 58221
rect 70838 58119 70872 58153
rect 70838 58051 70872 58085
rect 70838 57983 70872 58017
rect 70838 57915 70872 57949
rect 70838 57847 70872 57881
rect 70838 57779 70872 57813
rect 70838 57711 70872 57745
rect 70838 57643 70872 57677
rect 70838 57575 70872 57609
rect 70838 57507 70872 57541
rect 70838 57439 70872 57473
rect 70838 57371 70872 57405
rect 70838 57303 70872 57337
rect 70838 57235 70872 57269
rect 70838 57167 70872 57201
rect 70838 57099 70872 57133
rect 70838 57031 70872 57065
rect 70838 56963 70872 56997
rect 70838 56895 70872 56929
rect 70838 56827 70872 56861
rect 70838 56759 70872 56793
rect 70838 56691 70872 56725
rect 70838 56623 70872 56657
rect 70838 56555 70872 56589
rect 70838 56487 70872 56521
rect 70838 56419 70872 56453
rect 70838 56351 70872 56385
rect 70838 56283 70872 56317
rect 70838 56215 70872 56249
rect 70838 56147 70872 56181
rect 70838 56079 70872 56113
rect 70838 56011 70872 56045
rect 70838 55943 70872 55977
rect 70838 55875 70872 55909
rect 70838 55807 70872 55841
rect 70838 55739 70872 55773
rect 70838 55671 70872 55705
rect 70838 55603 70872 55637
rect 70838 55535 70872 55569
rect 70838 55467 70872 55501
rect 70838 55399 70872 55433
rect 70838 55331 70872 55365
rect 70838 55263 70872 55297
rect 70838 55195 70872 55229
rect 70838 55127 70872 55161
rect 70838 55059 70872 55093
rect 70838 54991 70872 55025
rect 70838 54923 70872 54957
rect 70838 54855 70872 54889
rect 70838 54787 70872 54821
rect 70838 54719 70872 54753
rect 70838 54651 70872 54685
rect 70838 54583 70872 54617
rect 70838 54515 70872 54549
rect 70838 54447 70872 54481
rect 70838 54379 70872 54413
rect 70838 54311 70872 54345
rect 70838 54243 70872 54277
rect 70838 54175 70872 54209
rect 70838 54107 70872 54141
rect 70838 54039 70872 54073
rect 70838 53971 70872 54005
rect 70838 53903 70872 53937
rect 70838 53835 70872 53869
rect 70838 53767 70872 53801
rect 70838 53699 70872 53733
rect 70838 53631 70872 53665
rect 70838 53563 70872 53597
rect 70838 53495 70872 53529
rect 70838 53427 70872 53461
rect 70838 53359 70872 53393
rect 70838 53291 70872 53325
rect 70838 53223 70872 53257
rect 70838 53155 70872 53189
rect 70838 53087 70872 53121
rect 70838 53019 70872 53053
rect 70838 52951 70872 52985
rect 70838 52883 70872 52917
rect 70838 52815 70872 52849
rect 70838 52747 70872 52781
rect 70838 52679 70872 52713
rect 70838 52611 70872 52645
rect 70838 52543 70872 52577
rect 70838 52475 70872 52509
rect 70838 52407 70872 52441
rect 70838 52339 70872 52373
rect 70838 52271 70872 52305
rect 70838 52203 70872 52237
rect 70838 52135 70872 52169
rect 70838 52067 70872 52101
rect 70838 51999 70872 52033
rect 70838 51931 70872 51965
rect 70838 51863 70872 51897
rect 70838 51795 70872 51829
rect 70838 51727 70872 51761
rect 70838 51659 70872 51693
rect 70838 51591 70872 51625
rect 70838 51523 70872 51557
rect 70838 51455 70872 51489
rect 70838 51387 70872 51421
rect 70838 51319 70872 51353
rect 70838 51251 70872 51285
rect 70838 51183 70872 51217
rect 70838 51115 70872 51149
rect 70838 51047 70872 51081
rect 70838 50979 70872 51013
rect 70838 50911 70872 50945
rect 70838 50843 70872 50877
rect 70838 50775 70872 50809
rect 70838 50707 70872 50741
rect 70838 50639 70872 50673
rect 70838 50571 70872 50605
rect 70838 50503 70872 50537
rect 70838 50435 70872 50469
rect 70838 50367 70872 50401
rect 70838 50299 70872 50333
rect 70838 50231 70872 50265
rect 70838 50163 70872 50197
rect 70838 50095 70872 50129
rect 70838 50027 70872 50061
rect 70838 49959 70872 49993
rect 70838 49891 70872 49925
rect 70838 49823 70872 49857
rect 70838 49755 70872 49789
rect 70838 49687 70872 49721
rect 70838 49619 70872 49653
rect 70838 49551 70872 49585
rect 70838 49483 70872 49517
rect 70838 49415 70872 49449
rect 70838 49347 70872 49381
rect 70838 49279 70872 49313
rect 70838 49211 70872 49245
rect 70838 49143 70872 49177
rect 70838 49075 70872 49109
rect 70838 49007 70872 49041
rect 70838 48939 70872 48973
rect 70838 48871 70872 48905
rect 70838 48803 70872 48837
rect 70838 48735 70872 48769
rect 70838 48667 70872 48701
rect 70838 48599 70872 48633
rect 70838 48531 70872 48565
rect 70838 48463 70872 48497
rect 70838 48395 70872 48429
rect 70838 48327 70872 48361
rect 70838 48259 70872 48293
rect 70838 48191 70872 48225
rect 70838 48123 70872 48157
rect 70838 48055 70872 48089
rect 70838 47987 70872 48021
rect 70838 47919 70872 47953
rect 70838 47851 70872 47885
rect 70838 47783 70872 47817
rect 70838 47715 70872 47749
rect 70838 47647 70872 47681
rect 70838 47579 70872 47613
rect 70838 47511 70872 47545
rect 70838 47443 70872 47477
rect 70838 47375 70872 47409
rect 70838 47307 70872 47341
rect 70838 47239 70872 47273
rect 70838 47171 70872 47205
rect 70838 47103 70872 47137
rect 70838 47035 70872 47069
rect 70838 46967 70872 47001
rect 70838 46899 70872 46933
rect 70838 46831 70872 46865
rect 70838 46763 70872 46797
rect 70838 46695 70872 46729
rect 70838 46627 70872 46661
rect 70838 46559 70872 46593
rect 70838 46491 70872 46525
rect 70838 46423 70872 46457
rect 70838 46355 70872 46389
rect 70838 46287 70872 46321
rect 70838 46219 70872 46253
rect 70838 46151 70872 46185
rect 70838 46083 70872 46117
rect 70838 46015 70872 46049
rect 70838 45947 70872 45981
rect 59191 45886 59225 45920
rect 59259 45886 59293 45920
rect 59327 45886 59361 45920
rect 59395 45886 59429 45920
rect 59463 45886 59497 45920
rect 59531 45886 59565 45920
rect 59599 45886 59633 45920
rect 59667 45886 59701 45920
rect 59735 45886 59769 45920
rect 59803 45886 59837 45920
rect 59871 45886 59905 45920
rect 59939 45886 59973 45920
rect 60007 45886 60041 45920
rect 60075 45886 60109 45920
rect 60143 45886 60177 45920
rect 60211 45886 60245 45920
rect 60279 45886 60313 45920
rect 60347 45886 60381 45920
rect 60415 45886 60449 45920
rect 60483 45886 60517 45920
rect 60551 45886 60585 45920
rect 60619 45886 60653 45920
rect 60687 45886 60721 45920
rect 60755 45886 60789 45920
rect 60823 45886 60857 45920
rect 60891 45886 60925 45920
rect 60959 45886 60993 45920
rect 61027 45886 61061 45920
rect 61095 45886 61129 45920
rect 61163 45886 61197 45920
rect 61231 45886 61265 45920
rect 61299 45886 61333 45920
rect 61367 45886 61401 45920
rect 61435 45886 61469 45920
rect 61503 45886 61537 45920
rect 61571 45886 61605 45920
rect 61639 45886 61673 45920
rect 61707 45886 61741 45920
rect 61775 45886 61809 45920
rect 61843 45886 61877 45920
rect 61911 45886 61945 45920
rect 61979 45886 62013 45920
rect 62047 45886 62081 45920
rect 62115 45886 62149 45920
rect 62183 45886 62217 45920
rect 62251 45886 62285 45920
rect 62319 45886 62353 45920
rect 62387 45886 62421 45920
rect 62455 45886 62489 45920
rect 62523 45886 62557 45920
rect 62591 45886 62625 45920
rect 62659 45886 62693 45920
rect 62727 45886 62761 45920
rect 62795 45886 62829 45920
rect 62863 45886 62897 45920
rect 62931 45886 62965 45920
rect 62999 45886 63033 45920
rect 63067 45886 63101 45920
rect 63135 45886 63169 45920
rect 63203 45886 63237 45920
rect 63271 45886 63305 45920
rect 63339 45886 63373 45920
rect 63407 45886 63441 45920
rect 63475 45886 63509 45920
rect 63543 45886 63577 45920
rect 63611 45886 63645 45920
rect 63679 45886 63713 45920
rect 63747 45886 63781 45920
rect 63815 45886 63849 45920
rect 63883 45886 63917 45920
rect 63951 45886 63985 45920
rect 64019 45886 64053 45920
rect 64087 45886 64121 45920
rect 64155 45886 64189 45920
rect 64223 45886 64257 45920
rect 64291 45886 64325 45920
rect 64359 45886 64393 45920
rect 64427 45886 64461 45920
rect 64495 45886 64529 45920
rect 64563 45886 64597 45920
rect 64631 45886 64665 45920
rect 64699 45886 64733 45920
rect 64767 45886 64801 45920
rect 64835 45886 64869 45920
rect 64903 45886 64937 45920
rect 64971 45886 65005 45920
rect 65039 45886 65073 45920
rect 65107 45886 65141 45920
rect 65175 45886 65209 45920
rect 65243 45886 65277 45920
rect 65311 45886 65345 45920
rect 65379 45886 65413 45920
rect 65447 45886 65481 45920
rect 65515 45886 65549 45920
rect 65583 45886 65617 45920
rect 65651 45886 65685 45920
rect 65719 45886 65753 45920
rect 65787 45886 65821 45920
rect 65855 45886 65889 45920
rect 65923 45886 65957 45920
rect 65991 45886 66025 45920
rect 66059 45886 66093 45920
rect 66127 45886 66161 45920
rect 66195 45886 66229 45920
rect 66263 45886 66297 45920
rect 66331 45886 66365 45920
rect 66399 45886 66433 45920
rect 66467 45886 66501 45920
rect 66535 45886 66569 45920
rect 66603 45886 66637 45920
rect 66671 45886 66705 45920
rect 66739 45886 66773 45920
rect 66807 45886 66841 45920
rect 66875 45886 66909 45920
rect 66943 45886 66977 45920
rect 67011 45886 67045 45920
rect 67079 45886 67113 45920
rect 67147 45886 67181 45920
rect 67215 45886 67249 45920
rect 67283 45886 67317 45920
rect 67351 45886 67385 45920
rect 67419 45886 67453 45920
rect 67487 45886 67521 45920
rect 67555 45886 67589 45920
rect 67623 45886 67657 45920
rect 67691 45886 67725 45920
rect 67759 45886 67793 45920
rect 67827 45886 67861 45920
rect 67895 45886 67929 45920
rect 67963 45886 67997 45920
rect 68031 45886 68065 45920
rect 68099 45886 68133 45920
rect 68167 45886 68201 45920
rect 68235 45886 68269 45920
rect 68303 45886 68337 45920
rect 68371 45886 68405 45920
rect 68439 45886 68473 45920
rect 68507 45886 68541 45920
rect 68575 45886 68609 45920
rect 68643 45886 68677 45920
rect 68711 45886 68745 45920
rect 68779 45886 68813 45920
rect 68847 45886 68881 45920
rect 68915 45886 68949 45920
rect 68983 45886 69017 45920
rect 69051 45886 69085 45920
rect 69119 45886 69153 45920
rect 69187 45886 69221 45920
rect 69255 45886 69289 45920
rect 69323 45886 69357 45920
rect 69391 45886 69425 45920
rect 69459 45886 69493 45920
rect 69527 45886 69561 45920
rect 69595 45886 69629 45920
rect 69663 45886 69697 45920
rect 69731 45886 69765 45920
rect 69799 45886 69833 45920
rect 69867 45886 69901 45920
rect 69935 45886 69969 45920
rect 70003 45886 70037 45920
rect 70071 45886 70105 45920
rect 70139 45886 70173 45920
rect 70207 45886 70241 45920
rect 70275 45886 70309 45920
rect 70343 45886 70377 45920
rect 70411 45886 70445 45920
rect 70479 45886 70513 45920
rect 70547 45886 70581 45920
rect 70615 45886 70649 45920
rect 70683 45886 70717 45920
rect 70751 45886 70785 45920
rect -3718 45830 -3684 45864
rect -3718 45762 -3684 45796
rect -3718 45694 -3684 45728
rect -3718 45626 -3684 45660
rect -3718 45558 -3684 45592
rect -3718 45490 -3684 45524
rect -3718 45422 -3684 45456
rect -3718 45354 -3684 45388
rect -3718 45286 -3684 45320
rect -3718 45218 -3684 45252
rect -3718 45150 -3684 45184
rect -3718 45082 -3684 45116
rect -3718 45014 -3684 45048
rect -3718 44946 -3684 44980
rect -3718 44878 -3684 44912
rect -3718 44810 -3684 44844
rect -3718 44742 -3684 44776
rect -3718 44674 -3684 44708
rect -3718 44606 -3684 44640
rect -3718 44538 -3684 44572
rect -3718 44470 -3684 44504
rect -3718 44402 -3684 44436
rect -3718 44334 -3684 44368
rect -10609 44246 -10575 44280
rect -10541 44246 -10507 44280
rect -10473 44246 -10439 44280
rect -10405 44246 -10371 44280
rect -10337 44246 -10303 44280
rect -10269 44246 -10235 44280
rect -10201 44246 -10167 44280
rect -10133 44246 -10099 44280
rect -10065 44246 -10031 44280
rect -9997 44246 -9963 44280
rect -9929 44246 -9895 44280
rect -9861 44246 -9827 44280
rect -9793 44246 -9759 44280
rect -9725 44246 -9691 44280
rect -9657 44246 -9623 44280
rect -9589 44246 -9555 44280
rect -9521 44246 -9487 44280
rect -9453 44246 -9419 44280
rect -9385 44246 -9351 44280
rect -9317 44246 -9283 44280
rect -9249 44246 -9215 44280
rect -9181 44246 -9147 44280
rect -9113 44246 -9079 44280
rect -9045 44246 -9011 44280
rect -8977 44246 -8943 44280
rect -8909 44246 -8875 44280
rect -8841 44246 -8807 44280
rect -8773 44246 -8739 44280
rect -8705 44246 -8671 44280
rect -8637 44246 -8603 44280
rect -8569 44246 -8535 44280
rect -8501 44246 -8467 44280
rect -8433 44246 -8399 44280
rect -8365 44246 -8331 44280
rect -8297 44246 -8263 44280
rect -8229 44246 -8195 44280
rect -8161 44246 -8127 44280
rect -8093 44246 -8059 44280
rect -8025 44246 -7991 44280
rect -7957 44246 -7923 44280
rect -7889 44246 -7855 44280
rect -7821 44246 -7787 44280
rect -7753 44246 -7719 44280
rect -7685 44246 -7651 44280
rect -7617 44246 -7583 44280
rect -7549 44246 -7515 44280
rect -7481 44246 -7447 44280
rect -7413 44246 -7379 44280
rect -7345 44246 -7311 44280
rect -7277 44246 -7243 44280
rect -7209 44246 -7175 44280
rect -7141 44246 -7107 44280
rect -7073 44246 -7039 44280
rect -7005 44246 -6971 44280
rect -6937 44246 -6903 44280
rect -6869 44246 -6835 44280
rect -6801 44246 -6767 44280
rect -6733 44246 -6699 44280
rect -6665 44246 -6631 44280
rect -6597 44246 -6563 44280
rect -6529 44246 -6495 44280
rect -6461 44246 -6427 44280
rect -6393 44246 -6359 44280
rect -6325 44246 -6291 44280
rect -6257 44246 -6223 44280
rect -6189 44246 -6155 44280
rect -6121 44246 -6087 44280
rect -6053 44246 -6019 44280
rect -5985 44246 -5951 44280
rect -5917 44246 -5883 44280
rect -5849 44246 -5815 44280
rect -5781 44246 -5747 44280
rect -5713 44246 -5679 44280
rect -5645 44246 -5611 44280
rect -5577 44246 -5543 44280
rect -5509 44246 -5475 44280
rect -5441 44246 -5407 44280
rect -5373 44246 -5339 44280
rect -5305 44246 -5271 44280
rect -5237 44246 -5203 44280
rect -5169 44246 -5135 44280
rect -5101 44246 -5067 44280
rect -5033 44246 -4999 44280
rect -4965 44246 -4931 44280
rect -4897 44246 -4863 44280
rect -4829 44246 -4795 44280
rect -4761 44246 -4727 44280
rect -4693 44246 -4659 44280
rect -4625 44246 -4591 44280
rect -4557 44246 -4523 44280
rect -4489 44246 -4455 44280
rect -4421 44246 -4387 44280
rect -4353 44246 -4319 44280
rect -4285 44246 -4251 44280
rect -4217 44246 -4183 44280
rect -4149 44246 -4115 44280
rect -4081 44246 -4047 44280
rect -4013 44246 -3979 44280
rect -3945 44246 -3911 44280
rect -3877 44246 -3843 44280
rect -3809 44246 -3775 44280
rect -2318 19487 -2284 19521
rect -2250 19487 -2216 19521
rect -2182 19487 -2148 19521
rect -2114 19487 -2080 19521
rect -2046 19487 -2012 19521
rect -1978 19487 -1944 19521
rect -1910 19487 -1876 19521
rect -1842 19487 -1808 19521
rect -1774 19487 -1740 19521
rect -1706 19487 -1672 19521
rect -1638 19487 -1604 19521
rect -1570 19487 -1536 19521
rect -1502 19487 -1468 19521
rect -1434 19487 -1400 19521
rect -1366 19487 -1332 19521
rect -1298 19487 -1264 19521
rect -1230 19487 -1196 19521
rect -1162 19487 -1128 19521
rect -1094 19487 -1060 19521
rect -1026 19487 -992 19521
rect -958 19487 -924 19521
rect -890 19487 -856 19521
rect -822 19487 -788 19521
rect -754 19487 -720 19521
rect -686 19487 -652 19521
rect -618 19487 -584 19521
rect -550 19487 -516 19521
rect -482 19487 -448 19521
rect -414 19487 -380 19521
rect -346 19487 -312 19521
rect -278 19487 -244 19521
rect -210 19487 -176 19521
rect -142 19487 -108 19521
rect -74 19487 -40 19521
rect -6 19487 28 19521
rect 62 19487 96 19521
rect 130 19487 164 19521
rect 198 19487 232 19521
rect 266 19487 300 19521
rect 334 19487 368 19521
rect 402 19487 436 19521
rect 470 19487 504 19521
rect 538 19487 572 19521
rect 606 19487 640 19521
rect 674 19487 708 19521
rect 742 19487 776 19521
rect 810 19487 844 19521
rect 878 19487 912 19521
rect 946 19487 980 19521
rect 1014 19487 1048 19521
rect 1082 19487 1116 19521
rect 1150 19487 1184 19521
rect 1218 19487 1252 19521
rect 1286 19487 1320 19521
rect 1354 19487 1388 19521
rect 1422 19487 1456 19521
rect 1490 19487 1524 19521
rect 1558 19487 1592 19521
rect 1626 19487 1660 19521
rect 1694 19487 1728 19521
rect 1762 19487 1796 19521
rect 1830 19487 1864 19521
rect 1898 19487 1932 19521
rect 1966 19487 2000 19521
rect 2034 19487 2068 19521
rect 2102 19487 2136 19521
rect 2170 19487 2204 19521
rect 2238 19487 2272 19521
rect 2306 19487 2340 19521
rect 2374 19487 2408 19521
rect 2442 19487 2476 19521
rect 2510 19487 2544 19521
rect 2578 19487 2612 19521
rect 2646 19487 2680 19521
rect 2714 19487 2748 19521
rect 2782 19487 2816 19521
rect 2850 19487 2884 19521
rect 2918 19487 2952 19521
rect 2986 19487 3020 19521
rect 3054 19487 3088 19521
rect 3122 19487 3156 19521
rect 3190 19487 3224 19521
rect 3258 19487 3292 19521
rect 3326 19487 3360 19521
rect 3394 19487 3428 19521
rect 3462 19487 3496 19521
rect 3530 19487 3564 19521
rect 3598 19487 3632 19521
rect 3666 19487 3700 19521
rect 3734 19487 3768 19521
rect 3802 19487 3836 19521
rect 3870 19487 3904 19521
rect 3938 19487 3972 19521
rect 4006 19487 4040 19521
rect 4074 19487 4108 19521
rect 4142 19487 4176 19521
rect 4210 19487 4244 19521
rect 4278 19487 4312 19521
rect 4346 19487 4380 19521
rect 4414 19487 4448 19521
rect 4482 19487 4516 19521
rect 4550 19487 4584 19521
rect 4618 19487 4652 19521
rect 4686 19487 4720 19521
rect 4754 19487 4788 19521
rect 4822 19487 4856 19521
rect 4890 19487 4924 19521
rect 4958 19487 4992 19521
rect 5026 19487 5060 19521
rect 5094 19487 5128 19521
rect 5162 19487 5196 19521
rect 5230 19487 5264 19521
rect 5298 19487 5332 19521
rect 5366 19487 5400 19521
rect 5434 19487 5468 19521
rect 5502 19487 5536 19521
rect 5570 19487 5604 19521
rect 5638 19487 5672 19521
rect 5706 19487 5740 19521
rect 5774 19487 5808 19521
rect 5842 19487 5876 19521
rect 5910 19487 5944 19521
rect 5978 19487 6012 19521
rect 6046 19487 6080 19521
rect 6114 19487 6148 19521
rect 6182 19487 6216 19521
rect 6250 19487 6284 19521
rect 6318 19487 6352 19521
rect 6386 19487 6420 19521
rect 6454 19487 6488 19521
rect 6522 19487 6556 19521
rect 6590 19487 6624 19521
rect 6658 19487 6692 19521
rect 6726 19487 6760 19521
rect 6794 19487 6828 19521
rect 6862 19487 6896 19521
rect 6930 19487 6964 19521
rect 6998 19487 7032 19521
rect 7066 19487 7100 19521
rect 7134 19487 7168 19521
rect 7202 19487 7236 19521
rect 7270 19487 7304 19521
rect 7338 19487 7372 19521
rect 7406 19487 7440 19521
rect 7474 19487 7508 19521
rect 7542 19487 7576 19521
rect 7610 19487 7644 19521
rect 7678 19487 7712 19521
rect 7746 19487 7780 19521
rect 7814 19487 7848 19521
rect 7882 19487 7916 19521
rect 7950 19487 7984 19521
rect 8018 19487 8052 19521
rect 8086 19487 8120 19521
rect 8154 19487 8188 19521
rect 8222 19487 8256 19521
rect 8290 19487 8324 19521
rect 8358 19487 8392 19521
rect 8426 19487 8460 19521
rect 8494 19487 8528 19521
rect 8562 19487 8596 19521
rect 8630 19487 8664 19521
rect 8698 19487 8732 19521
rect 8766 19487 8800 19521
rect 8834 19487 8868 19521
rect 8902 19487 8936 19521
rect 8970 19487 9004 19521
rect 9038 19487 9072 19521
rect 9106 19487 9140 19521
rect 9174 19487 9208 19521
rect 9242 19487 9276 19521
rect 9310 19487 9344 19521
rect 9378 19487 9412 19521
rect 9446 19487 9480 19521
rect 9514 19487 9548 19521
rect 9582 19487 9616 19521
rect 9650 19487 9684 19521
rect 9718 19487 9752 19521
rect 9786 19487 9820 19521
rect 9854 19487 9888 19521
rect 9922 19487 9956 19521
rect 9990 19487 10024 19521
rect 10058 19487 10092 19521
rect 10126 19487 10160 19521
rect 10194 19487 10228 19521
rect 10262 19487 10296 19521
rect 10330 19487 10364 19521
rect 10398 19487 10432 19521
rect 10466 19487 10500 19521
rect 10534 19487 10568 19521
rect 10602 19487 10636 19521
rect 10670 19487 10704 19521
rect 10738 19487 10772 19521
rect 10806 19487 10840 19521
rect 10874 19487 10908 19521
rect 10942 19487 10976 19521
rect 11010 19487 11044 19521
rect 11078 19487 11112 19521
rect 11146 19487 11180 19521
rect 11214 19487 11248 19521
rect 11282 19487 11316 19521
rect 11350 19487 11384 19521
rect 11418 19487 11452 19521
rect 11486 19487 11520 19521
rect 11554 19487 11588 19521
rect 11622 19487 11656 19521
rect 11690 19487 11724 19521
rect 11758 19487 11792 19521
rect 11826 19487 11860 19521
rect 11894 19487 11928 19521
rect 11962 19487 11996 19521
rect 12030 19487 12064 19521
rect 12098 19487 12132 19521
rect 12166 19487 12200 19521
rect 12234 19487 12268 19521
rect 12302 19487 12336 19521
rect 12370 19487 12404 19521
rect 12438 19487 12472 19521
rect 12506 19487 12540 19521
rect 12574 19487 12608 19521
rect 12642 19487 12676 19521
rect 12710 19487 12744 19521
rect 12778 19487 12812 19521
rect 12846 19487 12880 19521
rect 12914 19487 12948 19521
rect 12982 19487 13016 19521
rect 13050 19487 13084 19521
rect 13118 19487 13152 19521
rect 13186 19487 13220 19521
rect 13254 19487 13288 19521
rect 13322 19487 13356 19521
rect 13390 19487 13424 19521
rect 13458 19487 13492 19521
rect 13526 19487 13560 19521
rect 13594 19487 13628 19521
rect 13662 19487 13696 19521
rect 13730 19487 13764 19521
rect 13798 19487 13832 19521
rect 13866 19487 13900 19521
rect 13934 19487 13968 19521
rect 14002 19487 14036 19521
rect 14070 19487 14104 19521
rect 14138 19487 14172 19521
rect 14206 19487 14240 19521
rect 14274 19487 14308 19521
rect 14342 19487 14376 19521
rect 14410 19487 14444 19521
rect 14478 19487 14512 19521
rect 14546 19487 14580 19521
rect 14614 19487 14648 19521
rect 14682 19487 14716 19521
rect 14750 19487 14784 19521
rect 14818 19487 14852 19521
rect 14886 19487 14920 19521
rect 14954 19487 14988 19521
rect 15022 19487 15056 19521
rect 15090 19487 15124 19521
rect 15158 19487 15192 19521
rect 15226 19487 15260 19521
rect 15294 19487 15328 19521
rect 15362 19487 15396 19521
rect 15430 19487 15464 19521
rect 15498 19487 15532 19521
rect 15566 19487 15600 19521
rect 15634 19487 15668 19521
rect 15702 19487 15736 19521
rect 15770 19487 15804 19521
rect 15838 19487 15872 19521
rect 15906 19487 15940 19521
rect 15974 19487 16008 19521
rect 16042 19487 16076 19521
rect 16110 19487 16144 19521
rect 16178 19487 16212 19521
rect 16246 19487 16280 19521
rect 16314 19487 16348 19521
rect 16382 19487 16416 19521
rect 16450 19487 16484 19521
rect 16518 19487 16552 19521
rect 16586 19487 16620 19521
rect 16654 19487 16688 19521
rect 16722 19487 16756 19521
rect 16790 19487 16824 19521
rect 16858 19487 16892 19521
rect 16926 19487 16960 19521
rect 16994 19487 17028 19521
rect 17062 19487 17096 19521
rect 17130 19487 17164 19521
rect 17198 19487 17232 19521
rect 17266 19487 17300 19521
rect 17334 19487 17368 19521
rect 17402 19487 17436 19521
rect 17470 19487 17504 19521
rect 17538 19487 17572 19521
rect 17606 19487 17640 19521
rect 17674 19487 17708 19521
rect 17742 19487 17776 19521
rect 17810 19487 17844 19521
rect 17878 19487 17912 19521
rect 17946 19487 17980 19521
rect 18014 19487 18048 19521
rect 18082 19487 18116 19521
rect 18150 19487 18184 19521
rect 18218 19487 18252 19521
rect 18286 19487 18320 19521
rect 18354 19487 18388 19521
rect 18422 19487 18456 19521
rect 18490 19487 18524 19521
rect 18558 19487 18592 19521
rect 18626 19487 18660 19521
rect 18694 19487 18728 19521
rect 18762 19487 18796 19521
rect 18830 19487 18864 19521
rect 18898 19487 18932 19521
rect 18966 19487 19000 19521
rect 19034 19487 19068 19521
rect 19102 19487 19136 19521
rect 19170 19487 19204 19521
rect 19238 19487 19272 19521
rect 19306 19487 19340 19521
rect 19374 19487 19408 19521
rect 19442 19487 19476 19521
rect 19510 19487 19544 19521
rect 19578 19487 19612 19521
rect 19646 19487 19680 19521
rect 19714 19487 19748 19521
rect 19782 19487 19816 19521
rect 19850 19487 19884 19521
rect 19918 19487 19952 19521
rect 19986 19487 20020 19521
rect 20054 19487 20088 19521
rect 20122 19487 20156 19521
rect 20190 19487 20224 19521
rect 20258 19487 20292 19521
rect 20326 19487 20360 19521
rect 20394 19487 20428 19521
rect 20462 19487 20496 19521
rect 20530 19487 20564 19521
rect 20598 19487 20632 19521
rect 20666 19487 20700 19521
rect 20734 19487 20768 19521
rect 20802 19487 20836 19521
rect 20870 19487 20904 19521
rect 20938 19487 20972 19521
rect 21006 19487 21040 19521
rect 21074 19487 21108 19521
rect 21142 19487 21176 19521
rect 21210 19487 21244 19521
rect 21278 19487 21312 19521
rect 21346 19487 21380 19521
rect 21414 19487 21448 19521
rect 21482 19487 21516 19521
rect 21550 19487 21584 19521
rect 21618 19487 21652 19521
rect 21686 19487 21720 19521
rect 21754 19487 21788 19521
rect 21822 19487 21856 19521
rect 21890 19487 21924 19521
rect 21958 19487 21992 19521
rect 22026 19487 22060 19521
rect 22094 19487 22128 19521
rect 22162 19487 22196 19521
rect 22230 19487 22264 19521
rect 22298 19487 22332 19521
rect 22366 19487 22400 19521
rect 22434 19487 22468 19521
rect 22502 19487 22536 19521
rect 22570 19487 22604 19521
rect 22638 19487 22672 19521
rect 22706 19487 22740 19521
rect 22774 19487 22808 19521
rect 22842 19487 22876 19521
rect 22910 19487 22944 19521
rect 22978 19487 23012 19521
rect 23046 19487 23080 19521
rect 23114 19487 23148 19521
rect 23182 19487 23216 19521
rect 23250 19487 23284 19521
rect 23318 19487 23352 19521
rect 23386 19487 23420 19521
rect 23454 19487 23488 19521
rect 23522 19487 23556 19521
rect 23590 19487 23624 19521
rect 23658 19487 23692 19521
rect 23726 19487 23760 19521
rect 23794 19487 23828 19521
rect 23862 19487 23896 19521
rect 23930 19487 23964 19521
rect 23998 19487 24032 19521
rect 24066 19487 24100 19521
rect 24134 19487 24168 19521
rect 24202 19487 24236 19521
rect 24270 19487 24304 19521
rect 24338 19487 24372 19521
rect 24406 19487 24440 19521
rect 24474 19487 24508 19521
rect 24542 19487 24576 19521
rect 24610 19487 24644 19521
rect 24678 19487 24712 19521
rect 24746 19487 24780 19521
rect 24814 19487 24848 19521
rect 24882 19487 24916 19521
rect 24950 19487 24984 19521
rect 25018 19487 25052 19521
rect 25086 19487 25120 19521
rect 25154 19487 25188 19521
rect 25222 19487 25256 19521
rect 25290 19487 25324 19521
rect 25358 19487 25392 19521
rect 25426 19487 25460 19521
rect 25494 19487 25528 19521
rect 25562 19487 25596 19521
rect 25630 19487 25664 19521
rect 25698 19487 25732 19521
rect 25766 19487 25800 19521
rect 25834 19487 25868 19521
rect 25902 19487 25936 19521
rect 25970 19487 26004 19521
rect 26038 19487 26072 19521
rect 26106 19487 26140 19521
rect 26174 19487 26208 19521
rect 26242 19487 26276 19521
rect 26310 19487 26344 19521
rect 26378 19487 26412 19521
rect 26446 19487 26480 19521
rect 26514 19487 26548 19521
rect 26582 19487 26616 19521
rect 26650 19487 26684 19521
rect 26718 19487 26752 19521
rect 26786 19487 26820 19521
rect 26854 19487 26888 19521
rect 26922 19487 26956 19521
rect 26990 19487 27024 19521
rect 27058 19487 27092 19521
rect 27126 19487 27160 19521
rect 27194 19487 27228 19521
rect 27262 19487 27296 19521
rect 27330 19487 27364 19521
rect 27398 19487 27432 19521
rect 27466 19487 27500 19521
rect 27534 19487 27568 19521
rect 27602 19487 27636 19521
rect 27670 19487 27704 19521
rect 27738 19487 27772 19521
rect 27806 19487 27840 19521
rect 27874 19487 27908 19521
rect 27942 19487 27976 19521
rect 28010 19487 28044 19521
rect 28078 19487 28112 19521
rect 28146 19487 28180 19521
rect 28214 19487 28248 19521
rect 28282 19487 28316 19521
rect 28350 19487 28384 19521
rect 28418 19487 28452 19521
rect 28486 19487 28520 19521
rect 28554 19487 28588 19521
rect 28622 19487 28656 19521
rect 28690 19487 28724 19521
rect 28758 19487 28792 19521
rect 28826 19487 28860 19521
rect 28894 19487 28928 19521
rect 28962 19487 28996 19521
rect 29030 19487 29064 19521
rect 29098 19487 29132 19521
rect 29166 19487 29200 19521
rect 29234 19487 29268 19521
rect 29302 19487 29336 19521
rect 29370 19487 29404 19521
rect 29438 19487 29472 19521
rect 29506 19487 29540 19521
rect 29574 19487 29608 19521
rect 29642 19487 29676 19521
rect 29710 19487 29744 19521
rect 29778 19487 29812 19521
rect 29846 19487 29880 19521
rect 29914 19487 29948 19521
rect 29982 19487 30016 19521
rect 30050 19487 30084 19521
rect 30118 19487 30152 19521
rect 30186 19487 30220 19521
rect 30254 19487 30288 19521
rect 30322 19487 30356 19521
rect 30390 19487 30424 19521
rect 30458 19487 30492 19521
rect 30526 19487 30560 19521
rect 30594 19487 30628 19521
rect 30662 19487 30696 19521
rect 30730 19487 30764 19521
rect 30798 19487 30832 19521
rect 30866 19487 30900 19521
rect 30934 19487 30968 19521
rect 31002 19487 31036 19521
rect 31070 19487 31104 19521
rect 31138 19487 31172 19521
rect 31206 19487 31240 19521
rect 31274 19487 31308 19521
rect 31342 19487 31376 19521
rect 31410 19487 31444 19521
rect 31478 19487 31512 19521
rect 31546 19487 31580 19521
rect 31614 19487 31648 19521
rect 31682 19487 31716 19521
rect 31750 19487 31784 19521
rect 31818 19487 31852 19521
rect 31886 19487 31920 19521
rect 31954 19487 31988 19521
rect 32022 19487 32056 19521
rect 32090 19487 32124 19521
rect 32158 19487 32192 19521
rect 32226 19487 32260 19521
rect 32294 19487 32328 19521
rect 32362 19487 32396 19521
rect 32430 19487 32464 19521
rect 32498 19487 32532 19521
rect 32566 19487 32600 19521
rect 32634 19487 32668 19521
rect 32702 19487 32736 19521
rect 32770 19487 32804 19521
rect 32838 19487 32872 19521
rect 32906 19487 32940 19521
rect 32974 19487 33008 19521
rect 33042 19487 33076 19521
rect 33110 19487 33144 19521
rect 33178 19487 33212 19521
rect 33246 19487 33280 19521
rect 33314 19487 33348 19521
rect 33382 19487 33416 19521
rect 33450 19487 33484 19521
rect 33518 19487 33552 19521
rect 33586 19487 33620 19521
rect 33654 19487 33688 19521
rect 33722 19487 33756 19521
rect 33790 19487 33824 19521
rect 33858 19487 33892 19521
rect 33926 19487 33960 19521
rect 33994 19487 34028 19521
rect 34062 19487 34096 19521
rect 34130 19487 34164 19521
rect 34198 19487 34232 19521
rect 34266 19487 34300 19521
rect 34334 19487 34368 19521
rect 34402 19487 34436 19521
rect 34470 19487 34504 19521
rect 34538 19487 34572 19521
rect 34606 19487 34640 19521
rect 34674 19487 34708 19521
rect 34742 19487 34776 19521
rect 34810 19487 34844 19521
rect 34878 19487 34912 19521
rect 34946 19487 34980 19521
rect 35014 19487 35048 19521
rect 35082 19487 35116 19521
rect 35150 19487 35184 19521
rect 35218 19487 35252 19521
rect 35286 19487 35320 19521
rect 35354 19487 35388 19521
rect 35422 19487 35456 19521
rect 35490 19487 35524 19521
rect 35558 19487 35592 19521
rect 35626 19487 35660 19521
rect 35694 19487 35728 19521
rect 35762 19487 35796 19521
rect 35830 19487 35864 19521
rect 35898 19487 35932 19521
rect 35966 19487 36000 19521
rect 36034 19487 36068 19521
rect 36102 19487 36136 19521
rect 36170 19487 36204 19521
rect 36238 19487 36272 19521
rect 36306 19487 36340 19521
rect 36374 19487 36408 19521
rect 36442 19487 36476 19521
rect 36510 19487 36544 19521
rect 36578 19487 36612 19521
rect 36646 19487 36680 19521
rect 36714 19487 36748 19521
rect 36782 19487 36816 19521
rect 36850 19487 36884 19521
rect 36918 19487 36952 19521
rect 36986 19487 37020 19521
rect 37054 19487 37088 19521
rect 37122 19487 37156 19521
rect 37190 19487 37224 19521
rect 37258 19487 37292 19521
rect 37326 19487 37360 19521
rect 37394 19487 37428 19521
rect 37462 19487 37496 19521
rect 37530 19487 37564 19521
rect 37598 19487 37632 19521
rect 37666 19487 37700 19521
rect 37734 19487 37768 19521
rect 37802 19487 37836 19521
rect 37870 19487 37904 19521
rect 37938 19487 37972 19521
rect 38006 19487 38040 19521
rect 38074 19487 38108 19521
rect 38142 19487 38176 19521
rect 38210 19487 38244 19521
rect 38278 19487 38312 19521
rect 38346 19487 38380 19521
rect 38414 19487 38448 19521
rect 38482 19487 38516 19521
rect 38550 19487 38584 19521
rect 38618 19487 38652 19521
rect 38686 19487 38720 19521
rect 38754 19487 38788 19521
rect 38822 19487 38856 19521
rect 38890 19487 38924 19521
rect 38958 19487 38992 19521
rect 39026 19487 39060 19521
rect 39094 19487 39128 19521
rect 39162 19487 39196 19521
rect 39230 19487 39264 19521
rect 39298 19487 39332 19521
rect 39366 19487 39400 19521
rect 39434 19487 39468 19521
rect 39502 19487 39536 19521
rect 39570 19487 39604 19521
rect 39638 19487 39672 19521
rect 39706 19487 39740 19521
rect 39774 19487 39808 19521
rect 39842 19487 39876 19521
rect 39910 19487 39944 19521
rect 39978 19487 40012 19521
rect 40046 19487 40080 19521
rect 40114 19487 40148 19521
rect 40182 19487 40216 19521
rect 40250 19487 40284 19521
rect 40318 19487 40352 19521
rect 40386 19487 40420 19521
rect 40454 19487 40488 19521
rect 40522 19487 40556 19521
rect 40590 19487 40624 19521
rect 40658 19487 40692 19521
rect 40726 19487 40760 19521
rect 40794 19487 40828 19521
rect 40862 19487 40896 19521
rect 40930 19487 40964 19521
rect 40998 19487 41032 19521
rect 41066 19487 41100 19521
rect 41134 19487 41168 19521
rect 41202 19487 41236 19521
rect 41270 19487 41304 19521
rect 41338 19487 41372 19521
rect 41406 19487 41440 19521
rect 41474 19487 41508 19521
rect 41542 19487 41576 19521
rect 41610 19487 41644 19521
rect 41678 19487 41712 19521
rect 41746 19487 41780 19521
rect 41814 19487 41848 19521
rect 41882 19487 41916 19521
rect 41950 19487 41984 19521
rect 42018 19487 42052 19521
rect 42086 19487 42120 19521
rect 42154 19487 42188 19521
rect 42222 19487 42256 19521
rect 42290 19487 42324 19521
rect 42358 19487 42392 19521
rect 42426 19487 42460 19521
rect 42494 19487 42528 19521
rect 42562 19487 42596 19521
rect 42630 19487 42664 19521
rect 42698 19487 42732 19521
rect 42766 19487 42800 19521
rect 42834 19487 42868 19521
rect 42902 19487 42936 19521
rect 42970 19487 43004 19521
rect 43038 19487 43072 19521
rect 43106 19487 43140 19521
rect 43174 19487 43208 19521
rect 43242 19487 43276 19521
rect 43310 19487 43344 19521
rect 43378 19487 43412 19521
rect 43446 19487 43480 19521
rect 43514 19487 43548 19521
rect 43582 19487 43616 19521
rect 43650 19487 43684 19521
rect 43718 19487 43752 19521
rect 43786 19487 43820 19521
rect 43854 19487 43888 19521
rect 43922 19487 43956 19521
rect 43990 19487 44024 19521
rect 44058 19487 44092 19521
rect 44126 19487 44160 19521
rect 44194 19487 44228 19521
rect 44262 19487 44296 19521
rect 44330 19487 44364 19521
rect 44398 19487 44432 19521
rect 44466 19487 44500 19521
rect 44534 19487 44568 19521
rect 44602 19487 44636 19521
rect 44670 19487 44704 19521
rect 44738 19487 44772 19521
rect 44806 19487 44840 19521
rect 44874 19487 44908 19521
rect 44942 19487 44976 19521
rect 45010 19487 45044 19521
rect 45078 19487 45112 19521
rect 45146 19487 45180 19521
rect 45214 19487 45248 19521
rect 45282 19487 45316 19521
rect 45350 19487 45384 19521
rect 45418 19487 45452 19521
rect 45486 19487 45520 19521
rect 45554 19487 45588 19521
rect 45622 19487 45656 19521
rect 45690 19487 45724 19521
rect 45758 19487 45792 19521
rect 45826 19487 45860 19521
rect 45894 19487 45928 19521
rect 45962 19487 45996 19521
rect 46030 19487 46064 19521
rect 46098 19487 46132 19521
rect 46166 19487 46200 19521
rect 46234 19487 46268 19521
rect 46302 19487 46336 19521
rect 46370 19487 46404 19521
rect 46438 19487 46472 19521
rect 46506 19487 46540 19521
rect 46574 19487 46608 19521
rect 46642 19487 46676 19521
rect 46710 19487 46744 19521
rect 46778 19487 46812 19521
rect 46846 19487 46880 19521
rect 46914 19487 46948 19521
rect 46982 19487 47016 19521
rect 47050 19487 47084 19521
rect 47118 19487 47152 19521
rect -2396 19400 -2362 19434
rect -2396 19332 -2362 19366
rect -2396 19264 -2362 19298
rect -2396 19196 -2362 19230
rect -2396 19128 -2362 19162
rect -2396 19060 -2362 19094
rect -2396 18992 -2362 19026
rect -2396 18924 -2362 18958
rect -2396 18856 -2362 18890
rect -2396 18788 -2362 18822
rect -2396 18720 -2362 18754
rect -2396 18652 -2362 18686
rect -2396 18584 -2362 18618
rect -2396 18516 -2362 18550
rect -2396 18448 -2362 18482
rect -2396 18380 -2362 18414
rect -2396 18312 -2362 18346
rect -2396 18244 -2362 18278
rect -2396 18176 -2362 18210
rect -2396 18108 -2362 18142
rect -2396 18040 -2362 18074
rect -2396 17972 -2362 18006
rect -2396 17904 -2362 17938
rect -2396 17836 -2362 17870
rect -2396 17768 -2362 17802
rect -2396 17700 -2362 17734
rect -2396 17632 -2362 17666
rect -2396 17564 -2362 17598
rect -2396 17496 -2362 17530
rect -2396 17428 -2362 17462
rect -2396 17360 -2362 17394
rect -2396 17292 -2362 17326
rect -2396 17224 -2362 17258
rect -2396 17156 -2362 17190
rect -2396 17088 -2362 17122
rect -2396 17020 -2362 17054
rect -2396 16952 -2362 16986
rect -2396 16884 -2362 16918
rect -2396 16816 -2362 16850
rect -2396 16748 -2362 16782
rect -2396 16680 -2362 16714
rect -2396 16612 -2362 16646
rect -2396 16544 -2362 16578
rect -2396 16476 -2362 16510
rect -2396 16408 -2362 16442
rect -2396 16340 -2362 16374
rect -2396 16272 -2362 16306
rect -2396 16204 -2362 16238
rect -2396 16136 -2362 16170
rect -2396 16068 -2362 16102
rect -2396 16000 -2362 16034
rect -2396 15932 -2362 15966
rect -2396 15864 -2362 15898
rect -2396 15796 -2362 15830
rect -2396 15728 -2362 15762
rect -2396 15660 -2362 15694
rect -2396 15592 -2362 15626
rect -2396 15524 -2362 15558
rect -2396 15456 -2362 15490
rect -2396 15388 -2362 15422
rect -2396 15320 -2362 15354
rect -2396 15252 -2362 15286
rect -2396 15184 -2362 15218
rect -2396 15116 -2362 15150
rect -2396 15048 -2362 15082
rect -2396 14980 -2362 15014
rect -2396 14912 -2362 14946
rect -2396 14844 -2362 14878
rect -2396 14776 -2362 14810
rect -2396 14708 -2362 14742
rect -2396 14640 -2362 14674
rect -2396 14572 -2362 14606
rect -2396 14504 -2362 14538
rect -2396 14436 -2362 14470
rect -2396 14368 -2362 14402
rect -2396 14300 -2362 14334
rect -2396 14232 -2362 14266
rect -2396 14164 -2362 14198
rect -2396 14096 -2362 14130
rect -2396 14028 -2362 14062
rect -2396 13960 -2362 13994
rect -2396 13892 -2362 13926
rect -2396 13824 -2362 13858
rect -2396 13756 -2362 13790
rect -2396 13688 -2362 13722
rect -2396 13620 -2362 13654
rect -2396 13552 -2362 13586
rect -2396 13484 -2362 13518
rect -2396 13416 -2362 13450
rect -2396 13348 -2362 13382
rect -2396 13280 -2362 13314
rect -2396 13212 -2362 13246
rect -2396 13144 -2362 13178
rect -2396 13076 -2362 13110
rect -2396 13008 -2362 13042
rect -2396 12940 -2362 12974
rect -2396 12872 -2362 12906
rect -2396 12804 -2362 12838
rect -2396 12736 -2362 12770
rect -2396 12668 -2362 12702
rect -2396 12600 -2362 12634
rect -2396 12532 -2362 12566
rect -2396 12464 -2362 12498
rect -2396 12396 -2362 12430
rect -2396 12328 -2362 12362
rect -2396 12260 -2362 12294
rect -2396 12192 -2362 12226
rect -2396 12124 -2362 12158
rect -2396 12056 -2362 12090
rect -2396 11988 -2362 12022
rect -2396 11920 -2362 11954
rect -2396 11852 -2362 11886
rect -2396 11784 -2362 11818
rect -2396 11716 -2362 11750
rect -2396 11648 -2362 11682
rect -2396 11580 -2362 11614
rect -2396 11512 -2362 11546
rect -2396 11444 -2362 11478
rect -2396 11376 -2362 11410
rect -2396 11308 -2362 11342
rect -2396 11240 -2362 11274
rect -2396 11172 -2362 11206
rect -2396 11104 -2362 11138
rect -2396 11036 -2362 11070
rect -2396 10968 -2362 11002
rect -2396 10900 -2362 10934
rect -2396 10832 -2362 10866
rect -2396 10764 -2362 10798
rect -2396 10696 -2362 10730
rect -2396 10628 -2362 10662
rect -2396 10560 -2362 10594
rect -2396 10492 -2362 10526
rect -2396 10424 -2362 10458
rect -2396 10356 -2362 10390
rect -2396 10288 -2362 10322
rect -2396 10220 -2362 10254
rect -2396 10152 -2362 10186
rect -2396 10084 -2362 10118
rect -2396 10016 -2362 10050
rect -2396 9948 -2362 9982
rect -2396 9880 -2362 9914
rect -2396 9812 -2362 9846
rect -2396 9744 -2362 9778
rect -2396 9676 -2362 9710
rect -2396 9608 -2362 9642
rect -2396 9540 -2362 9574
rect -2396 9472 -2362 9506
rect -2396 9404 -2362 9438
rect -2396 9336 -2362 9370
rect -2396 9268 -2362 9302
rect -2396 9200 -2362 9234
rect -2396 9132 -2362 9166
rect -2396 9064 -2362 9098
rect -2396 8996 -2362 9030
rect -2396 8928 -2362 8962
rect -2396 8860 -2362 8894
rect -2396 8792 -2362 8826
rect -2396 8724 -2362 8758
rect -2396 8656 -2362 8690
rect -2396 8588 -2362 8622
rect -2396 8520 -2362 8554
rect -2396 8452 -2362 8486
rect -2396 8384 -2362 8418
rect -2396 8316 -2362 8350
rect -2396 8248 -2362 8282
rect -2396 8180 -2362 8214
rect -2396 8112 -2362 8146
rect -2396 8044 -2362 8078
rect -2396 7976 -2362 8010
rect -2396 7908 -2362 7942
rect -2396 7840 -2362 7874
rect -2396 7772 -2362 7806
rect -2396 7704 -2362 7738
rect -2396 7636 -2362 7670
rect -2396 7568 -2362 7602
rect -2396 7500 -2362 7534
rect -2396 7432 -2362 7466
rect -2396 7364 -2362 7398
rect -2396 7296 -2362 7330
rect -2396 7228 -2362 7262
rect -2396 7160 -2362 7194
rect -2396 7092 -2362 7126
rect -2396 7024 -2362 7058
rect -2396 6956 -2362 6990
rect -2396 6888 -2362 6922
rect -2396 6820 -2362 6854
rect -2396 6752 -2362 6786
rect -2396 6684 -2362 6718
rect -2396 6616 -2362 6650
rect -2396 6548 -2362 6582
rect -2396 6480 -2362 6514
rect -2396 6412 -2362 6446
rect -2396 6344 -2362 6378
rect -2396 6276 -2362 6310
rect -2396 6208 -2362 6242
rect -2396 6140 -2362 6174
rect -2396 6072 -2362 6106
rect -2396 6004 -2362 6038
rect -2396 5936 -2362 5970
rect -2396 5868 -2362 5902
rect -2396 5800 -2362 5834
rect -2396 5732 -2362 5766
rect -2396 5664 -2362 5698
rect -2396 5596 -2362 5630
rect -2396 5528 -2362 5562
rect -2396 5460 -2362 5494
rect -2396 5392 -2362 5426
rect -2396 5324 -2362 5358
rect -2396 5256 -2362 5290
rect -2396 5188 -2362 5222
rect -2396 5120 -2362 5154
rect -2396 5052 -2362 5086
rect -2396 4984 -2362 5018
rect -2396 4916 -2362 4950
rect -2396 4848 -2362 4882
rect -2396 4780 -2362 4814
rect -2396 4712 -2362 4746
rect -2396 4644 -2362 4678
rect -2396 4576 -2362 4610
rect -2396 4508 -2362 4542
rect -2396 4440 -2362 4474
rect -2396 4372 -2362 4406
rect -2396 4304 -2362 4338
rect -2396 4236 -2362 4270
rect -2396 4168 -2362 4202
rect -2396 4100 -2362 4134
rect -2396 4032 -2362 4066
rect -2396 3964 -2362 3998
rect -2396 3896 -2362 3930
rect -2396 3828 -2362 3862
rect -2396 3760 -2362 3794
rect -2396 3692 -2362 3726
rect 47196 19400 47230 19434
rect 47196 19332 47230 19366
rect 47196 19264 47230 19298
rect 47196 19196 47230 19230
rect 47196 19128 47230 19162
rect 47196 19060 47230 19094
rect 47196 18992 47230 19026
rect 47196 18924 47230 18958
rect 47196 18856 47230 18890
rect 47196 18788 47230 18822
rect 47196 18720 47230 18754
rect 47196 18652 47230 18686
rect 47196 18584 47230 18618
rect 47196 18516 47230 18550
rect 47196 18448 47230 18482
rect 47196 18380 47230 18414
rect 47196 18312 47230 18346
rect 47196 18244 47230 18278
rect 47196 18176 47230 18210
rect 47196 18108 47230 18142
rect 47196 18040 47230 18074
rect 47196 17972 47230 18006
rect 47196 17904 47230 17938
rect 47196 17836 47230 17870
rect 47196 17768 47230 17802
rect 47196 17700 47230 17734
rect 47196 17632 47230 17666
rect 47196 17564 47230 17598
rect 47196 17496 47230 17530
rect 47196 17428 47230 17462
rect 47196 17360 47230 17394
rect 47196 17292 47230 17326
rect 47196 17224 47230 17258
rect 47196 17156 47230 17190
rect 47196 17088 47230 17122
rect 47196 17020 47230 17054
rect 47196 16952 47230 16986
rect 47196 16884 47230 16918
rect 47196 16816 47230 16850
rect 47196 16748 47230 16782
rect 47196 16680 47230 16714
rect 47196 16612 47230 16646
rect 47196 16544 47230 16578
rect 47196 16476 47230 16510
rect 47196 16408 47230 16442
rect 47196 16340 47230 16374
rect 47196 16272 47230 16306
rect 47196 16204 47230 16238
rect 47196 16136 47230 16170
rect 47196 16068 47230 16102
rect 47196 16000 47230 16034
rect 47196 15932 47230 15966
rect 47196 15864 47230 15898
rect 47196 15796 47230 15830
rect 47196 15728 47230 15762
rect 47196 15660 47230 15694
rect 47196 15592 47230 15626
rect 47196 15524 47230 15558
rect 47196 15456 47230 15490
rect 47196 15388 47230 15422
rect 47196 15320 47230 15354
rect 47196 15252 47230 15286
rect 47196 15184 47230 15218
rect 47196 15116 47230 15150
rect 47196 15048 47230 15082
rect 47196 14980 47230 15014
rect 47196 14912 47230 14946
rect 47196 14844 47230 14878
rect 47196 14776 47230 14810
rect 47196 14708 47230 14742
rect 47196 14640 47230 14674
rect 47196 14572 47230 14606
rect 47196 14504 47230 14538
rect 47196 14436 47230 14470
rect 47196 14368 47230 14402
rect 47196 14300 47230 14334
rect 47196 14232 47230 14266
rect 47196 14164 47230 14198
rect 47196 14096 47230 14130
rect 47196 14028 47230 14062
rect 47196 13960 47230 13994
rect 47196 13892 47230 13926
rect 47196 13824 47230 13858
rect 47196 13756 47230 13790
rect 47196 13688 47230 13722
rect 47196 13620 47230 13654
rect 47196 13552 47230 13586
rect 47196 13484 47230 13518
rect 47196 13416 47230 13450
rect 47196 13348 47230 13382
rect 47196 13280 47230 13314
rect 47196 13212 47230 13246
rect 47196 13144 47230 13178
rect 47196 13076 47230 13110
rect 47196 13008 47230 13042
rect 47196 12940 47230 12974
rect 47196 12872 47230 12906
rect 47196 12804 47230 12838
rect 47196 12736 47230 12770
rect 47196 12668 47230 12702
rect 47196 12600 47230 12634
rect 47196 12532 47230 12566
rect 47196 12464 47230 12498
rect 47196 12396 47230 12430
rect 47196 12328 47230 12362
rect 47196 12260 47230 12294
rect 47196 12192 47230 12226
rect 47196 12124 47230 12158
rect 47196 12056 47230 12090
rect 47196 11988 47230 12022
rect 47196 11920 47230 11954
rect 47196 11852 47230 11886
rect 47196 11784 47230 11818
rect 47196 11716 47230 11750
rect 47196 11648 47230 11682
rect 47196 11580 47230 11614
rect 47196 11512 47230 11546
rect 47196 11444 47230 11478
rect 47196 11376 47230 11410
rect 47196 11308 47230 11342
rect 47196 11240 47230 11274
rect 47196 11172 47230 11206
rect 47196 11104 47230 11138
rect 47196 11036 47230 11070
rect 47196 10968 47230 11002
rect 47196 10900 47230 10934
rect 47196 10832 47230 10866
rect 47196 10764 47230 10798
rect 47196 10696 47230 10730
rect 47196 10628 47230 10662
rect 47196 10560 47230 10594
rect 47196 10492 47230 10526
rect 47196 10424 47230 10458
rect 47196 10356 47230 10390
rect 47196 10288 47230 10322
rect 47196 10220 47230 10254
rect 47196 10152 47230 10186
rect 47196 10084 47230 10118
rect 47196 10016 47230 10050
rect 47196 9948 47230 9982
rect 47196 9880 47230 9914
rect 47196 9812 47230 9846
rect 47196 9744 47230 9778
rect 47196 9676 47230 9710
rect 47196 9608 47230 9642
rect 47196 9540 47230 9574
rect 47196 9472 47230 9506
rect 47196 9404 47230 9438
rect 47196 9336 47230 9370
rect 47196 9268 47230 9302
rect 47196 9200 47230 9234
rect 47196 9132 47230 9166
rect 47196 9064 47230 9098
rect 47196 8996 47230 9030
rect 47196 8928 47230 8962
rect 47196 8860 47230 8894
rect 47196 8792 47230 8826
rect 47196 8724 47230 8758
rect 47196 8656 47230 8690
rect 47196 8588 47230 8622
rect 47196 8520 47230 8554
rect 47196 8452 47230 8486
rect 47196 8384 47230 8418
rect 47196 8316 47230 8350
rect 47196 8248 47230 8282
rect 47196 8180 47230 8214
rect 47196 8112 47230 8146
rect 47196 8044 47230 8078
rect 47196 7976 47230 8010
rect 47196 7908 47230 7942
rect 47196 7840 47230 7874
rect 47196 7772 47230 7806
rect 47196 7704 47230 7738
rect 47196 7636 47230 7670
rect 47196 7568 47230 7602
rect 47196 7500 47230 7534
rect 47196 7432 47230 7466
rect 47196 7364 47230 7398
rect 47196 7296 47230 7330
rect 47196 7228 47230 7262
rect 47196 7160 47230 7194
rect 47196 7092 47230 7126
rect 47196 7024 47230 7058
rect 47196 6956 47230 6990
rect 47196 6888 47230 6922
rect 47196 6820 47230 6854
rect 47196 6752 47230 6786
rect 47196 6684 47230 6718
rect 47196 6616 47230 6650
rect 47196 6548 47230 6582
rect 47196 6480 47230 6514
rect 47196 6412 47230 6446
rect 47196 6344 47230 6378
rect 47196 6276 47230 6310
rect 47196 6208 47230 6242
rect 47196 6140 47230 6174
rect 47196 6072 47230 6106
rect 47196 6004 47230 6038
rect 47196 5936 47230 5970
rect 47196 5868 47230 5902
rect 47196 5800 47230 5834
rect 47196 5732 47230 5766
rect 47196 5664 47230 5698
rect 47196 5596 47230 5630
rect 47196 5528 47230 5562
rect 47196 5460 47230 5494
rect 47196 5392 47230 5426
rect 47196 5324 47230 5358
rect 47196 5256 47230 5290
rect 47196 5188 47230 5222
rect 47196 5120 47230 5154
rect 47196 5052 47230 5086
rect 47196 4984 47230 5018
rect 47196 4916 47230 4950
rect 47196 4848 47230 4882
rect 47196 4780 47230 4814
rect 47196 4712 47230 4746
rect 47196 4644 47230 4678
rect 47196 4576 47230 4610
rect 47196 4508 47230 4542
rect 47196 4440 47230 4474
rect 47196 4372 47230 4406
rect 47196 4304 47230 4338
rect 47196 4236 47230 4270
rect 47196 4168 47230 4202
rect 47196 4100 47230 4134
rect 47196 4032 47230 4066
rect 47196 3964 47230 3998
rect 47196 3896 47230 3930
rect 47196 3828 47230 3862
rect 47196 3760 47230 3794
rect 47196 3692 47230 3726
rect -2318 3606 -2284 3640
rect -2250 3606 -2216 3640
rect -2182 3606 -2148 3640
rect -2114 3606 -2080 3640
rect -2046 3606 -2012 3640
rect -1978 3606 -1944 3640
rect -1910 3606 -1876 3640
rect -1842 3606 -1808 3640
rect -1774 3606 -1740 3640
rect -1706 3606 -1672 3640
rect -1638 3606 -1604 3640
rect -1570 3606 -1536 3640
rect -1502 3606 -1468 3640
rect -1434 3606 -1400 3640
rect -1366 3606 -1332 3640
rect -1298 3606 -1264 3640
rect -1230 3606 -1196 3640
rect -1162 3606 -1128 3640
rect -1094 3606 -1060 3640
rect -1026 3606 -992 3640
rect -958 3606 -924 3640
rect -890 3606 -856 3640
rect -822 3606 -788 3640
rect -754 3606 -720 3640
rect -686 3606 -652 3640
rect -618 3606 -584 3640
rect -550 3606 -516 3640
rect -482 3606 -448 3640
rect -414 3606 -380 3640
rect -346 3606 -312 3640
rect -278 3606 -244 3640
rect -210 3606 -176 3640
rect -142 3606 -108 3640
rect -74 3606 -40 3640
rect -6 3606 28 3640
rect 62 3606 96 3640
rect 130 3606 164 3640
rect 198 3606 232 3640
rect 266 3606 300 3640
rect 334 3606 368 3640
rect 402 3606 436 3640
rect 470 3606 504 3640
rect 538 3606 572 3640
rect 606 3606 640 3640
rect 674 3606 708 3640
rect 742 3606 776 3640
rect 810 3606 844 3640
rect 878 3606 912 3640
rect 946 3606 980 3640
rect 1014 3606 1048 3640
rect 1082 3606 1116 3640
rect 1150 3606 1184 3640
rect 1218 3606 1252 3640
rect 1286 3606 1320 3640
rect 1354 3606 1388 3640
rect 1422 3606 1456 3640
rect 1490 3606 1524 3640
rect 1558 3606 1592 3640
rect 1626 3606 1660 3640
rect 1694 3606 1728 3640
rect 1762 3606 1796 3640
rect 1830 3606 1864 3640
rect 1898 3606 1932 3640
rect 1966 3606 2000 3640
rect 2034 3606 2068 3640
rect 2102 3606 2136 3640
rect 2170 3606 2204 3640
rect 2238 3606 2272 3640
rect 2306 3606 2340 3640
rect 2374 3606 2408 3640
rect 2442 3606 2476 3640
rect 2510 3606 2544 3640
rect 2578 3606 2612 3640
rect 2646 3606 2680 3640
rect 2714 3606 2748 3640
rect 2782 3606 2816 3640
rect 2850 3606 2884 3640
rect 2918 3606 2952 3640
rect 2986 3606 3020 3640
rect 3054 3606 3088 3640
rect 3122 3606 3156 3640
rect 3190 3606 3224 3640
rect 3258 3606 3292 3640
rect 3326 3606 3360 3640
rect 3394 3606 3428 3640
rect 3462 3606 3496 3640
rect 3530 3606 3564 3640
rect 3598 3606 3632 3640
rect 3666 3606 3700 3640
rect 3734 3606 3768 3640
rect 3802 3606 3836 3640
rect 3870 3606 3904 3640
rect 3938 3606 3972 3640
rect 4006 3606 4040 3640
rect 4074 3606 4108 3640
rect 4142 3606 4176 3640
rect 4210 3606 4244 3640
rect 4278 3606 4312 3640
rect 4346 3606 4380 3640
rect 4414 3606 4448 3640
rect 4482 3606 4516 3640
rect 4550 3606 4584 3640
rect 4618 3606 4652 3640
rect 4686 3606 4720 3640
rect 4754 3606 4788 3640
rect 4822 3606 4856 3640
rect 4890 3606 4924 3640
rect 4958 3606 4992 3640
rect 5026 3606 5060 3640
rect 5094 3606 5128 3640
rect 5162 3606 5196 3640
rect 5230 3606 5264 3640
rect 5298 3606 5332 3640
rect 5366 3606 5400 3640
rect 5434 3606 5468 3640
rect 5502 3606 5536 3640
rect 5570 3606 5604 3640
rect 5638 3606 5672 3640
rect 5706 3606 5740 3640
rect 5774 3606 5808 3640
rect 5842 3606 5876 3640
rect 5910 3606 5944 3640
rect 5978 3606 6012 3640
rect 6046 3606 6080 3640
rect 6114 3606 6148 3640
rect 6182 3606 6216 3640
rect 6250 3606 6284 3640
rect 6318 3606 6352 3640
rect 6386 3606 6420 3640
rect 6454 3606 6488 3640
rect 6522 3606 6556 3640
rect 6590 3606 6624 3640
rect 6658 3606 6692 3640
rect 6726 3606 6760 3640
rect 6794 3606 6828 3640
rect 6862 3606 6896 3640
rect 6930 3606 6964 3640
rect 6998 3606 7032 3640
rect 7066 3606 7100 3640
rect 7134 3606 7168 3640
rect 7202 3606 7236 3640
rect 7270 3606 7304 3640
rect 7338 3606 7372 3640
rect 7406 3606 7440 3640
rect 7474 3606 7508 3640
rect 7542 3606 7576 3640
rect 7610 3606 7644 3640
rect 7678 3606 7712 3640
rect 7746 3606 7780 3640
rect 7814 3606 7848 3640
rect 7882 3606 7916 3640
rect 7950 3606 7984 3640
rect 8018 3606 8052 3640
rect 8086 3606 8120 3640
rect 8154 3606 8188 3640
rect 8222 3606 8256 3640
rect 8290 3606 8324 3640
rect 8358 3606 8392 3640
rect 8426 3606 8460 3640
rect 8494 3606 8528 3640
rect 8562 3606 8596 3640
rect 8630 3606 8664 3640
rect 8698 3606 8732 3640
rect 8766 3606 8800 3640
rect 8834 3606 8868 3640
rect 8902 3606 8936 3640
rect 8970 3606 9004 3640
rect 9038 3606 9072 3640
rect 9106 3606 9140 3640
rect 9174 3606 9208 3640
rect 9242 3606 9276 3640
rect 9310 3606 9344 3640
rect 9378 3606 9412 3640
rect 9446 3606 9480 3640
rect 9514 3606 9548 3640
rect 9582 3606 9616 3640
rect 9650 3606 9684 3640
rect 9718 3606 9752 3640
rect 9786 3606 9820 3640
rect 9854 3606 9888 3640
rect 9922 3606 9956 3640
rect 9990 3606 10024 3640
rect 10058 3606 10092 3640
rect 10126 3606 10160 3640
rect 10194 3606 10228 3640
rect 10262 3606 10296 3640
rect 10330 3606 10364 3640
rect 10398 3606 10432 3640
rect 10466 3606 10500 3640
rect 10534 3606 10568 3640
rect 10602 3606 10636 3640
rect 10670 3606 10704 3640
rect 10738 3606 10772 3640
rect 10806 3606 10840 3640
rect 10874 3606 10908 3640
rect 10942 3606 10976 3640
rect 11010 3606 11044 3640
rect 11078 3606 11112 3640
rect 11146 3606 11180 3640
rect 11214 3606 11248 3640
rect 11282 3606 11316 3640
rect 11350 3606 11384 3640
rect 11418 3606 11452 3640
rect 11486 3606 11520 3640
rect 11554 3606 11588 3640
rect 11622 3606 11656 3640
rect 11690 3606 11724 3640
rect 11758 3606 11792 3640
rect 11826 3606 11860 3640
rect 11894 3606 11928 3640
rect 11962 3606 11996 3640
rect 12030 3606 12064 3640
rect 12098 3606 12132 3640
rect 12166 3606 12200 3640
rect 12234 3606 12268 3640
rect 12302 3606 12336 3640
rect 12370 3606 12404 3640
rect 12438 3606 12472 3640
rect 12506 3606 12540 3640
rect 12574 3606 12608 3640
rect 12642 3606 12676 3640
rect 12710 3606 12744 3640
rect 12778 3606 12812 3640
rect 12846 3606 12880 3640
rect 12914 3606 12948 3640
rect 12982 3606 13016 3640
rect 13050 3606 13084 3640
rect 13118 3606 13152 3640
rect 13186 3606 13220 3640
rect 13254 3606 13288 3640
rect 13322 3606 13356 3640
rect 13390 3606 13424 3640
rect 13458 3606 13492 3640
rect 13526 3606 13560 3640
rect 13594 3606 13628 3640
rect 13662 3606 13696 3640
rect 13730 3606 13764 3640
rect 13798 3606 13832 3640
rect 13866 3606 13900 3640
rect 13934 3606 13968 3640
rect 14002 3606 14036 3640
rect 14070 3606 14104 3640
rect 14138 3606 14172 3640
rect 14206 3606 14240 3640
rect 14274 3606 14308 3640
rect 14342 3606 14376 3640
rect 14410 3606 14444 3640
rect 14478 3606 14512 3640
rect 14546 3606 14580 3640
rect 14614 3606 14648 3640
rect 14682 3606 14716 3640
rect 14750 3606 14784 3640
rect 14818 3606 14852 3640
rect 14886 3606 14920 3640
rect 14954 3606 14988 3640
rect 15022 3606 15056 3640
rect 15090 3606 15124 3640
rect 15158 3606 15192 3640
rect 15226 3606 15260 3640
rect 15294 3606 15328 3640
rect 15362 3606 15396 3640
rect 15430 3606 15464 3640
rect 15498 3606 15532 3640
rect 15566 3606 15600 3640
rect 15634 3606 15668 3640
rect 15702 3606 15736 3640
rect 15770 3606 15804 3640
rect 15838 3606 15872 3640
rect 15906 3606 15940 3640
rect 15974 3606 16008 3640
rect 16042 3606 16076 3640
rect 16110 3606 16144 3640
rect 16178 3606 16212 3640
rect 16246 3606 16280 3640
rect 16314 3606 16348 3640
rect 16382 3606 16416 3640
rect 16450 3606 16484 3640
rect 16518 3606 16552 3640
rect 16586 3606 16620 3640
rect 16654 3606 16688 3640
rect 16722 3606 16756 3640
rect 16790 3606 16824 3640
rect 16858 3606 16892 3640
rect 16926 3606 16960 3640
rect 16994 3606 17028 3640
rect 17062 3606 17096 3640
rect 17130 3606 17164 3640
rect 17198 3606 17232 3640
rect 17266 3606 17300 3640
rect 17334 3606 17368 3640
rect 17402 3606 17436 3640
rect 17470 3606 17504 3640
rect 17538 3606 17572 3640
rect 17606 3606 17640 3640
rect 17674 3606 17708 3640
rect 17742 3606 17776 3640
rect 17810 3606 17844 3640
rect 17878 3606 17912 3640
rect 17946 3606 17980 3640
rect 18014 3606 18048 3640
rect 18082 3606 18116 3640
rect 18150 3606 18184 3640
rect 18218 3606 18252 3640
rect 18286 3606 18320 3640
rect 18354 3606 18388 3640
rect 18422 3606 18456 3640
rect 18490 3606 18524 3640
rect 18558 3606 18592 3640
rect 18626 3606 18660 3640
rect 18694 3606 18728 3640
rect 18762 3606 18796 3640
rect 18830 3606 18864 3640
rect 18898 3606 18932 3640
rect 18966 3606 19000 3640
rect 19034 3606 19068 3640
rect 19102 3606 19136 3640
rect 19170 3606 19204 3640
rect 19238 3606 19272 3640
rect 19306 3606 19340 3640
rect 19374 3606 19408 3640
rect 19442 3606 19476 3640
rect 19510 3606 19544 3640
rect 19578 3606 19612 3640
rect 19646 3606 19680 3640
rect 19714 3606 19748 3640
rect 19782 3606 19816 3640
rect 19850 3606 19884 3640
rect 19918 3606 19952 3640
rect 19986 3606 20020 3640
rect 20054 3606 20088 3640
rect 20122 3606 20156 3640
rect 20190 3606 20224 3640
rect 20258 3606 20292 3640
rect 20326 3606 20360 3640
rect 20394 3606 20428 3640
rect 20462 3606 20496 3640
rect 20530 3606 20564 3640
rect 20598 3606 20632 3640
rect 20666 3606 20700 3640
rect 20734 3606 20768 3640
rect 20802 3606 20836 3640
rect 20870 3606 20904 3640
rect 20938 3606 20972 3640
rect 21006 3606 21040 3640
rect 21074 3606 21108 3640
rect 21142 3606 21176 3640
rect 21210 3606 21244 3640
rect 21278 3606 21312 3640
rect 21346 3606 21380 3640
rect 21414 3606 21448 3640
rect 21482 3606 21516 3640
rect 21550 3606 21584 3640
rect 21618 3606 21652 3640
rect 21686 3606 21720 3640
rect 21754 3606 21788 3640
rect 21822 3606 21856 3640
rect 21890 3606 21924 3640
rect 21958 3606 21992 3640
rect 22026 3606 22060 3640
rect 22094 3606 22128 3640
rect 22162 3606 22196 3640
rect 22230 3606 22264 3640
rect 22298 3606 22332 3640
rect 22366 3606 22400 3640
rect 22434 3606 22468 3640
rect 22502 3606 22536 3640
rect 22570 3606 22604 3640
rect 22638 3606 22672 3640
rect 22706 3606 22740 3640
rect 22774 3606 22808 3640
rect 22842 3606 22876 3640
rect 22910 3606 22944 3640
rect 22978 3606 23012 3640
rect 23046 3606 23080 3640
rect 23114 3606 23148 3640
rect 23182 3606 23216 3640
rect 23250 3606 23284 3640
rect 23318 3606 23352 3640
rect 23386 3606 23420 3640
rect 23454 3606 23488 3640
rect 23522 3606 23556 3640
rect 23590 3606 23624 3640
rect 23658 3606 23692 3640
rect 23726 3606 23760 3640
rect 23794 3606 23828 3640
rect 23862 3606 23896 3640
rect 23930 3606 23964 3640
rect 23998 3606 24032 3640
rect 24066 3606 24100 3640
rect 24134 3606 24168 3640
rect 24202 3606 24236 3640
rect 24270 3606 24304 3640
rect 24338 3606 24372 3640
rect 24406 3606 24440 3640
rect 24474 3606 24508 3640
rect 24542 3606 24576 3640
rect 24610 3606 24644 3640
rect 24678 3606 24712 3640
rect 24746 3606 24780 3640
rect 24814 3606 24848 3640
rect 24882 3606 24916 3640
rect 24950 3606 24984 3640
rect 25018 3606 25052 3640
rect 25086 3606 25120 3640
rect 25154 3606 25188 3640
rect 25222 3606 25256 3640
rect 25290 3606 25324 3640
rect 25358 3606 25392 3640
rect 25426 3606 25460 3640
rect 25494 3606 25528 3640
rect 25562 3606 25596 3640
rect 25630 3606 25664 3640
rect 25698 3606 25732 3640
rect 25766 3606 25800 3640
rect 25834 3606 25868 3640
rect 25902 3606 25936 3640
rect 25970 3606 26004 3640
rect 26038 3606 26072 3640
rect 26106 3606 26140 3640
rect 26174 3606 26208 3640
rect 26242 3606 26276 3640
rect 26310 3606 26344 3640
rect 26378 3606 26412 3640
rect 26446 3606 26480 3640
rect 26514 3606 26548 3640
rect 26582 3606 26616 3640
rect 26650 3606 26684 3640
rect 26718 3606 26752 3640
rect 26786 3606 26820 3640
rect 26854 3606 26888 3640
rect 26922 3606 26956 3640
rect 26990 3606 27024 3640
rect 27058 3606 27092 3640
rect 27126 3606 27160 3640
rect 27194 3606 27228 3640
rect 27262 3606 27296 3640
rect 27330 3606 27364 3640
rect 27398 3606 27432 3640
rect 27466 3606 27500 3640
rect 27534 3606 27568 3640
rect 27602 3606 27636 3640
rect 27670 3606 27704 3640
rect 27738 3606 27772 3640
rect 27806 3606 27840 3640
rect 27874 3606 27908 3640
rect 27942 3606 27976 3640
rect 28010 3606 28044 3640
rect 28078 3606 28112 3640
rect 28146 3606 28180 3640
rect 28214 3606 28248 3640
rect 28282 3606 28316 3640
rect 28350 3606 28384 3640
rect 28418 3606 28452 3640
rect 28486 3606 28520 3640
rect 28554 3606 28588 3640
rect 28622 3606 28656 3640
rect 28690 3606 28724 3640
rect 28758 3606 28792 3640
rect 28826 3606 28860 3640
rect 28894 3606 28928 3640
rect 28962 3606 28996 3640
rect 29030 3606 29064 3640
rect 29098 3606 29132 3640
rect 29166 3606 29200 3640
rect 29234 3606 29268 3640
rect 29302 3606 29336 3640
rect 29370 3606 29404 3640
rect 29438 3606 29472 3640
rect 29506 3606 29540 3640
rect 29574 3606 29608 3640
rect 29642 3606 29676 3640
rect 29710 3606 29744 3640
rect 29778 3606 29812 3640
rect 29846 3606 29880 3640
rect 29914 3606 29948 3640
rect 29982 3606 30016 3640
rect 30050 3606 30084 3640
rect 30118 3606 30152 3640
rect 30186 3606 30220 3640
rect 30254 3606 30288 3640
rect 30322 3606 30356 3640
rect 30390 3606 30424 3640
rect 30458 3606 30492 3640
rect 30526 3606 30560 3640
rect 30594 3606 30628 3640
rect 30662 3606 30696 3640
rect 30730 3606 30764 3640
rect 30798 3606 30832 3640
rect 30866 3606 30900 3640
rect 30934 3606 30968 3640
rect 31002 3606 31036 3640
rect 31070 3606 31104 3640
rect 31138 3606 31172 3640
rect 31206 3606 31240 3640
rect 31274 3606 31308 3640
rect 31342 3606 31376 3640
rect 31410 3606 31444 3640
rect 31478 3606 31512 3640
rect 31546 3606 31580 3640
rect 31614 3606 31648 3640
rect 31682 3606 31716 3640
rect 31750 3606 31784 3640
rect 31818 3606 31852 3640
rect 31886 3606 31920 3640
rect 31954 3606 31988 3640
rect 32022 3606 32056 3640
rect 32090 3606 32124 3640
rect 32158 3606 32192 3640
rect 32226 3606 32260 3640
rect 32294 3606 32328 3640
rect 32362 3606 32396 3640
rect 32430 3606 32464 3640
rect 32498 3606 32532 3640
rect 32566 3606 32600 3640
rect 32634 3606 32668 3640
rect 32702 3606 32736 3640
rect 32770 3606 32804 3640
rect 32838 3606 32872 3640
rect 32906 3606 32940 3640
rect 32974 3606 33008 3640
rect 33042 3606 33076 3640
rect 33110 3606 33144 3640
rect 33178 3606 33212 3640
rect 33246 3606 33280 3640
rect 33314 3606 33348 3640
rect 33382 3606 33416 3640
rect 33450 3606 33484 3640
rect 33518 3606 33552 3640
rect 33586 3606 33620 3640
rect 33654 3606 33688 3640
rect 33722 3606 33756 3640
rect 33790 3606 33824 3640
rect 33858 3606 33892 3640
rect 33926 3606 33960 3640
rect 33994 3606 34028 3640
rect 34062 3606 34096 3640
rect 34130 3606 34164 3640
rect 34198 3606 34232 3640
rect 34266 3606 34300 3640
rect 34334 3606 34368 3640
rect 34402 3606 34436 3640
rect 34470 3606 34504 3640
rect 34538 3606 34572 3640
rect 34606 3606 34640 3640
rect 34674 3606 34708 3640
rect 34742 3606 34776 3640
rect 34810 3606 34844 3640
rect 34878 3606 34912 3640
rect 34946 3606 34980 3640
rect 35014 3606 35048 3640
rect 35082 3606 35116 3640
rect 35150 3606 35184 3640
rect 35218 3606 35252 3640
rect 35286 3606 35320 3640
rect 35354 3606 35388 3640
rect 35422 3606 35456 3640
rect 35490 3606 35524 3640
rect 35558 3606 35592 3640
rect 35626 3606 35660 3640
rect 35694 3606 35728 3640
rect 35762 3606 35796 3640
rect 35830 3606 35864 3640
rect 35898 3606 35932 3640
rect 35966 3606 36000 3640
rect 36034 3606 36068 3640
rect 36102 3606 36136 3640
rect 36170 3606 36204 3640
rect 36238 3606 36272 3640
rect 36306 3606 36340 3640
rect 36374 3606 36408 3640
rect 36442 3606 36476 3640
rect 36510 3606 36544 3640
rect 36578 3606 36612 3640
rect 36646 3606 36680 3640
rect 36714 3606 36748 3640
rect 36782 3606 36816 3640
rect 36850 3606 36884 3640
rect 36918 3606 36952 3640
rect 36986 3606 37020 3640
rect 37054 3606 37088 3640
rect 37122 3606 37156 3640
rect 37190 3606 37224 3640
rect 37258 3606 37292 3640
rect 37326 3606 37360 3640
rect 37394 3606 37428 3640
rect 37462 3606 37496 3640
rect 37530 3606 37564 3640
rect 37598 3606 37632 3640
rect 37666 3606 37700 3640
rect 37734 3606 37768 3640
rect 37802 3606 37836 3640
rect 37870 3606 37904 3640
rect 37938 3606 37972 3640
rect 38006 3606 38040 3640
rect 38074 3606 38108 3640
rect 38142 3606 38176 3640
rect 38210 3606 38244 3640
rect 38278 3606 38312 3640
rect 38346 3606 38380 3640
rect 38414 3606 38448 3640
rect 38482 3606 38516 3640
rect 38550 3606 38584 3640
rect 38618 3606 38652 3640
rect 38686 3606 38720 3640
rect 38754 3606 38788 3640
rect 38822 3606 38856 3640
rect 38890 3606 38924 3640
rect 38958 3606 38992 3640
rect 39026 3606 39060 3640
rect 39094 3606 39128 3640
rect 39162 3606 39196 3640
rect 39230 3606 39264 3640
rect 39298 3606 39332 3640
rect 39366 3606 39400 3640
rect 39434 3606 39468 3640
rect 39502 3606 39536 3640
rect 39570 3606 39604 3640
rect 39638 3606 39672 3640
rect 39706 3606 39740 3640
rect 39774 3606 39808 3640
rect 39842 3606 39876 3640
rect 39910 3606 39944 3640
rect 39978 3606 40012 3640
rect 40046 3606 40080 3640
rect 40114 3606 40148 3640
rect 40182 3606 40216 3640
rect 40250 3606 40284 3640
rect 40318 3606 40352 3640
rect 40386 3606 40420 3640
rect 40454 3606 40488 3640
rect 40522 3606 40556 3640
rect 40590 3606 40624 3640
rect 40658 3606 40692 3640
rect 40726 3606 40760 3640
rect 40794 3606 40828 3640
rect 40862 3606 40896 3640
rect 40930 3606 40964 3640
rect 40998 3606 41032 3640
rect 41066 3606 41100 3640
rect 41134 3606 41168 3640
rect 41202 3606 41236 3640
rect 41270 3606 41304 3640
rect 41338 3606 41372 3640
rect 41406 3606 41440 3640
rect 41474 3606 41508 3640
rect 41542 3606 41576 3640
rect 41610 3606 41644 3640
rect 41678 3606 41712 3640
rect 41746 3606 41780 3640
rect 41814 3606 41848 3640
rect 41882 3606 41916 3640
rect 41950 3606 41984 3640
rect 42018 3606 42052 3640
rect 42086 3606 42120 3640
rect 42154 3606 42188 3640
rect 42222 3606 42256 3640
rect 42290 3606 42324 3640
rect 42358 3606 42392 3640
rect 42426 3606 42460 3640
rect 42494 3606 42528 3640
rect 42562 3606 42596 3640
rect 42630 3606 42664 3640
rect 42698 3606 42732 3640
rect 42766 3606 42800 3640
rect 42834 3606 42868 3640
rect 42902 3606 42936 3640
rect 42970 3606 43004 3640
rect 43038 3606 43072 3640
rect 43106 3606 43140 3640
rect 43174 3606 43208 3640
rect 43242 3606 43276 3640
rect 43310 3606 43344 3640
rect 43378 3606 43412 3640
rect 43446 3606 43480 3640
rect 43514 3606 43548 3640
rect 43582 3606 43616 3640
rect 43650 3606 43684 3640
rect 43718 3606 43752 3640
rect 43786 3606 43820 3640
rect 43854 3606 43888 3640
rect 43922 3606 43956 3640
rect 43990 3606 44024 3640
rect 44058 3606 44092 3640
rect 44126 3606 44160 3640
rect 44194 3606 44228 3640
rect 44262 3606 44296 3640
rect 44330 3606 44364 3640
rect 44398 3606 44432 3640
rect 44466 3606 44500 3640
rect 44534 3606 44568 3640
rect 44602 3606 44636 3640
rect 44670 3606 44704 3640
rect 44738 3606 44772 3640
rect 44806 3606 44840 3640
rect 44874 3606 44908 3640
rect 44942 3606 44976 3640
rect 45010 3606 45044 3640
rect 45078 3606 45112 3640
rect 45146 3606 45180 3640
rect 45214 3606 45248 3640
rect 45282 3606 45316 3640
rect 45350 3606 45384 3640
rect 45418 3606 45452 3640
rect 45486 3606 45520 3640
rect 45554 3606 45588 3640
rect 45622 3606 45656 3640
rect 45690 3606 45724 3640
rect 45758 3606 45792 3640
rect 45826 3606 45860 3640
rect 45894 3606 45928 3640
rect 45962 3606 45996 3640
rect 46030 3606 46064 3640
rect 46098 3606 46132 3640
rect 46166 3606 46200 3640
rect 46234 3606 46268 3640
rect 46302 3606 46336 3640
rect 46370 3606 46404 3640
rect 46438 3606 46472 3640
rect 46506 3606 46540 3640
rect 46574 3606 46608 3640
rect 46642 3606 46676 3640
rect 46710 3606 46744 3640
rect 46778 3606 46812 3640
rect 46846 3606 46880 3640
rect 46914 3606 46948 3640
rect 46982 3606 47016 3640
rect 47050 3606 47084 3640
rect 47118 3606 47152 3640
<< locali >>
rect -2396 116750 -2318 116784
rect -2284 116750 -2250 116784
rect -2216 116750 -2182 116784
rect -2148 116750 -2114 116784
rect -2080 116750 -2046 116784
rect -2012 116750 -1978 116784
rect -1944 116750 -1910 116784
rect -1876 116750 -1842 116784
rect -1808 116750 -1774 116784
rect -1740 116750 -1706 116784
rect -1672 116750 -1638 116784
rect -1604 116750 -1570 116784
rect -1536 116750 -1502 116784
rect -1468 116750 -1434 116784
rect -1400 116750 -1366 116784
rect -1332 116750 -1298 116784
rect -1264 116750 -1230 116784
rect -1196 116750 -1162 116784
rect -1128 116750 -1094 116784
rect -1060 116750 -1026 116784
rect -992 116750 -958 116784
rect -924 116750 -890 116784
rect -856 116750 -822 116784
rect -788 116750 -754 116784
rect -720 116750 -686 116784
rect -652 116750 -618 116784
rect -584 116750 -550 116784
rect -516 116750 -482 116784
rect -448 116750 -414 116784
rect -380 116750 -346 116784
rect -312 116750 -278 116784
rect -244 116750 -210 116784
rect -176 116750 -142 116784
rect -108 116750 -74 116784
rect -40 116750 -6 116784
rect 28 116750 62 116784
rect 96 116750 130 116784
rect 164 116750 198 116784
rect 232 116750 266 116784
rect 300 116750 334 116784
rect 368 116750 402 116784
rect 436 116750 470 116784
rect 504 116750 538 116784
rect 572 116750 606 116784
rect 640 116750 674 116784
rect 708 116750 742 116784
rect 776 116750 810 116784
rect 844 116750 878 116784
rect 912 116750 946 116784
rect 980 116750 1014 116784
rect 1048 116750 1082 116784
rect 1116 116750 1150 116784
rect 1184 116750 1218 116784
rect 1252 116750 1286 116784
rect 1320 116750 1354 116784
rect 1388 116750 1422 116784
rect 1456 116750 1490 116784
rect 1524 116750 1558 116784
rect 1592 116750 1626 116784
rect 1660 116750 1694 116784
rect 1728 116750 1762 116784
rect 1796 116750 1830 116784
rect 1864 116750 1898 116784
rect 1932 116750 1966 116784
rect 2000 116750 2034 116784
rect 2068 116750 2102 116784
rect 2136 116750 2170 116784
rect 2204 116750 2238 116784
rect 2272 116750 2306 116784
rect 2340 116750 2374 116784
rect 2408 116750 2442 116784
rect 2476 116750 2510 116784
rect 2544 116750 2578 116784
rect 2612 116750 2646 116784
rect 2680 116750 2714 116784
rect 2748 116750 2782 116784
rect 2816 116750 2850 116784
rect 2884 116750 2918 116784
rect 2952 116750 2986 116784
rect 3020 116750 3054 116784
rect 3088 116750 3122 116784
rect 3156 116750 3190 116784
rect 3224 116750 3258 116784
rect 3292 116750 3326 116784
rect 3360 116750 3394 116784
rect 3428 116750 3462 116784
rect 3496 116750 3530 116784
rect 3564 116750 3598 116784
rect 3632 116750 3666 116784
rect 3700 116750 3734 116784
rect 3768 116750 3802 116784
rect 3836 116750 3870 116784
rect 3904 116750 3938 116784
rect 3972 116750 4006 116784
rect 4040 116750 4074 116784
rect 4108 116750 4142 116784
rect 4176 116750 4210 116784
rect 4244 116750 4278 116784
rect 4312 116750 4346 116784
rect 4380 116750 4414 116784
rect 4448 116750 4482 116784
rect 4516 116750 4550 116784
rect 4584 116750 4618 116784
rect 4652 116750 4686 116784
rect 4720 116750 4754 116784
rect 4788 116750 4822 116784
rect 4856 116750 4890 116784
rect 4924 116750 4958 116784
rect 4992 116750 5026 116784
rect 5060 116750 5094 116784
rect 5128 116750 5162 116784
rect 5196 116750 5230 116784
rect 5264 116750 5298 116784
rect 5332 116750 5366 116784
rect 5400 116750 5434 116784
rect 5468 116750 5502 116784
rect 5536 116750 5570 116784
rect 5604 116750 5638 116784
rect 5672 116750 5706 116784
rect 5740 116750 5774 116784
rect 5808 116750 5842 116784
rect 5876 116750 5910 116784
rect 5944 116750 5978 116784
rect 6012 116750 6046 116784
rect 6080 116750 6114 116784
rect 6148 116750 6182 116784
rect 6216 116750 6250 116784
rect 6284 116750 6318 116784
rect 6352 116750 6386 116784
rect 6420 116750 6454 116784
rect 6488 116750 6522 116784
rect 6556 116750 6590 116784
rect 6624 116750 6658 116784
rect 6692 116750 6726 116784
rect 6760 116750 6794 116784
rect 6828 116750 6862 116784
rect 6896 116750 6930 116784
rect 6964 116750 6998 116784
rect 7032 116750 7066 116784
rect 7100 116750 7134 116784
rect 7168 116750 7202 116784
rect 7236 116750 7270 116784
rect 7304 116750 7338 116784
rect 7372 116750 7406 116784
rect 7440 116750 7474 116784
rect 7508 116750 7542 116784
rect 7576 116750 7610 116784
rect 7644 116750 7678 116784
rect 7712 116750 7746 116784
rect 7780 116750 7814 116784
rect 7848 116750 7882 116784
rect 7916 116750 7950 116784
rect 7984 116750 8018 116784
rect 8052 116750 8086 116784
rect 8120 116750 8154 116784
rect 8188 116750 8222 116784
rect 8256 116750 8290 116784
rect 8324 116750 8358 116784
rect 8392 116750 8426 116784
rect 8460 116750 8494 116784
rect 8528 116750 8562 116784
rect 8596 116750 8630 116784
rect 8664 116750 8698 116784
rect 8732 116750 8766 116784
rect 8800 116750 8834 116784
rect 8868 116750 8902 116784
rect 8936 116750 8970 116784
rect 9004 116750 9038 116784
rect 9072 116750 9106 116784
rect 9140 116750 9174 116784
rect 9208 116750 9242 116784
rect 9276 116750 9310 116784
rect 9344 116750 9378 116784
rect 9412 116750 9446 116784
rect 9480 116750 9514 116784
rect 9548 116750 9582 116784
rect 9616 116750 9650 116784
rect 9684 116750 9718 116784
rect 9752 116750 9786 116784
rect 9820 116750 9854 116784
rect 9888 116750 9922 116784
rect 9956 116750 9990 116784
rect 10024 116750 10058 116784
rect 10092 116750 10126 116784
rect 10160 116750 10194 116784
rect 10228 116750 10262 116784
rect 10296 116750 10330 116784
rect 10364 116750 10398 116784
rect 10432 116750 10466 116784
rect 10500 116750 10534 116784
rect 10568 116750 10602 116784
rect 10636 116750 10670 116784
rect 10704 116750 10738 116784
rect 10772 116750 10806 116784
rect 10840 116750 10874 116784
rect 10908 116750 10942 116784
rect 10976 116750 11010 116784
rect 11044 116750 11078 116784
rect 11112 116750 11146 116784
rect 11180 116750 11214 116784
rect 11248 116750 11282 116784
rect 11316 116750 11350 116784
rect 11384 116750 11418 116784
rect 11452 116750 11486 116784
rect 11520 116750 11554 116784
rect 11588 116750 11622 116784
rect 11656 116750 11690 116784
rect 11724 116750 11758 116784
rect 11792 116750 11826 116784
rect 11860 116750 11894 116784
rect 11928 116750 11962 116784
rect 11996 116750 12030 116784
rect 12064 116750 12098 116784
rect 12132 116750 12166 116784
rect 12200 116750 12234 116784
rect 12268 116750 12302 116784
rect 12336 116750 12370 116784
rect 12404 116750 12438 116784
rect 12472 116750 12506 116784
rect 12540 116750 12574 116784
rect 12608 116750 12642 116784
rect 12676 116750 12710 116784
rect 12744 116750 12778 116784
rect 12812 116750 12846 116784
rect 12880 116750 12914 116784
rect 12948 116750 12982 116784
rect 13016 116750 13050 116784
rect 13084 116750 13118 116784
rect 13152 116750 13186 116784
rect 13220 116750 13254 116784
rect 13288 116750 13322 116784
rect 13356 116750 13390 116784
rect 13424 116750 13458 116784
rect 13492 116750 13526 116784
rect 13560 116750 13594 116784
rect 13628 116750 13662 116784
rect 13696 116750 13730 116784
rect 13764 116750 13798 116784
rect 13832 116750 13866 116784
rect 13900 116750 13934 116784
rect 13968 116750 14002 116784
rect 14036 116750 14070 116784
rect 14104 116750 14138 116784
rect 14172 116750 14206 116784
rect 14240 116750 14274 116784
rect 14308 116750 14342 116784
rect 14376 116750 14410 116784
rect 14444 116750 14478 116784
rect 14512 116750 14546 116784
rect 14580 116750 14614 116784
rect 14648 116750 14682 116784
rect 14716 116750 14750 116784
rect 14784 116750 14818 116784
rect 14852 116750 14886 116784
rect 14920 116750 14954 116784
rect 14988 116750 15022 116784
rect 15056 116750 15090 116784
rect 15124 116750 15158 116784
rect 15192 116750 15226 116784
rect 15260 116750 15294 116784
rect 15328 116750 15362 116784
rect 15396 116750 15430 116784
rect 15464 116750 15498 116784
rect 15532 116750 15566 116784
rect 15600 116750 15634 116784
rect 15668 116750 15702 116784
rect 15736 116750 15770 116784
rect 15804 116750 15838 116784
rect 15872 116750 15906 116784
rect 15940 116750 15974 116784
rect 16008 116750 16042 116784
rect 16076 116750 16110 116784
rect 16144 116750 16178 116784
rect 16212 116750 16246 116784
rect 16280 116750 16314 116784
rect 16348 116750 16382 116784
rect 16416 116750 16450 116784
rect 16484 116750 16518 116784
rect 16552 116750 16586 116784
rect 16620 116750 16654 116784
rect 16688 116750 16722 116784
rect 16756 116750 16790 116784
rect 16824 116750 16858 116784
rect 16892 116750 16926 116784
rect 16960 116750 16994 116784
rect 17028 116750 17062 116784
rect 17096 116750 17130 116784
rect 17164 116750 17198 116784
rect 17232 116750 17266 116784
rect 17300 116750 17334 116784
rect 17368 116750 17402 116784
rect 17436 116750 17470 116784
rect 17504 116750 17538 116784
rect 17572 116750 17606 116784
rect 17640 116750 17674 116784
rect 17708 116750 17742 116784
rect 17776 116750 17810 116784
rect 17844 116750 17878 116784
rect 17912 116750 17946 116784
rect 17980 116750 18014 116784
rect 18048 116750 18082 116784
rect 18116 116750 18150 116784
rect 18184 116750 18218 116784
rect 18252 116750 18286 116784
rect 18320 116750 18354 116784
rect 18388 116750 18422 116784
rect 18456 116750 18490 116784
rect 18524 116750 18558 116784
rect 18592 116750 18626 116784
rect 18660 116750 18694 116784
rect 18728 116750 18762 116784
rect 18796 116750 18830 116784
rect 18864 116750 18898 116784
rect 18932 116750 18966 116784
rect 19000 116750 19034 116784
rect 19068 116750 19102 116784
rect 19136 116750 19170 116784
rect 19204 116750 19238 116784
rect 19272 116750 19306 116784
rect 19340 116750 19374 116784
rect 19408 116750 19442 116784
rect 19476 116750 19510 116784
rect 19544 116750 19578 116784
rect 19612 116750 19646 116784
rect 19680 116750 19714 116784
rect 19748 116750 19782 116784
rect 19816 116750 19850 116784
rect 19884 116750 19918 116784
rect 19952 116750 19986 116784
rect 20020 116750 20054 116784
rect 20088 116750 20122 116784
rect 20156 116750 20190 116784
rect 20224 116750 20258 116784
rect 20292 116750 20326 116784
rect 20360 116750 20394 116784
rect 20428 116750 20462 116784
rect 20496 116750 20530 116784
rect 20564 116750 20598 116784
rect 20632 116750 20666 116784
rect 20700 116750 20734 116784
rect 20768 116750 20802 116784
rect 20836 116750 20870 116784
rect 20904 116750 20938 116784
rect 20972 116750 21006 116784
rect 21040 116750 21074 116784
rect 21108 116750 21142 116784
rect 21176 116750 21210 116784
rect 21244 116750 21278 116784
rect 21312 116750 21346 116784
rect 21380 116750 21414 116784
rect 21448 116750 21482 116784
rect 21516 116750 21550 116784
rect 21584 116750 21618 116784
rect 21652 116750 21686 116784
rect 21720 116750 21754 116784
rect 21788 116750 21822 116784
rect 21856 116750 21890 116784
rect 21924 116750 21958 116784
rect 21992 116750 22026 116784
rect 22060 116750 22094 116784
rect 22128 116750 22162 116784
rect 22196 116750 22230 116784
rect 22264 116750 22298 116784
rect 22332 116750 22366 116784
rect 22400 116750 22434 116784
rect 22468 116750 22502 116784
rect 22536 116750 22570 116784
rect 22604 116750 22638 116784
rect 22672 116750 22706 116784
rect 22740 116750 22774 116784
rect 22808 116750 22842 116784
rect 22876 116750 22910 116784
rect 22944 116750 22978 116784
rect 23012 116750 23046 116784
rect 23080 116750 23114 116784
rect 23148 116750 23182 116784
rect 23216 116750 23250 116784
rect 23284 116750 23318 116784
rect 23352 116750 23386 116784
rect 23420 116750 23454 116784
rect 23488 116750 23522 116784
rect 23556 116750 23590 116784
rect 23624 116750 23658 116784
rect 23692 116750 23726 116784
rect 23760 116750 23794 116784
rect 23828 116750 23862 116784
rect 23896 116750 23930 116784
rect 23964 116750 23998 116784
rect 24032 116750 24066 116784
rect 24100 116750 24134 116784
rect 24168 116750 24202 116784
rect 24236 116750 24270 116784
rect 24304 116750 24338 116784
rect 24372 116750 24406 116784
rect 24440 116750 24474 116784
rect 24508 116750 24542 116784
rect 24576 116750 24610 116784
rect 24644 116750 24678 116784
rect 24712 116750 24746 116784
rect 24780 116750 24814 116784
rect 24848 116750 24882 116784
rect 24916 116750 24950 116784
rect 24984 116750 25018 116784
rect 25052 116750 25086 116784
rect 25120 116750 25154 116784
rect 25188 116750 25222 116784
rect 25256 116750 25290 116784
rect 25324 116750 25358 116784
rect 25392 116750 25426 116784
rect 25460 116750 25494 116784
rect 25528 116750 25562 116784
rect 25596 116750 25630 116784
rect 25664 116750 25698 116784
rect 25732 116750 25766 116784
rect 25800 116750 25834 116784
rect 25868 116750 25902 116784
rect 25936 116750 25970 116784
rect 26004 116750 26038 116784
rect 26072 116750 26106 116784
rect 26140 116750 26174 116784
rect 26208 116750 26242 116784
rect 26276 116750 26310 116784
rect 26344 116750 26378 116784
rect 26412 116750 26446 116784
rect 26480 116750 26514 116784
rect 26548 116750 26582 116784
rect 26616 116750 26650 116784
rect 26684 116750 26718 116784
rect 26752 116750 26786 116784
rect 26820 116750 26854 116784
rect 26888 116750 26922 116784
rect 26956 116750 26990 116784
rect 27024 116750 27058 116784
rect 27092 116750 27126 116784
rect 27160 116750 27194 116784
rect 27228 116750 27262 116784
rect 27296 116750 27330 116784
rect 27364 116750 27398 116784
rect 27432 116750 27466 116784
rect 27500 116750 27534 116784
rect 27568 116750 27602 116784
rect 27636 116750 27670 116784
rect 27704 116750 27738 116784
rect 27772 116750 27806 116784
rect 27840 116750 27874 116784
rect 27908 116750 27942 116784
rect 27976 116750 28010 116784
rect 28044 116750 28078 116784
rect 28112 116750 28146 116784
rect 28180 116750 28214 116784
rect 28248 116750 28282 116784
rect 28316 116750 28350 116784
rect 28384 116750 28418 116784
rect 28452 116750 28486 116784
rect 28520 116750 28554 116784
rect 28588 116750 28622 116784
rect 28656 116750 28690 116784
rect 28724 116750 28758 116784
rect 28792 116750 28826 116784
rect 28860 116750 28894 116784
rect 28928 116750 28962 116784
rect 28996 116750 29030 116784
rect 29064 116750 29098 116784
rect 29132 116750 29166 116784
rect 29200 116750 29234 116784
rect 29268 116750 29302 116784
rect 29336 116750 29370 116784
rect 29404 116750 29438 116784
rect 29472 116750 29506 116784
rect 29540 116750 29574 116784
rect 29608 116750 29642 116784
rect 29676 116750 29710 116784
rect 29744 116750 29778 116784
rect 29812 116750 29846 116784
rect 29880 116750 29914 116784
rect 29948 116750 29982 116784
rect 30016 116750 30050 116784
rect 30084 116750 30118 116784
rect 30152 116750 30186 116784
rect 30220 116750 30254 116784
rect 30288 116750 30322 116784
rect 30356 116750 30390 116784
rect 30424 116750 30458 116784
rect 30492 116750 30526 116784
rect 30560 116750 30594 116784
rect 30628 116750 30662 116784
rect 30696 116750 30730 116784
rect 30764 116750 30798 116784
rect 30832 116750 30866 116784
rect 30900 116750 30934 116784
rect 30968 116750 31002 116784
rect 31036 116750 31070 116784
rect 31104 116750 31138 116784
rect 31172 116750 31206 116784
rect 31240 116750 31274 116784
rect 31308 116750 31342 116784
rect 31376 116750 31410 116784
rect 31444 116750 31478 116784
rect 31512 116750 31546 116784
rect 31580 116750 31614 116784
rect 31648 116750 31682 116784
rect 31716 116750 31750 116784
rect 31784 116750 31818 116784
rect 31852 116750 31886 116784
rect 31920 116750 31954 116784
rect 31988 116750 32022 116784
rect 32056 116750 32090 116784
rect 32124 116750 32158 116784
rect 32192 116750 32226 116784
rect 32260 116750 32294 116784
rect 32328 116750 32362 116784
rect 32396 116750 32430 116784
rect 32464 116750 32498 116784
rect 32532 116750 32566 116784
rect 32600 116750 32634 116784
rect 32668 116750 32702 116784
rect 32736 116750 32770 116784
rect 32804 116750 32838 116784
rect 32872 116750 32906 116784
rect 32940 116750 32974 116784
rect 33008 116750 33042 116784
rect 33076 116750 33110 116784
rect 33144 116750 33178 116784
rect 33212 116750 33246 116784
rect 33280 116750 33314 116784
rect 33348 116750 33382 116784
rect 33416 116750 33450 116784
rect 33484 116750 33518 116784
rect 33552 116750 33586 116784
rect 33620 116750 33654 116784
rect 33688 116750 33722 116784
rect 33756 116750 33790 116784
rect 33824 116750 33858 116784
rect 33892 116750 33926 116784
rect 33960 116750 33994 116784
rect 34028 116750 34062 116784
rect 34096 116750 34130 116784
rect 34164 116750 34198 116784
rect 34232 116750 34266 116784
rect 34300 116750 34334 116784
rect 34368 116750 34402 116784
rect 34436 116750 34470 116784
rect 34504 116750 34538 116784
rect 34572 116750 34606 116784
rect 34640 116750 34674 116784
rect 34708 116750 34742 116784
rect 34776 116750 34810 116784
rect 34844 116750 34878 116784
rect 34912 116750 34946 116784
rect 34980 116750 35014 116784
rect 35048 116750 35082 116784
rect 35116 116750 35150 116784
rect 35184 116750 35218 116784
rect 35252 116750 35286 116784
rect 35320 116750 35354 116784
rect 35388 116750 35422 116784
rect 35456 116750 35490 116784
rect 35524 116750 35558 116784
rect 35592 116750 35626 116784
rect 35660 116750 35694 116784
rect 35728 116750 35762 116784
rect 35796 116750 35830 116784
rect 35864 116750 35898 116784
rect 35932 116750 35966 116784
rect 36000 116750 36034 116784
rect 36068 116750 36102 116784
rect 36136 116750 36170 116784
rect 36204 116750 36238 116784
rect 36272 116750 36306 116784
rect 36340 116750 36374 116784
rect 36408 116750 36442 116784
rect 36476 116750 36510 116784
rect 36544 116750 36578 116784
rect 36612 116750 36646 116784
rect 36680 116750 36714 116784
rect 36748 116750 36782 116784
rect 36816 116750 36850 116784
rect 36884 116750 36918 116784
rect 36952 116750 36986 116784
rect 37020 116750 37054 116784
rect 37088 116750 37122 116784
rect 37156 116750 37190 116784
rect 37224 116750 37258 116784
rect 37292 116750 37326 116784
rect 37360 116750 37394 116784
rect 37428 116750 37462 116784
rect 37496 116750 37530 116784
rect 37564 116750 37598 116784
rect 37632 116750 37666 116784
rect 37700 116750 37734 116784
rect 37768 116750 37802 116784
rect 37836 116750 37870 116784
rect 37904 116750 37938 116784
rect 37972 116750 38006 116784
rect 38040 116750 38074 116784
rect 38108 116750 38142 116784
rect 38176 116750 38210 116784
rect 38244 116750 38278 116784
rect 38312 116750 38346 116784
rect 38380 116750 38414 116784
rect 38448 116750 38482 116784
rect 38516 116750 38550 116784
rect 38584 116750 38618 116784
rect 38652 116750 38686 116784
rect 38720 116750 38754 116784
rect 38788 116750 38822 116784
rect 38856 116750 38890 116784
rect 38924 116750 38958 116784
rect 38992 116750 39026 116784
rect 39060 116750 39094 116784
rect 39128 116750 39162 116784
rect 39196 116750 39230 116784
rect 39264 116750 39298 116784
rect 39332 116750 39366 116784
rect 39400 116750 39434 116784
rect 39468 116750 39502 116784
rect 39536 116750 39570 116784
rect 39604 116750 39638 116784
rect 39672 116750 39706 116784
rect 39740 116750 39774 116784
rect 39808 116750 39842 116784
rect 39876 116750 39910 116784
rect 39944 116750 39978 116784
rect 40012 116750 40046 116784
rect 40080 116750 40114 116784
rect 40148 116750 40182 116784
rect 40216 116750 40250 116784
rect 40284 116750 40318 116784
rect 40352 116750 40386 116784
rect 40420 116750 40454 116784
rect 40488 116750 40522 116784
rect 40556 116750 40590 116784
rect 40624 116750 40658 116784
rect 40692 116750 40726 116784
rect 40760 116750 40794 116784
rect 40828 116750 40862 116784
rect 40896 116750 40930 116784
rect 40964 116750 40998 116784
rect 41032 116750 41066 116784
rect 41100 116750 41134 116784
rect 41168 116750 41202 116784
rect 41236 116750 41270 116784
rect 41304 116750 41338 116784
rect 41372 116750 41406 116784
rect 41440 116750 41474 116784
rect 41508 116750 41542 116784
rect 41576 116750 41610 116784
rect 41644 116750 41678 116784
rect 41712 116750 41746 116784
rect 41780 116750 41814 116784
rect 41848 116750 41882 116784
rect 41916 116750 41950 116784
rect 41984 116750 42018 116784
rect 42052 116750 42086 116784
rect 42120 116750 42154 116784
rect 42188 116750 42222 116784
rect 42256 116750 42290 116784
rect 42324 116750 42358 116784
rect 42392 116750 42426 116784
rect 42460 116750 42494 116784
rect 42528 116750 42562 116784
rect 42596 116750 42630 116784
rect 42664 116750 42698 116784
rect 42732 116750 42766 116784
rect 42800 116750 42834 116784
rect 42868 116750 42902 116784
rect 42936 116750 42970 116784
rect 43004 116750 43038 116784
rect 43072 116750 43106 116784
rect 43140 116750 43174 116784
rect 43208 116750 43242 116784
rect 43276 116750 43310 116784
rect 43344 116750 43378 116784
rect 43412 116750 43446 116784
rect 43480 116750 43514 116784
rect 43548 116750 43582 116784
rect 43616 116750 43650 116784
rect 43684 116750 43718 116784
rect 43752 116750 43786 116784
rect 43820 116750 43854 116784
rect 43888 116750 43922 116784
rect 43956 116750 43990 116784
rect 44024 116750 44058 116784
rect 44092 116750 44126 116784
rect 44160 116750 44194 116784
rect 44228 116750 44262 116784
rect 44296 116750 44330 116784
rect 44364 116750 44398 116784
rect 44432 116750 44466 116784
rect 44500 116750 44534 116784
rect 44568 116750 44602 116784
rect 44636 116750 44670 116784
rect 44704 116750 44738 116784
rect 44772 116750 44806 116784
rect 44840 116750 44874 116784
rect 44908 116750 44942 116784
rect 44976 116750 45010 116784
rect 45044 116750 45078 116784
rect 45112 116750 45146 116784
rect 45180 116750 45214 116784
rect 45248 116750 45282 116784
rect 45316 116750 45350 116784
rect 45384 116750 45418 116784
rect 45452 116750 45486 116784
rect 45520 116750 45554 116784
rect 45588 116750 45622 116784
rect 45656 116750 45690 116784
rect 45724 116750 45758 116784
rect 45792 116750 45826 116784
rect 45860 116750 45894 116784
rect 45928 116750 45962 116784
rect 45996 116750 46030 116784
rect 46064 116750 46098 116784
rect 46132 116750 46166 116784
rect 46200 116750 46234 116784
rect 46268 116750 46302 116784
rect 46336 116750 46370 116784
rect 46404 116750 46438 116784
rect 46472 116750 46506 116784
rect 46540 116750 46574 116784
rect 46608 116750 46642 116784
rect 46676 116750 46710 116784
rect 46744 116750 46778 116784
rect 46812 116750 46846 116784
rect 46880 116750 46914 116784
rect 46948 116750 46982 116784
rect 47016 116750 47050 116784
rect 47084 116750 47118 116784
rect 47152 116750 47230 116784
rect -2396 116697 -2362 116750
rect -2396 116629 -2362 116663
rect -2396 116561 -2362 116595
rect -2396 116493 -2362 116527
rect -2396 116425 -2362 116459
rect -2396 116357 -2362 116391
rect -2396 116289 -2362 116323
rect -2396 116221 -2362 116255
rect -2396 116153 -2362 116187
rect -2396 116085 -2362 116119
rect -2396 116017 -2362 116051
rect -2396 115949 -2362 115983
rect -2396 115881 -2362 115915
rect -2396 115813 -2362 115847
rect -2396 115745 -2362 115779
rect -2396 115677 -2362 115711
rect -2396 115609 -2362 115643
rect -2396 115541 -2362 115575
rect -2396 115473 -2362 115507
rect -2396 115405 -2362 115439
rect -2396 115337 -2362 115371
rect -2396 115269 -2362 115303
rect -2396 115201 -2362 115235
rect -2396 115133 -2362 115167
rect -2396 115065 -2362 115099
rect -2396 114997 -2362 115031
rect -2396 114929 -2362 114963
rect -2396 114861 -2362 114895
rect -2396 114793 -2362 114827
rect -2396 114725 -2362 114759
rect -2396 114657 -2362 114691
rect -2396 114589 -2362 114623
rect -2396 114521 -2362 114555
rect -2396 114453 -2362 114487
rect -2396 114385 -2362 114419
rect -2396 114317 -2362 114351
rect -2396 114249 -2362 114283
rect -2396 114181 -2362 114215
rect -2396 114113 -2362 114147
rect -2396 114045 -2362 114079
rect -2396 113977 -2362 114011
rect -2396 113909 -2362 113943
rect -2396 113841 -2362 113875
rect -2396 113773 -2362 113807
rect -2396 113705 -2362 113739
rect -2396 113637 -2362 113671
rect -2396 113569 -2362 113603
rect -2396 113501 -2362 113535
rect -2396 113433 -2362 113467
rect -2396 113365 -2362 113399
rect -2396 113297 -2362 113331
rect -2396 113229 -2362 113263
rect -2396 113161 -2362 113195
rect -2396 113093 -2362 113127
rect -2396 113025 -2362 113059
rect -2396 112957 -2362 112991
rect -2396 112889 -2362 112923
rect -2396 112821 -2362 112855
rect -2396 112753 -2362 112787
rect -2396 112685 -2362 112719
rect -2396 112617 -2362 112651
rect -2396 112549 -2362 112583
rect -2396 112481 -2362 112515
rect -2396 112413 -2362 112447
rect -2396 112345 -2362 112379
rect -2396 112277 -2362 112311
rect -2396 112209 -2362 112243
rect -2396 112141 -2362 112175
rect -2396 112073 -2362 112107
rect -2396 112005 -2362 112039
rect -2396 111937 -2362 111971
rect -2396 111869 -2362 111903
rect -2396 111801 -2362 111835
rect -2396 111733 -2362 111767
rect -2396 111665 -2362 111699
rect -2396 111597 -2362 111631
rect -2396 111529 -2362 111563
rect -2396 111461 -2362 111495
rect -2396 111393 -2362 111427
rect -2396 111325 -2362 111359
rect -2396 111257 -2362 111291
rect -2396 111189 -2362 111223
rect -2396 111121 -2362 111155
rect -2396 111053 -2362 111087
rect -2396 110985 -2362 111019
rect -2396 110917 -2362 110951
rect -2396 110849 -2362 110883
rect -2396 110781 -2362 110815
rect -2396 110713 -2362 110747
rect -2396 110645 -2362 110679
rect -2396 110577 -2362 110611
rect -2396 110509 -2362 110543
rect -2396 110441 -2362 110475
rect -2396 110373 -2362 110407
rect -2396 110305 -2362 110339
rect -2396 110237 -2362 110271
rect -2396 110169 -2362 110203
rect -2396 110101 -2362 110135
rect -2396 110033 -2362 110067
rect -2396 109965 -2362 109999
rect -2396 109897 -2362 109931
rect -2396 109829 -2362 109863
rect -2396 109761 -2362 109795
rect -2396 109693 -2362 109727
rect -2396 109625 -2362 109659
rect -2396 109557 -2362 109591
rect -2396 109489 -2362 109523
rect -2396 109421 -2362 109455
rect -2396 109353 -2362 109387
rect -2396 109285 -2362 109319
rect -2396 109217 -2362 109251
rect -2396 109149 -2362 109183
rect -2396 109081 -2362 109115
rect -2396 109013 -2362 109047
rect -2396 108945 -2362 108979
rect -2396 108877 -2362 108911
rect -2396 108809 -2362 108843
rect -2396 108741 -2362 108775
rect -2396 108673 -2362 108707
rect -2396 108605 -2362 108639
rect -2396 108537 -2362 108571
rect -2396 108469 -2362 108503
rect -2396 108401 -2362 108435
rect -2396 108333 -2362 108367
rect -2396 108265 -2362 108299
rect -2396 108197 -2362 108231
rect -2396 108129 -2362 108163
rect -2396 108061 -2362 108095
rect -2396 107993 -2362 108027
rect -2396 107925 -2362 107959
rect -2396 107857 -2362 107891
rect -2396 107789 -2362 107823
rect -2396 107721 -2362 107755
rect -2396 107653 -2362 107687
rect -2396 107585 -2362 107619
rect -2396 107517 -2362 107551
rect -2396 107449 -2362 107483
rect -2396 107381 -2362 107415
rect -2396 107313 -2362 107347
rect -2396 107245 -2362 107279
rect -2396 107177 -2362 107211
rect -2396 107109 -2362 107143
rect -2396 107041 -2362 107075
rect -2396 106973 -2362 107007
rect -2396 106905 -2362 106939
rect -2396 106837 -2362 106871
rect -2396 106769 -2362 106803
rect -2396 106701 -2362 106735
rect -2396 106633 -2362 106667
rect -2396 106565 -2362 106599
rect -2396 106497 -2362 106531
rect -2396 106429 -2362 106463
rect -2396 106361 -2362 106395
rect -2396 106293 -2362 106327
rect -2396 106225 -2362 106259
rect -2396 106157 -2362 106191
rect -2396 106089 -2362 106123
rect -2396 106021 -2362 106055
rect -2396 105953 -2362 105987
rect -2396 105885 -2362 105919
rect -2396 105817 -2362 105851
rect -2396 105749 -2362 105783
rect -2396 105681 -2362 105715
rect -2396 105613 -2362 105647
rect -2396 105545 -2362 105579
rect -2396 105477 -2362 105511
rect -2396 105409 -2362 105443
rect -2396 105341 -2362 105375
rect -2396 105273 -2362 105307
rect -2396 105205 -2362 105239
rect -2396 105137 -2362 105171
rect -2396 105069 -2362 105103
rect -2396 105001 -2362 105035
rect -2396 104933 -2362 104967
rect -2396 104865 -2362 104899
rect -2396 104797 -2362 104831
rect -2396 104729 -2362 104763
rect -2396 104661 -2362 104695
rect -2396 104593 -2362 104627
rect -2396 104525 -2362 104559
rect -2396 104457 -2362 104491
rect -2396 104389 -2362 104423
rect -2396 104321 -2362 104355
rect -2396 104253 -2362 104287
rect -2396 104185 -2362 104219
rect -2396 104117 -2362 104151
rect -2396 104049 -2362 104083
rect -2396 103981 -2362 104015
rect -2396 103913 -2362 103947
rect -2396 103845 -2362 103879
rect -2396 103777 -2362 103811
rect -2396 103709 -2362 103743
rect -2396 103641 -2362 103675
rect -2396 103573 -2362 103607
rect -2396 103505 -2362 103539
rect -2396 103437 -2362 103471
rect -2396 103369 -2362 103403
rect -2396 103301 -2362 103335
rect -2396 103233 -2362 103267
rect -2396 103165 -2362 103199
rect -2396 103097 -2362 103131
rect -2396 103029 -2362 103063
rect -2396 102961 -2362 102995
rect -2396 102893 -2362 102927
rect -2396 102825 -2362 102859
rect -2396 102757 -2362 102791
rect -2396 102689 -2362 102723
rect -2396 102621 -2362 102655
rect -2396 102553 -2362 102587
rect -2396 102485 -2362 102519
rect -2396 102417 -2362 102451
rect -2396 102349 -2362 102383
rect -2396 102281 -2362 102315
rect -2396 102213 -2362 102247
rect -2396 102145 -2362 102179
rect -2396 102077 -2362 102111
rect -2396 102009 -2362 102043
rect -2396 101941 -2362 101975
rect -2396 101873 -2362 101907
rect -2396 101805 -2362 101839
rect -2396 101737 -2362 101771
rect -2396 101669 -2362 101703
rect -2396 101601 -2362 101635
rect -2396 101533 -2362 101567
rect -2396 101465 -2362 101499
rect -2396 101397 -2362 101431
rect -2396 101329 -2362 101363
rect -2396 101261 -2362 101295
rect -2396 101193 -2362 101227
rect -2396 101125 -2362 101159
rect -2396 101057 -2362 101091
rect -2396 100989 -2362 101023
rect -2396 100903 -2362 100955
rect 47196 116697 47230 116750
rect 47196 116629 47230 116663
rect 47196 116561 47230 116595
rect 47196 116493 47230 116527
rect 47196 116425 47230 116459
rect 47196 116357 47230 116391
rect 47196 116289 47230 116323
rect 47196 116221 47230 116255
rect 47196 116153 47230 116187
rect 47196 116085 47230 116119
rect 47196 116017 47230 116051
rect 47196 115949 47230 115983
rect 47196 115881 47230 115915
rect 47196 115813 47230 115847
rect 47196 115745 47230 115779
rect 47196 115677 47230 115711
rect 47196 115609 47230 115643
rect 47196 115541 47230 115575
rect 47196 115473 47230 115507
rect 47196 115405 47230 115439
rect 47196 115337 47230 115371
rect 47196 115269 47230 115303
rect 47196 115201 47230 115235
rect 47196 115133 47230 115167
rect 47196 115065 47230 115099
rect 47196 114997 47230 115031
rect 47196 114929 47230 114963
rect 47196 114861 47230 114895
rect 47196 114793 47230 114827
rect 47196 114725 47230 114759
rect 47196 114657 47230 114691
rect 47196 114589 47230 114623
rect 47196 114521 47230 114555
rect 47196 114453 47230 114487
rect 47196 114385 47230 114419
rect 47196 114317 47230 114351
rect 47196 114249 47230 114283
rect 47196 114181 47230 114215
rect 47196 114113 47230 114147
rect 47196 114045 47230 114079
rect 47196 113977 47230 114011
rect 47196 113909 47230 113943
rect 47196 113841 47230 113875
rect 47196 113773 47230 113807
rect 47196 113705 47230 113739
rect 47196 113637 47230 113671
rect 47196 113569 47230 113603
rect 47196 113501 47230 113535
rect 47196 113433 47230 113467
rect 47196 113365 47230 113399
rect 47196 113297 47230 113331
rect 47196 113229 47230 113263
rect 47196 113161 47230 113195
rect 47196 113093 47230 113127
rect 47196 113025 47230 113059
rect 47196 112957 47230 112991
rect 47196 112889 47230 112923
rect 47196 112821 47230 112855
rect 47196 112753 47230 112787
rect 47196 112685 47230 112719
rect 47196 112617 47230 112651
rect 47196 112549 47230 112583
rect 47196 112481 47230 112515
rect 47196 112413 47230 112447
rect 47196 112345 47230 112379
rect 47196 112277 47230 112311
rect 47196 112209 47230 112243
rect 47196 112141 47230 112175
rect 47196 112073 47230 112107
rect 47196 112005 47230 112039
rect 47196 111937 47230 111971
rect 47196 111869 47230 111903
rect 47196 111801 47230 111835
rect 47196 111733 47230 111767
rect 47196 111665 47230 111699
rect 47196 111597 47230 111631
rect 47196 111529 47230 111563
rect 47196 111461 47230 111495
rect 47196 111393 47230 111427
rect 47196 111325 47230 111359
rect 47196 111257 47230 111291
rect 47196 111189 47230 111223
rect 47196 111121 47230 111155
rect 47196 111053 47230 111087
rect 47196 110985 47230 111019
rect 47196 110917 47230 110951
rect 47196 110849 47230 110883
rect 47196 110781 47230 110815
rect 47196 110713 47230 110747
rect 47196 110645 47230 110679
rect 47196 110577 47230 110611
rect 47196 110509 47230 110543
rect 47196 110441 47230 110475
rect 47196 110373 47230 110407
rect 47196 110305 47230 110339
rect 47196 110237 47230 110271
rect 47196 110169 47230 110203
rect 47196 110101 47230 110135
rect 47196 110033 47230 110067
rect 47196 109965 47230 109999
rect 47196 109897 47230 109931
rect 47196 109829 47230 109863
rect 47196 109761 47230 109795
rect 47196 109693 47230 109727
rect 47196 109625 47230 109659
rect 47196 109557 47230 109591
rect 47196 109489 47230 109523
rect 47196 109421 47230 109455
rect 47196 109353 47230 109387
rect 47196 109285 47230 109319
rect 47196 109217 47230 109251
rect 47196 109149 47230 109183
rect 47196 109081 47230 109115
rect 47196 109013 47230 109047
rect 47196 108945 47230 108979
rect 47196 108877 47230 108911
rect 47196 108809 47230 108843
rect 47196 108741 47230 108775
rect 47196 108673 47230 108707
rect 47196 108605 47230 108639
rect 47196 108537 47230 108571
rect 47196 108469 47230 108503
rect 47196 108401 47230 108435
rect 47196 108333 47230 108367
rect 47196 108265 47230 108299
rect 47196 108197 47230 108231
rect 47196 108129 47230 108163
rect 47196 108061 47230 108095
rect 47196 107993 47230 108027
rect 47196 107925 47230 107959
rect 47196 107857 47230 107891
rect 47196 107789 47230 107823
rect 47196 107721 47230 107755
rect 47196 107653 47230 107687
rect 47196 107585 47230 107619
rect 47196 107517 47230 107551
rect 47196 107449 47230 107483
rect 47196 107381 47230 107415
rect 47196 107313 47230 107347
rect 47196 107245 47230 107279
rect 47196 107177 47230 107211
rect 47196 107109 47230 107143
rect 47196 107041 47230 107075
rect 47196 106973 47230 107007
rect 47196 106905 47230 106939
rect 47196 106837 47230 106871
rect 47196 106769 47230 106803
rect 47196 106701 47230 106735
rect 47196 106633 47230 106667
rect 47196 106565 47230 106599
rect 47196 106497 47230 106531
rect 47196 106429 47230 106463
rect 47196 106361 47230 106395
rect 47196 106293 47230 106327
rect 47196 106225 47230 106259
rect 47196 106157 47230 106191
rect 47196 106089 47230 106123
rect 47196 106021 47230 106055
rect 47196 105953 47230 105987
rect 47196 105885 47230 105919
rect 47196 105817 47230 105851
rect 47196 105749 47230 105783
rect 47196 105681 47230 105715
rect 47196 105613 47230 105647
rect 47196 105545 47230 105579
rect 47196 105477 47230 105511
rect 47196 105409 47230 105443
rect 47196 105341 47230 105375
rect 47196 105273 47230 105307
rect 47196 105205 47230 105239
rect 47196 105137 47230 105171
rect 47196 105069 47230 105103
rect 47196 105001 47230 105035
rect 47196 104933 47230 104967
rect 47196 104865 47230 104899
rect 47196 104797 47230 104831
rect 47196 104729 47230 104763
rect 47196 104661 47230 104695
rect 47196 104593 47230 104627
rect 47196 104525 47230 104559
rect 47196 104457 47230 104491
rect 47196 104389 47230 104423
rect 47196 104321 47230 104355
rect 47196 104253 47230 104287
rect 47196 104185 47230 104219
rect 47196 104117 47230 104151
rect 47196 104049 47230 104083
rect 47196 103981 47230 104015
rect 47196 103913 47230 103947
rect 47196 103845 47230 103879
rect 47196 103777 47230 103811
rect 47196 103709 47230 103743
rect 47196 103641 47230 103675
rect 47196 103573 47230 103607
rect 47196 103505 47230 103539
rect 47196 103437 47230 103471
rect 47196 103369 47230 103403
rect 47196 103301 47230 103335
rect 47196 103233 47230 103267
rect 47196 103165 47230 103199
rect 47196 103097 47230 103131
rect 47196 103029 47230 103063
rect 47196 102961 47230 102995
rect 47196 102893 47230 102927
rect 47196 102825 47230 102859
rect 47196 102757 47230 102791
rect 47196 102689 47230 102723
rect 47196 102621 47230 102655
rect 47196 102553 47230 102587
rect 47196 102485 47230 102519
rect 47196 102417 47230 102451
rect 47196 102349 47230 102383
rect 47196 102281 47230 102315
rect 47196 102213 47230 102247
rect 47196 102145 47230 102179
rect 47196 102077 47230 102111
rect 47196 102009 47230 102043
rect 47196 101941 47230 101975
rect 47196 101873 47230 101907
rect 47196 101805 47230 101839
rect 47196 101737 47230 101771
rect 47196 101669 47230 101703
rect 47196 101601 47230 101635
rect 47196 101533 47230 101567
rect 47196 101465 47230 101499
rect 47196 101397 47230 101431
rect 47196 101329 47230 101363
rect 47196 101261 47230 101295
rect 47196 101193 47230 101227
rect 47196 101125 47230 101159
rect 47196 101057 47230 101091
rect 47196 100989 47230 101023
rect 47196 100903 47230 100955
rect -2396 100869 -2318 100903
rect -2284 100869 -2250 100903
rect -2216 100869 -2182 100903
rect -2148 100869 -2114 100903
rect -2080 100869 -2046 100903
rect -2012 100869 -1978 100903
rect -1944 100869 -1910 100903
rect -1876 100869 -1842 100903
rect -1808 100869 -1774 100903
rect -1740 100869 -1706 100903
rect -1672 100869 -1638 100903
rect -1604 100869 -1570 100903
rect -1536 100869 -1502 100903
rect -1468 100869 -1434 100903
rect -1400 100869 -1366 100903
rect -1332 100869 -1298 100903
rect -1264 100869 -1230 100903
rect -1196 100869 -1162 100903
rect -1128 100869 -1094 100903
rect -1060 100869 -1026 100903
rect -992 100869 -958 100903
rect -924 100869 -890 100903
rect -856 100869 -822 100903
rect -788 100869 -754 100903
rect -720 100869 -686 100903
rect -652 100869 -618 100903
rect -584 100869 -550 100903
rect -516 100869 -482 100903
rect -448 100869 -414 100903
rect -380 100869 -346 100903
rect -312 100869 -278 100903
rect -244 100869 -210 100903
rect -176 100869 -142 100903
rect -108 100869 -74 100903
rect -40 100869 -6 100903
rect 28 100869 62 100903
rect 96 100869 130 100903
rect 164 100869 198 100903
rect 232 100869 266 100903
rect 300 100869 334 100903
rect 368 100869 402 100903
rect 436 100869 470 100903
rect 504 100869 538 100903
rect 572 100869 606 100903
rect 640 100869 674 100903
rect 708 100869 742 100903
rect 776 100869 810 100903
rect 844 100869 878 100903
rect 912 100869 946 100903
rect 980 100869 1014 100903
rect 1048 100869 1082 100903
rect 1116 100869 1150 100903
rect 1184 100869 1218 100903
rect 1252 100869 1286 100903
rect 1320 100869 1354 100903
rect 1388 100869 1422 100903
rect 1456 100869 1490 100903
rect 1524 100869 1558 100903
rect 1592 100869 1626 100903
rect 1660 100869 1694 100903
rect 1728 100869 1762 100903
rect 1796 100869 1830 100903
rect 1864 100869 1898 100903
rect 1932 100869 1966 100903
rect 2000 100869 2034 100903
rect 2068 100869 2102 100903
rect 2136 100869 2170 100903
rect 2204 100869 2238 100903
rect 2272 100869 2306 100903
rect 2340 100869 2374 100903
rect 2408 100869 2442 100903
rect 2476 100869 2510 100903
rect 2544 100869 2578 100903
rect 2612 100869 2646 100903
rect 2680 100869 2714 100903
rect 2748 100869 2782 100903
rect 2816 100869 2850 100903
rect 2884 100869 2918 100903
rect 2952 100869 2986 100903
rect 3020 100869 3054 100903
rect 3088 100869 3122 100903
rect 3156 100869 3190 100903
rect 3224 100869 3258 100903
rect 3292 100869 3326 100903
rect 3360 100869 3394 100903
rect 3428 100869 3462 100903
rect 3496 100869 3530 100903
rect 3564 100869 3598 100903
rect 3632 100869 3666 100903
rect 3700 100869 3734 100903
rect 3768 100869 3802 100903
rect 3836 100869 3870 100903
rect 3904 100869 3938 100903
rect 3972 100869 4006 100903
rect 4040 100869 4074 100903
rect 4108 100869 4142 100903
rect 4176 100869 4210 100903
rect 4244 100869 4278 100903
rect 4312 100869 4346 100903
rect 4380 100869 4414 100903
rect 4448 100869 4482 100903
rect 4516 100869 4550 100903
rect 4584 100869 4618 100903
rect 4652 100869 4686 100903
rect 4720 100869 4754 100903
rect 4788 100869 4822 100903
rect 4856 100869 4890 100903
rect 4924 100869 4958 100903
rect 4992 100869 5026 100903
rect 5060 100869 5094 100903
rect 5128 100869 5162 100903
rect 5196 100869 5230 100903
rect 5264 100869 5298 100903
rect 5332 100869 5366 100903
rect 5400 100869 5434 100903
rect 5468 100869 5502 100903
rect 5536 100869 5570 100903
rect 5604 100869 5638 100903
rect 5672 100869 5706 100903
rect 5740 100869 5774 100903
rect 5808 100869 5842 100903
rect 5876 100869 5910 100903
rect 5944 100869 5978 100903
rect 6012 100869 6046 100903
rect 6080 100869 6114 100903
rect 6148 100869 6182 100903
rect 6216 100869 6250 100903
rect 6284 100869 6318 100903
rect 6352 100869 6386 100903
rect 6420 100869 6454 100903
rect 6488 100869 6522 100903
rect 6556 100869 6590 100903
rect 6624 100869 6658 100903
rect 6692 100869 6726 100903
rect 6760 100869 6794 100903
rect 6828 100869 6862 100903
rect 6896 100869 6930 100903
rect 6964 100869 6998 100903
rect 7032 100869 7066 100903
rect 7100 100869 7134 100903
rect 7168 100869 7202 100903
rect 7236 100869 7270 100903
rect 7304 100869 7338 100903
rect 7372 100869 7406 100903
rect 7440 100869 7474 100903
rect 7508 100869 7542 100903
rect 7576 100869 7610 100903
rect 7644 100869 7678 100903
rect 7712 100869 7746 100903
rect 7780 100869 7814 100903
rect 7848 100869 7882 100903
rect 7916 100869 7950 100903
rect 7984 100869 8018 100903
rect 8052 100869 8086 100903
rect 8120 100869 8154 100903
rect 8188 100869 8222 100903
rect 8256 100869 8290 100903
rect 8324 100869 8358 100903
rect 8392 100869 8426 100903
rect 8460 100869 8494 100903
rect 8528 100869 8562 100903
rect 8596 100869 8630 100903
rect 8664 100869 8698 100903
rect 8732 100869 8766 100903
rect 8800 100869 8834 100903
rect 8868 100869 8902 100903
rect 8936 100869 8970 100903
rect 9004 100869 9038 100903
rect 9072 100869 9106 100903
rect 9140 100869 9174 100903
rect 9208 100869 9242 100903
rect 9276 100869 9310 100903
rect 9344 100869 9378 100903
rect 9412 100869 9446 100903
rect 9480 100869 9514 100903
rect 9548 100869 9582 100903
rect 9616 100869 9650 100903
rect 9684 100869 9718 100903
rect 9752 100869 9786 100903
rect 9820 100869 9854 100903
rect 9888 100869 9922 100903
rect 9956 100869 9990 100903
rect 10024 100869 10058 100903
rect 10092 100869 10126 100903
rect 10160 100869 10194 100903
rect 10228 100869 10262 100903
rect 10296 100869 10330 100903
rect 10364 100869 10398 100903
rect 10432 100869 10466 100903
rect 10500 100869 10534 100903
rect 10568 100869 10602 100903
rect 10636 100869 10670 100903
rect 10704 100869 10738 100903
rect 10772 100869 10806 100903
rect 10840 100869 10874 100903
rect 10908 100869 10942 100903
rect 10976 100869 11010 100903
rect 11044 100869 11078 100903
rect 11112 100869 11146 100903
rect 11180 100869 11214 100903
rect 11248 100869 11282 100903
rect 11316 100869 11350 100903
rect 11384 100869 11418 100903
rect 11452 100869 11486 100903
rect 11520 100869 11554 100903
rect 11588 100869 11622 100903
rect 11656 100869 11690 100903
rect 11724 100869 11758 100903
rect 11792 100869 11826 100903
rect 11860 100869 11894 100903
rect 11928 100869 11962 100903
rect 11996 100869 12030 100903
rect 12064 100869 12098 100903
rect 12132 100869 12166 100903
rect 12200 100869 12234 100903
rect 12268 100869 12302 100903
rect 12336 100869 12370 100903
rect 12404 100869 12438 100903
rect 12472 100869 12506 100903
rect 12540 100869 12574 100903
rect 12608 100869 12642 100903
rect 12676 100869 12710 100903
rect 12744 100869 12778 100903
rect 12812 100869 12846 100903
rect 12880 100869 12914 100903
rect 12948 100869 12982 100903
rect 13016 100869 13050 100903
rect 13084 100869 13118 100903
rect 13152 100869 13186 100903
rect 13220 100869 13254 100903
rect 13288 100869 13322 100903
rect 13356 100869 13390 100903
rect 13424 100869 13458 100903
rect 13492 100869 13526 100903
rect 13560 100869 13594 100903
rect 13628 100869 13662 100903
rect 13696 100869 13730 100903
rect 13764 100869 13798 100903
rect 13832 100869 13866 100903
rect 13900 100869 13934 100903
rect 13968 100869 14002 100903
rect 14036 100869 14070 100903
rect 14104 100869 14138 100903
rect 14172 100869 14206 100903
rect 14240 100869 14274 100903
rect 14308 100869 14342 100903
rect 14376 100869 14410 100903
rect 14444 100869 14478 100903
rect 14512 100869 14546 100903
rect 14580 100869 14614 100903
rect 14648 100869 14682 100903
rect 14716 100869 14750 100903
rect 14784 100869 14818 100903
rect 14852 100869 14886 100903
rect 14920 100869 14954 100903
rect 14988 100869 15022 100903
rect 15056 100869 15090 100903
rect 15124 100869 15158 100903
rect 15192 100869 15226 100903
rect 15260 100869 15294 100903
rect 15328 100869 15362 100903
rect 15396 100869 15430 100903
rect 15464 100869 15498 100903
rect 15532 100869 15566 100903
rect 15600 100869 15634 100903
rect 15668 100869 15702 100903
rect 15736 100869 15770 100903
rect 15804 100869 15838 100903
rect 15872 100869 15906 100903
rect 15940 100869 15974 100903
rect 16008 100869 16042 100903
rect 16076 100869 16110 100903
rect 16144 100869 16178 100903
rect 16212 100869 16246 100903
rect 16280 100869 16314 100903
rect 16348 100869 16382 100903
rect 16416 100869 16450 100903
rect 16484 100869 16518 100903
rect 16552 100869 16586 100903
rect 16620 100869 16654 100903
rect 16688 100869 16722 100903
rect 16756 100869 16790 100903
rect 16824 100869 16858 100903
rect 16892 100869 16926 100903
rect 16960 100869 16994 100903
rect 17028 100869 17062 100903
rect 17096 100869 17130 100903
rect 17164 100869 17198 100903
rect 17232 100869 17266 100903
rect 17300 100869 17334 100903
rect 17368 100869 17402 100903
rect 17436 100869 17470 100903
rect 17504 100869 17538 100903
rect 17572 100869 17606 100903
rect 17640 100869 17674 100903
rect 17708 100869 17742 100903
rect 17776 100869 17810 100903
rect 17844 100869 17878 100903
rect 17912 100869 17946 100903
rect 17980 100869 18014 100903
rect 18048 100869 18082 100903
rect 18116 100869 18150 100903
rect 18184 100869 18218 100903
rect 18252 100869 18286 100903
rect 18320 100869 18354 100903
rect 18388 100869 18422 100903
rect 18456 100869 18490 100903
rect 18524 100869 18558 100903
rect 18592 100869 18626 100903
rect 18660 100869 18694 100903
rect 18728 100869 18762 100903
rect 18796 100869 18830 100903
rect 18864 100869 18898 100903
rect 18932 100869 18966 100903
rect 19000 100869 19034 100903
rect 19068 100869 19102 100903
rect 19136 100869 19170 100903
rect 19204 100869 19238 100903
rect 19272 100869 19306 100903
rect 19340 100869 19374 100903
rect 19408 100869 19442 100903
rect 19476 100869 19510 100903
rect 19544 100869 19578 100903
rect 19612 100869 19646 100903
rect 19680 100869 19714 100903
rect 19748 100869 19782 100903
rect 19816 100869 19850 100903
rect 19884 100869 19918 100903
rect 19952 100869 19986 100903
rect 20020 100869 20054 100903
rect 20088 100869 20122 100903
rect 20156 100869 20190 100903
rect 20224 100869 20258 100903
rect 20292 100869 20326 100903
rect 20360 100869 20394 100903
rect 20428 100869 20462 100903
rect 20496 100869 20530 100903
rect 20564 100869 20598 100903
rect 20632 100869 20666 100903
rect 20700 100869 20734 100903
rect 20768 100869 20802 100903
rect 20836 100869 20870 100903
rect 20904 100869 20938 100903
rect 20972 100869 21006 100903
rect 21040 100869 21074 100903
rect 21108 100869 21142 100903
rect 21176 100869 21210 100903
rect 21244 100869 21278 100903
rect 21312 100869 21346 100903
rect 21380 100869 21414 100903
rect 21448 100869 21482 100903
rect 21516 100869 21550 100903
rect 21584 100869 21618 100903
rect 21652 100869 21686 100903
rect 21720 100869 21754 100903
rect 21788 100869 21822 100903
rect 21856 100869 21890 100903
rect 21924 100869 21958 100903
rect 21992 100869 22026 100903
rect 22060 100869 22094 100903
rect 22128 100869 22162 100903
rect 22196 100869 22230 100903
rect 22264 100869 22298 100903
rect 22332 100869 22366 100903
rect 22400 100869 22434 100903
rect 22468 100869 22502 100903
rect 22536 100869 22570 100903
rect 22604 100869 22638 100903
rect 22672 100869 22706 100903
rect 22740 100869 22774 100903
rect 22808 100869 22842 100903
rect 22876 100869 22910 100903
rect 22944 100869 22978 100903
rect 23012 100869 23046 100903
rect 23080 100869 23114 100903
rect 23148 100869 23182 100903
rect 23216 100869 23250 100903
rect 23284 100869 23318 100903
rect 23352 100869 23386 100903
rect 23420 100869 23454 100903
rect 23488 100869 23522 100903
rect 23556 100869 23590 100903
rect 23624 100869 23658 100903
rect 23692 100869 23726 100903
rect 23760 100869 23794 100903
rect 23828 100869 23862 100903
rect 23896 100869 23930 100903
rect 23964 100869 23998 100903
rect 24032 100869 24066 100903
rect 24100 100869 24134 100903
rect 24168 100869 24202 100903
rect 24236 100869 24270 100903
rect 24304 100869 24338 100903
rect 24372 100869 24406 100903
rect 24440 100869 24474 100903
rect 24508 100869 24542 100903
rect 24576 100869 24610 100903
rect 24644 100869 24678 100903
rect 24712 100869 24746 100903
rect 24780 100869 24814 100903
rect 24848 100869 24882 100903
rect 24916 100869 24950 100903
rect 24984 100869 25018 100903
rect 25052 100869 25086 100903
rect 25120 100869 25154 100903
rect 25188 100869 25222 100903
rect 25256 100869 25290 100903
rect 25324 100869 25358 100903
rect 25392 100869 25426 100903
rect 25460 100869 25494 100903
rect 25528 100869 25562 100903
rect 25596 100869 25630 100903
rect 25664 100869 25698 100903
rect 25732 100869 25766 100903
rect 25800 100869 25834 100903
rect 25868 100869 25902 100903
rect 25936 100869 25970 100903
rect 26004 100869 26038 100903
rect 26072 100869 26106 100903
rect 26140 100869 26174 100903
rect 26208 100869 26242 100903
rect 26276 100869 26310 100903
rect 26344 100869 26378 100903
rect 26412 100869 26446 100903
rect 26480 100869 26514 100903
rect 26548 100869 26582 100903
rect 26616 100869 26650 100903
rect 26684 100869 26718 100903
rect 26752 100869 26786 100903
rect 26820 100869 26854 100903
rect 26888 100869 26922 100903
rect 26956 100869 26990 100903
rect 27024 100869 27058 100903
rect 27092 100869 27126 100903
rect 27160 100869 27194 100903
rect 27228 100869 27262 100903
rect 27296 100869 27330 100903
rect 27364 100869 27398 100903
rect 27432 100869 27466 100903
rect 27500 100869 27534 100903
rect 27568 100869 27602 100903
rect 27636 100869 27670 100903
rect 27704 100869 27738 100903
rect 27772 100869 27806 100903
rect 27840 100869 27874 100903
rect 27908 100869 27942 100903
rect 27976 100869 28010 100903
rect 28044 100869 28078 100903
rect 28112 100869 28146 100903
rect 28180 100869 28214 100903
rect 28248 100869 28282 100903
rect 28316 100869 28350 100903
rect 28384 100869 28418 100903
rect 28452 100869 28486 100903
rect 28520 100869 28554 100903
rect 28588 100869 28622 100903
rect 28656 100869 28690 100903
rect 28724 100869 28758 100903
rect 28792 100869 28826 100903
rect 28860 100869 28894 100903
rect 28928 100869 28962 100903
rect 28996 100869 29030 100903
rect 29064 100869 29098 100903
rect 29132 100869 29166 100903
rect 29200 100869 29234 100903
rect 29268 100869 29302 100903
rect 29336 100869 29370 100903
rect 29404 100869 29438 100903
rect 29472 100869 29506 100903
rect 29540 100869 29574 100903
rect 29608 100869 29642 100903
rect 29676 100869 29710 100903
rect 29744 100869 29778 100903
rect 29812 100869 29846 100903
rect 29880 100869 29914 100903
rect 29948 100869 29982 100903
rect 30016 100869 30050 100903
rect 30084 100869 30118 100903
rect 30152 100869 30186 100903
rect 30220 100869 30254 100903
rect 30288 100869 30322 100903
rect 30356 100869 30390 100903
rect 30424 100869 30458 100903
rect 30492 100869 30526 100903
rect 30560 100869 30594 100903
rect 30628 100869 30662 100903
rect 30696 100869 30730 100903
rect 30764 100869 30798 100903
rect 30832 100869 30866 100903
rect 30900 100869 30934 100903
rect 30968 100869 31002 100903
rect 31036 100869 31070 100903
rect 31104 100869 31138 100903
rect 31172 100869 31206 100903
rect 31240 100869 31274 100903
rect 31308 100869 31342 100903
rect 31376 100869 31410 100903
rect 31444 100869 31478 100903
rect 31512 100869 31546 100903
rect 31580 100869 31614 100903
rect 31648 100869 31682 100903
rect 31716 100869 31750 100903
rect 31784 100869 31818 100903
rect 31852 100869 31886 100903
rect 31920 100869 31954 100903
rect 31988 100869 32022 100903
rect 32056 100869 32090 100903
rect 32124 100869 32158 100903
rect 32192 100869 32226 100903
rect 32260 100869 32294 100903
rect 32328 100869 32362 100903
rect 32396 100869 32430 100903
rect 32464 100869 32498 100903
rect 32532 100869 32566 100903
rect 32600 100869 32634 100903
rect 32668 100869 32702 100903
rect 32736 100869 32770 100903
rect 32804 100869 32838 100903
rect 32872 100869 32906 100903
rect 32940 100869 32974 100903
rect 33008 100869 33042 100903
rect 33076 100869 33110 100903
rect 33144 100869 33178 100903
rect 33212 100869 33246 100903
rect 33280 100869 33314 100903
rect 33348 100869 33382 100903
rect 33416 100869 33450 100903
rect 33484 100869 33518 100903
rect 33552 100869 33586 100903
rect 33620 100869 33654 100903
rect 33688 100869 33722 100903
rect 33756 100869 33790 100903
rect 33824 100869 33858 100903
rect 33892 100869 33926 100903
rect 33960 100869 33994 100903
rect 34028 100869 34062 100903
rect 34096 100869 34130 100903
rect 34164 100869 34198 100903
rect 34232 100869 34266 100903
rect 34300 100869 34334 100903
rect 34368 100869 34402 100903
rect 34436 100869 34470 100903
rect 34504 100869 34538 100903
rect 34572 100869 34606 100903
rect 34640 100869 34674 100903
rect 34708 100869 34742 100903
rect 34776 100869 34810 100903
rect 34844 100869 34878 100903
rect 34912 100869 34946 100903
rect 34980 100869 35014 100903
rect 35048 100869 35082 100903
rect 35116 100869 35150 100903
rect 35184 100869 35218 100903
rect 35252 100869 35286 100903
rect 35320 100869 35354 100903
rect 35388 100869 35422 100903
rect 35456 100869 35490 100903
rect 35524 100869 35558 100903
rect 35592 100869 35626 100903
rect 35660 100869 35694 100903
rect 35728 100869 35762 100903
rect 35796 100869 35830 100903
rect 35864 100869 35898 100903
rect 35932 100869 35966 100903
rect 36000 100869 36034 100903
rect 36068 100869 36102 100903
rect 36136 100869 36170 100903
rect 36204 100869 36238 100903
rect 36272 100869 36306 100903
rect 36340 100869 36374 100903
rect 36408 100869 36442 100903
rect 36476 100869 36510 100903
rect 36544 100869 36578 100903
rect 36612 100869 36646 100903
rect 36680 100869 36714 100903
rect 36748 100869 36782 100903
rect 36816 100869 36850 100903
rect 36884 100869 36918 100903
rect 36952 100869 36986 100903
rect 37020 100869 37054 100903
rect 37088 100869 37122 100903
rect 37156 100869 37190 100903
rect 37224 100869 37258 100903
rect 37292 100869 37326 100903
rect 37360 100869 37394 100903
rect 37428 100869 37462 100903
rect 37496 100869 37530 100903
rect 37564 100869 37598 100903
rect 37632 100869 37666 100903
rect 37700 100869 37734 100903
rect 37768 100869 37802 100903
rect 37836 100869 37870 100903
rect 37904 100869 37938 100903
rect 37972 100869 38006 100903
rect 38040 100869 38074 100903
rect 38108 100869 38142 100903
rect 38176 100869 38210 100903
rect 38244 100869 38278 100903
rect 38312 100869 38346 100903
rect 38380 100869 38414 100903
rect 38448 100869 38482 100903
rect 38516 100869 38550 100903
rect 38584 100869 38618 100903
rect 38652 100869 38686 100903
rect 38720 100869 38754 100903
rect 38788 100869 38822 100903
rect 38856 100869 38890 100903
rect 38924 100869 38958 100903
rect 38992 100869 39026 100903
rect 39060 100869 39094 100903
rect 39128 100869 39162 100903
rect 39196 100869 39230 100903
rect 39264 100869 39298 100903
rect 39332 100869 39366 100903
rect 39400 100869 39434 100903
rect 39468 100869 39502 100903
rect 39536 100869 39570 100903
rect 39604 100869 39638 100903
rect 39672 100869 39706 100903
rect 39740 100869 39774 100903
rect 39808 100869 39842 100903
rect 39876 100869 39910 100903
rect 39944 100869 39978 100903
rect 40012 100869 40046 100903
rect 40080 100869 40114 100903
rect 40148 100869 40182 100903
rect 40216 100869 40250 100903
rect 40284 100869 40318 100903
rect 40352 100869 40386 100903
rect 40420 100869 40454 100903
rect 40488 100869 40522 100903
rect 40556 100869 40590 100903
rect 40624 100869 40658 100903
rect 40692 100869 40726 100903
rect 40760 100869 40794 100903
rect 40828 100869 40862 100903
rect 40896 100869 40930 100903
rect 40964 100869 40998 100903
rect 41032 100869 41066 100903
rect 41100 100869 41134 100903
rect 41168 100869 41202 100903
rect 41236 100869 41270 100903
rect 41304 100869 41338 100903
rect 41372 100869 41406 100903
rect 41440 100869 41474 100903
rect 41508 100869 41542 100903
rect 41576 100869 41610 100903
rect 41644 100869 41678 100903
rect 41712 100869 41746 100903
rect 41780 100869 41814 100903
rect 41848 100869 41882 100903
rect 41916 100869 41950 100903
rect 41984 100869 42018 100903
rect 42052 100869 42086 100903
rect 42120 100869 42154 100903
rect 42188 100869 42222 100903
rect 42256 100869 42290 100903
rect 42324 100869 42358 100903
rect 42392 100869 42426 100903
rect 42460 100869 42494 100903
rect 42528 100869 42562 100903
rect 42596 100869 42630 100903
rect 42664 100869 42698 100903
rect 42732 100869 42766 100903
rect 42800 100869 42834 100903
rect 42868 100869 42902 100903
rect 42936 100869 42970 100903
rect 43004 100869 43038 100903
rect 43072 100869 43106 100903
rect 43140 100869 43174 100903
rect 43208 100869 43242 100903
rect 43276 100869 43310 100903
rect 43344 100869 43378 100903
rect 43412 100869 43446 100903
rect 43480 100869 43514 100903
rect 43548 100869 43582 100903
rect 43616 100869 43650 100903
rect 43684 100869 43718 100903
rect 43752 100869 43786 100903
rect 43820 100869 43854 100903
rect 43888 100869 43922 100903
rect 43956 100869 43990 100903
rect 44024 100869 44058 100903
rect 44092 100869 44126 100903
rect 44160 100869 44194 100903
rect 44228 100869 44262 100903
rect 44296 100869 44330 100903
rect 44364 100869 44398 100903
rect 44432 100869 44466 100903
rect 44500 100869 44534 100903
rect 44568 100869 44602 100903
rect 44636 100869 44670 100903
rect 44704 100869 44738 100903
rect 44772 100869 44806 100903
rect 44840 100869 44874 100903
rect 44908 100869 44942 100903
rect 44976 100869 45010 100903
rect 45044 100869 45078 100903
rect 45112 100869 45146 100903
rect 45180 100869 45214 100903
rect 45248 100869 45282 100903
rect 45316 100869 45350 100903
rect 45384 100869 45418 100903
rect 45452 100869 45486 100903
rect 45520 100869 45554 100903
rect 45588 100869 45622 100903
rect 45656 100869 45690 100903
rect 45724 100869 45758 100903
rect 45792 100869 45826 100903
rect 45860 100869 45894 100903
rect 45928 100869 45962 100903
rect 45996 100869 46030 100903
rect 46064 100869 46098 100903
rect 46132 100869 46166 100903
rect 46200 100869 46234 100903
rect 46268 100869 46302 100903
rect 46336 100869 46370 100903
rect 46404 100869 46438 100903
rect 46472 100869 46506 100903
rect 46540 100869 46574 100903
rect 46608 100869 46642 100903
rect 46676 100869 46710 100903
rect 46744 100869 46778 100903
rect 46812 100869 46846 100903
rect 46880 100869 46914 100903
rect 46948 100869 46982 100903
rect 47016 100869 47050 100903
rect 47084 100869 47118 100903
rect 47152 100869 47230 100903
rect -10699 76110 -10609 76144
rect -10575 76110 -10541 76144
rect -10507 76110 -10473 76144
rect -10439 76110 -10405 76144
rect -10371 76110 -10337 76144
rect -10303 76110 -10269 76144
rect -10235 76110 -10201 76144
rect -10167 76110 -10133 76144
rect -10099 76110 -10065 76144
rect -10031 76110 -9997 76144
rect -9963 76110 -9929 76144
rect -9895 76110 -9861 76144
rect -9827 76110 -9793 76144
rect -9759 76110 -9725 76144
rect -9691 76110 -9657 76144
rect -9623 76110 -9589 76144
rect -9555 76110 -9521 76144
rect -9487 76110 -9453 76144
rect -9419 76110 -9385 76144
rect -9351 76110 -9317 76144
rect -9283 76110 -9249 76144
rect -9215 76110 -9181 76144
rect -9147 76110 -9113 76144
rect -9079 76110 -9045 76144
rect -9011 76110 -8977 76144
rect -8943 76110 -8909 76144
rect -8875 76110 -8841 76144
rect -8807 76110 -8773 76144
rect -8739 76110 -8705 76144
rect -8671 76110 -8637 76144
rect -8603 76110 -8569 76144
rect -8535 76110 -8501 76144
rect -8467 76110 -8433 76144
rect -8399 76110 -8365 76144
rect -8331 76110 -8297 76144
rect -8263 76110 -8229 76144
rect -8195 76110 -8161 76144
rect -8127 76110 -8093 76144
rect -8059 76110 -8025 76144
rect -7991 76110 -7957 76144
rect -7923 76110 -7889 76144
rect -7855 76110 -7821 76144
rect -7787 76110 -7753 76144
rect -7719 76110 -7685 76144
rect -7651 76110 -7617 76144
rect -7583 76110 -7549 76144
rect -7515 76110 -7481 76144
rect -7447 76110 -7413 76144
rect -7379 76110 -7345 76144
rect -7311 76110 -7277 76144
rect -7243 76110 -7209 76144
rect -7175 76110 -7141 76144
rect -7107 76110 -7073 76144
rect -7039 76110 -7005 76144
rect -6971 76110 -6937 76144
rect -6903 76110 -6869 76144
rect -6835 76110 -6801 76144
rect -6767 76110 -6733 76144
rect -6699 76110 -6665 76144
rect -6631 76110 -6597 76144
rect -6563 76110 -6529 76144
rect -6495 76110 -6461 76144
rect -6427 76110 -6393 76144
rect -6359 76110 -6325 76144
rect -6291 76110 -6257 76144
rect -6223 76110 -6189 76144
rect -6155 76110 -6121 76144
rect -6087 76110 -6053 76144
rect -6019 76110 -5985 76144
rect -5951 76110 -5917 76144
rect -5883 76110 -5849 76144
rect -5815 76110 -5781 76144
rect -5747 76110 -5713 76144
rect -5679 76110 -5645 76144
rect -5611 76110 -5577 76144
rect -5543 76110 -5509 76144
rect -5475 76110 -5441 76144
rect -5407 76110 -5373 76144
rect -5339 76110 -5305 76144
rect -5271 76110 -5237 76144
rect -5203 76110 -5169 76144
rect -5135 76110 -5101 76144
rect -5067 76110 -5033 76144
rect -4999 76110 -4965 76144
rect -4931 76110 -4897 76144
rect -4863 76110 -4829 76144
rect -4795 76110 -4761 76144
rect -4727 76110 -4693 76144
rect -4659 76110 -4625 76144
rect -4591 76110 -4557 76144
rect -4523 76110 -4489 76144
rect -4455 76110 -4421 76144
rect -4387 76110 -4353 76144
rect -4319 76110 -4285 76144
rect -4251 76110 -4217 76144
rect -4183 76110 -4149 76144
rect -4115 76110 -4081 76144
rect -4047 76110 -4013 76144
rect -3979 76110 -3945 76144
rect -3911 76110 -3877 76144
rect -3843 76110 -3809 76144
rect -3775 76110 -3684 76144
rect -10699 76084 -10665 76110
rect -10699 76016 -10665 76050
rect -10699 75948 -10665 75982
rect -10699 75880 -10665 75914
rect -10699 75812 -10665 75846
rect -10699 75744 -10665 75778
rect -10699 75676 -10665 75710
rect -10699 75608 -10665 75642
rect -10699 75540 -10665 75574
rect -10699 75472 -10665 75506
rect -10699 75404 -10665 75438
rect -10699 75336 -10665 75370
rect -10699 75268 -10665 75302
rect -10699 75200 -10665 75234
rect -10699 75132 -10665 75166
rect -10699 75064 -10665 75098
rect -10699 74996 -10665 75030
rect -10699 74928 -10665 74962
rect -10699 74860 -10665 74894
rect -10699 74792 -10665 74826
rect -10699 74724 -10665 74758
rect -10699 74656 -10665 74690
rect -10699 74588 -10665 74622
rect -10699 74520 -10665 74554
rect -10699 74452 -10665 74486
rect -10699 74384 -10665 74418
rect -10699 74316 -10665 74350
rect -10699 74248 -10665 74282
rect -10699 74180 -10665 74214
rect -10699 74112 -10665 74146
rect -10699 74044 -10665 74078
rect -10699 73976 -10665 74010
rect -10699 73908 -10665 73942
rect -10699 73840 -10665 73874
rect -10699 73772 -10665 73806
rect -10699 73704 -10665 73738
rect -10699 73636 -10665 73670
rect -10699 73568 -10665 73602
rect -10699 73500 -10665 73534
rect -10699 73432 -10665 73466
rect -10699 73364 -10665 73398
rect -10699 73296 -10665 73330
rect -10699 73228 -10665 73262
rect -10699 73160 -10665 73194
rect -10699 73092 -10665 73126
rect -10699 73024 -10665 73058
rect -10699 72956 -10665 72990
rect -10699 72888 -10665 72922
rect -10699 72820 -10665 72854
rect -10699 72752 -10665 72786
rect -10699 72684 -10665 72718
rect -10699 72616 -10665 72650
rect -10699 72548 -10665 72582
rect -10699 72480 -10665 72514
rect -10699 72412 -10665 72446
rect -10699 72344 -10665 72378
rect -10699 72276 -10665 72310
rect -10699 72208 -10665 72242
rect -10699 72140 -10665 72174
rect -10699 72072 -10665 72106
rect -10699 72004 -10665 72038
rect -10699 71936 -10665 71970
rect -10699 71868 -10665 71902
rect -10699 71800 -10665 71834
rect -10699 71732 -10665 71766
rect -10699 71664 -10665 71698
rect -10699 71596 -10665 71630
rect -10699 71528 -10665 71562
rect -10699 71460 -10665 71494
rect -10699 71392 -10665 71426
rect -10699 71324 -10665 71358
rect -10699 71256 -10665 71290
rect -10699 71188 -10665 71222
rect -10699 71120 -10665 71154
rect -10699 71052 -10665 71086
rect -10699 70984 -10665 71018
rect -10699 70916 -10665 70950
rect -10699 70848 -10665 70882
rect -10699 70780 -10665 70814
rect -10699 70712 -10665 70746
rect -10699 70644 -10665 70678
rect -10699 70576 -10665 70610
rect -10699 70508 -10665 70542
rect -10699 70440 -10665 70474
rect -10699 70372 -10665 70406
rect -10699 70304 -10665 70338
rect -10699 70236 -10665 70270
rect -10699 70168 -10665 70202
rect -10699 70100 -10665 70134
rect -10699 70032 -10665 70066
rect -10699 69964 -10665 69998
rect -10699 69896 -10665 69930
rect -10699 69828 -10665 69862
rect -10699 69760 -10665 69794
rect -10699 69692 -10665 69726
rect -10699 69624 -10665 69658
rect -10699 69556 -10665 69590
rect -10699 69488 -10665 69522
rect -10699 69420 -10665 69454
rect -10699 69352 -10665 69386
rect -10699 69284 -10665 69318
rect -10699 69216 -10665 69250
rect -10699 69148 -10665 69182
rect -10699 69080 -10665 69114
rect -10699 69012 -10665 69046
rect -10699 68944 -10665 68978
rect -10699 68876 -10665 68910
rect -10699 68808 -10665 68842
rect -10699 68740 -10665 68774
rect -10699 68672 -10665 68706
rect -10699 68604 -10665 68638
rect -10699 68536 -10665 68570
rect -10699 68468 -10665 68502
rect -10699 68400 -10665 68434
rect -10699 68332 -10665 68366
rect -10699 68264 -10665 68298
rect -10699 68196 -10665 68230
rect -10699 68128 -10665 68162
rect -10699 68060 -10665 68094
rect -10699 67992 -10665 68026
rect -10699 67924 -10665 67958
rect -10699 67856 -10665 67890
rect -10699 67788 -10665 67822
rect -10699 67720 -10665 67754
rect -10699 67652 -10665 67686
rect -10699 67584 -10665 67618
rect -10699 67516 -10665 67550
rect -10699 67448 -10665 67482
rect -10699 67380 -10665 67414
rect -10699 67312 -10665 67346
rect -10699 67244 -10665 67278
rect -10699 67176 -10665 67210
rect -10699 67108 -10665 67142
rect -10699 67040 -10665 67074
rect -10699 66972 -10665 67006
rect -10699 66904 -10665 66938
rect -10699 66836 -10665 66870
rect -10699 66768 -10665 66802
rect -10699 66700 -10665 66734
rect -10699 66632 -10665 66666
rect -10699 66564 -10665 66598
rect -10699 66496 -10665 66530
rect -10699 66428 -10665 66462
rect -10699 66360 -10665 66394
rect -10699 66292 -10665 66326
rect -10699 66224 -10665 66258
rect -10699 66156 -10665 66190
rect -10699 66088 -10665 66122
rect -10699 66020 -10665 66054
rect -10699 65952 -10665 65986
rect -10699 65884 -10665 65918
rect -10699 65816 -10665 65850
rect -10699 65748 -10665 65782
rect -10699 65680 -10665 65714
rect -10699 65612 -10665 65646
rect -10699 65544 -10665 65578
rect -10699 65476 -10665 65510
rect -10699 65408 -10665 65442
rect -10699 65340 -10665 65374
rect -10699 65272 -10665 65306
rect -10699 65204 -10665 65238
rect -10699 65136 -10665 65170
rect -10699 65068 -10665 65102
rect -10699 65000 -10665 65034
rect -10699 64932 -10665 64966
rect -10699 64864 -10665 64898
rect -10699 64796 -10665 64830
rect -10699 64728 -10665 64762
rect -10699 64660 -10665 64694
rect -10699 64592 -10665 64626
rect -10699 64524 -10665 64558
rect -10699 64456 -10665 64490
rect -10699 64388 -10665 64422
rect -10699 64320 -10665 64354
rect -10699 64252 -10665 64286
rect -10699 64184 -10665 64218
rect -10699 64120 -10665 64150
rect -3718 76056 -3684 76110
rect -3718 75988 -3684 76022
rect -3718 75920 -3684 75954
rect -3718 75852 -3684 75886
rect -3718 75784 -3684 75818
rect -3718 75716 -3684 75750
rect -3718 75648 -3684 75682
rect -3718 75580 -3684 75614
rect -3718 75512 -3684 75546
rect -3718 75444 -3684 75478
rect -3718 75376 -3684 75410
rect -3718 75308 -3684 75342
rect -3718 75240 -3684 75274
rect -3718 75172 -3684 75206
rect -3718 75104 -3684 75138
rect -3718 75036 -3684 75070
rect -3718 74968 -3684 75002
rect -3718 74900 -3684 74934
rect -3718 74832 -3684 74866
rect -3718 74764 -3684 74798
rect -3718 74696 -3684 74730
rect -3718 74628 -3684 74662
rect -3718 74560 -3684 74594
rect -3718 74492 -3684 74526
rect -3718 74424 -3684 74458
rect -3718 74356 -3684 74390
rect -3718 74288 -3684 74322
rect -3718 74220 -3684 74254
rect -3718 74152 -3684 74186
rect -3718 74084 -3684 74118
rect -3718 74016 -3684 74050
rect -3718 73948 -3684 73982
rect -3718 73880 -3684 73914
rect -3718 73812 -3684 73846
rect -3718 73744 -3684 73778
rect -3718 73676 -3684 73710
rect -3718 73608 -3684 73642
rect -3718 73540 -3684 73574
rect -3718 73472 -3684 73506
rect -3718 73404 -3684 73438
rect -3718 73336 -3684 73370
rect -3718 73268 -3684 73302
rect -3718 73200 -3684 73234
rect -3718 73132 -3684 73166
rect -3718 73064 -3684 73098
rect -3718 72996 -3684 73030
rect -3718 72928 -3684 72962
rect -3718 72860 -3684 72894
rect -3718 72792 -3684 72826
rect -3718 72724 -3684 72758
rect -3718 72656 -3684 72690
rect -3718 72588 -3684 72622
rect -3718 72520 -3684 72554
rect -3718 72452 -3684 72486
rect -3718 72384 -3684 72418
rect -3718 72316 -3684 72350
rect -3718 72248 -3684 72282
rect -3718 72180 -3684 72214
rect -3718 72112 -3684 72146
rect -3718 72044 -3684 72078
rect -3718 71976 -3684 72010
rect -3718 71908 -3684 71942
rect -3718 71840 -3684 71874
rect -3718 71772 -3684 71806
rect -3718 71704 -3684 71738
rect -3718 71636 -3684 71670
rect -3718 71568 -3684 71602
rect -3718 71500 -3684 71534
rect -3718 71432 -3684 71466
rect -3718 71364 -3684 71398
rect -3718 71296 -3684 71330
rect -3718 71228 -3684 71262
rect -3718 71160 -3684 71194
rect -3718 71092 -3684 71126
rect -3718 71024 -3684 71058
rect -3718 70956 -3684 70990
rect -3718 70888 -3684 70922
rect -3718 70820 -3684 70854
rect -3718 70752 -3684 70786
rect -3718 70684 -3684 70718
rect -3718 70616 -3684 70650
rect -3718 70548 -3684 70582
rect -3718 70480 -3684 70514
rect -3718 70412 -3684 70446
rect -3718 70344 -3684 70378
rect -3718 70276 -3684 70310
rect -3718 70208 -3684 70242
rect -3718 70140 -3684 70174
rect -3718 70072 -3684 70106
rect -3718 70004 -3684 70038
rect -3718 69936 -3684 69970
rect -3718 69868 -3684 69902
rect -3718 69800 -3684 69834
rect -3718 69732 -3684 69766
rect -3718 69664 -3684 69698
rect -3718 69596 -3684 69630
rect -3718 69528 -3684 69562
rect -3718 69460 -3684 69494
rect -3718 69392 -3684 69426
rect -3718 69324 -3684 69358
rect -3718 69256 -3684 69290
rect -3718 69188 -3684 69222
rect -3718 69120 -3684 69154
rect -3718 69052 -3684 69086
rect -3718 68984 -3684 69018
rect -3718 68916 -3684 68950
rect -3718 68848 -3684 68882
rect -3718 68780 -3684 68814
rect -3718 68712 -3684 68746
rect -3718 68644 -3684 68678
rect -3718 68576 -3684 68610
rect -3718 68508 -3684 68542
rect -3718 68440 -3684 68474
rect -3718 68372 -3684 68406
rect -3718 68304 -3684 68338
rect -3718 68236 -3684 68270
rect -3718 68168 -3684 68202
rect -3718 68100 -3684 68134
rect -3718 68032 -3684 68066
rect -3718 67964 -3684 67998
rect -3718 67896 -3684 67930
rect -3718 67828 -3684 67862
rect -3718 67760 -3684 67794
rect -3718 67692 -3684 67726
rect -3718 67624 -3684 67658
rect -3718 67556 -3684 67590
rect -3718 67488 -3684 67522
rect -3718 67420 -3684 67454
rect -3718 67352 -3684 67386
rect -3718 67284 -3684 67318
rect -3718 67216 -3684 67250
rect -3718 67148 -3684 67182
rect -3718 67080 -3684 67114
rect -3718 67012 -3684 67046
rect -3718 66944 -3684 66978
rect -3718 66876 -3684 66910
rect -3718 66808 -3684 66842
rect -3718 66740 -3684 66774
rect -3718 66672 -3684 66706
rect -3718 66604 -3684 66638
rect -3718 66536 -3684 66570
rect -3718 66468 -3684 66502
rect -3718 66400 -3684 66434
rect -3718 66332 -3684 66366
rect -3718 66264 -3684 66298
rect -3718 66196 -3684 66230
rect -3718 66128 -3684 66162
rect -3718 66060 -3684 66094
rect -3718 65992 -3684 66026
rect -3718 65924 -3684 65958
rect -3718 65856 -3684 65890
rect -3718 65788 -3684 65822
rect -3718 65720 -3684 65754
rect -3718 65652 -3684 65686
rect -3718 65584 -3684 65618
rect -3718 65516 -3684 65550
rect -3718 65448 -3684 65482
rect -3718 65380 -3684 65414
rect -3718 65312 -3684 65346
rect -3718 65244 -3684 65278
rect -3718 65176 -3684 65210
rect -3718 65108 -3684 65142
rect -3718 65040 -3684 65074
rect -3718 64972 -3684 65006
rect -3718 64904 -3684 64938
rect -3718 64836 -3684 64870
rect -3718 64768 -3684 64802
rect -3718 64700 -3684 64734
rect -3718 64632 -3684 64666
rect -3718 64564 -3684 64598
rect -3718 64496 -3684 64530
rect -3718 64428 -3684 64462
rect -3718 64360 -3684 64394
rect -3718 64292 -3684 64326
rect -3718 64224 -3684 64258
rect -3718 64156 -3684 64190
rect -10699 64086 -10624 64120
rect -10590 64086 -10556 64120
rect -10522 64086 -10488 64120
rect -10454 64086 -10420 64120
rect -10386 64086 -10352 64120
rect -10318 64086 -10284 64120
rect -10250 64086 -10216 64120
rect -10182 64086 -10148 64120
rect -10114 64086 -10080 64120
rect -10046 64086 -10012 64120
rect -9978 64086 -9944 64120
rect -9910 64086 -9876 64120
rect -9842 64086 -9808 64120
rect -9774 64086 -9740 64120
rect -9706 64086 -9672 64120
rect -9638 64086 -9604 64120
rect -9570 64086 -9536 64120
rect -9502 64086 -9468 64120
rect -9434 64086 -9400 64120
rect -9366 64086 -9332 64120
rect -9298 64086 -9264 64120
rect -9230 64086 -9196 64120
rect -9162 64086 -9128 64120
rect -9094 64086 -9060 64120
rect -9026 64086 -8992 64120
rect -8958 64086 -8924 64120
rect -8890 64086 -8856 64120
rect -8822 64086 -8788 64120
rect -8754 64086 -8720 64120
rect -8686 64086 -8652 64120
rect -8618 64086 -8584 64120
rect -8550 64086 -8516 64120
rect -8482 64086 -8448 64120
rect -8414 64086 -8380 64120
rect -8346 64086 -8312 64120
rect -8278 64086 -8244 64120
rect -8210 64086 -8176 64120
rect -8142 64086 -8108 64120
rect -8074 64086 -8040 64120
rect -8006 64086 -7972 64120
rect -7938 64086 -7904 64120
rect -7870 64086 -7836 64120
rect -7802 64086 -7768 64120
rect -7734 64086 -7700 64120
rect -7666 64086 -7632 64120
rect -7598 64086 -7564 64120
rect -7530 64086 -7496 64120
rect -7462 64086 -7428 64120
rect -7394 64086 -7360 64120
rect -7326 64086 -7292 64120
rect -7258 64086 -7173 64120
rect -7207 64059 -7173 64086
rect -7207 63991 -7173 64025
rect -7207 63923 -7173 63957
rect -7207 63855 -7173 63889
rect -7207 63787 -7173 63821
rect -7207 63719 -7173 63753
rect -7207 63651 -7173 63685
rect -7207 63583 -7173 63617
rect -7207 63515 -7173 63549
rect -7207 63447 -7173 63481
rect -7207 63379 -7173 63413
rect -7207 63311 -7173 63345
rect -7207 63243 -7173 63277
rect -7207 63175 -7173 63209
rect -7207 63107 -7173 63141
rect -7207 63039 -7173 63073
rect -7207 62971 -7173 63005
rect -7207 62903 -7173 62937
rect -7207 62835 -7173 62869
rect -7207 62767 -7173 62801
rect -7207 62699 -7173 62733
rect -7207 62631 -7173 62665
rect -7207 62563 -7173 62597
rect -7207 62495 -7173 62529
rect -7207 62427 -7173 62461
rect -7207 62359 -7173 62393
rect -7207 62291 -7173 62325
rect -7207 62223 -7173 62257
rect -7207 62155 -7173 62189
rect -7207 62087 -7173 62121
rect -7207 62019 -7173 62053
rect -7207 61951 -7173 61985
rect -7207 61883 -7173 61917
rect -7207 61815 -7173 61849
rect -7207 61747 -7173 61781
rect -7207 61679 -7173 61713
rect -7207 61611 -7173 61645
rect -7207 61543 -7173 61577
rect -7207 61475 -7173 61509
rect -7207 61407 -7173 61441
rect -7207 61339 -7173 61373
rect -7207 61271 -7173 61305
rect -7207 61203 -7173 61237
rect -7207 61135 -7173 61169
rect -7207 61067 -7173 61101
rect -7207 60999 -7173 61033
rect -7207 60931 -7173 60965
rect -7207 60863 -7173 60897
rect -7207 60795 -7173 60829
rect -7207 60727 -7173 60761
rect -7207 60659 -7173 60693
rect -7207 60591 -7173 60625
rect -7207 60523 -7173 60557
rect -7207 60455 -7173 60489
rect -7207 60387 -7173 60421
rect -7207 60319 -7173 60353
rect -7207 60251 -7173 60285
rect -7207 60183 -7173 60217
rect -7207 60115 -7173 60149
rect -7207 60047 -7173 60081
rect -7207 59979 -7173 60013
rect -7207 59911 -7173 59945
rect -7207 59843 -7173 59877
rect -7207 59775 -7173 59809
rect -7207 59707 -7173 59741
rect -7207 59639 -7173 59673
rect -7207 59571 -7173 59605
rect -7207 59503 -7173 59537
rect -7207 59435 -7173 59469
rect -7207 59367 -7173 59401
rect -7207 59299 -7173 59333
rect -7207 59231 -7173 59265
rect -7207 59163 -7173 59197
rect -7207 59095 -7173 59129
rect -7207 59027 -7173 59061
rect -7207 58959 -7173 58993
rect -7207 58891 -7173 58925
rect -7207 58823 -7173 58857
rect -7207 58755 -7173 58789
rect -7207 58687 -7173 58721
rect -7207 58619 -7173 58653
rect -7207 58551 -7173 58585
rect -7207 58483 -7173 58517
rect -7207 58415 -7173 58449
rect -7207 58347 -7173 58381
rect -7207 58279 -7173 58313
rect -7207 58211 -7173 58245
rect -7207 58143 -7173 58177
rect -7207 58075 -7173 58109
rect -7207 58007 -7173 58041
rect -7207 57939 -7173 57973
rect -7207 57871 -7173 57905
rect -7207 57803 -7173 57837
rect -7207 57735 -7173 57769
rect -7207 57667 -7173 57701
rect -7207 57599 -7173 57633
rect -7207 57531 -7173 57565
rect -7207 57463 -7173 57497
rect -7207 57395 -7173 57429
rect -7207 57327 -7173 57361
rect -7207 57259 -7173 57293
rect -7207 57191 -7173 57225
rect -7207 57123 -7173 57157
rect -7207 57055 -7173 57089
rect -7207 56987 -7173 57021
rect -7207 56919 -7173 56953
rect -7207 56851 -7173 56885
rect -7207 56783 -7173 56817
rect -7207 56715 -7173 56749
rect -7207 56647 -7173 56681
rect -7207 56579 -7173 56613
rect -7207 56511 -7173 56545
rect -7207 56443 -7173 56477
rect -7207 56375 -7173 56409
rect -7207 56304 -7173 56341
rect -10699 56270 -10614 56304
rect -10580 56270 -10546 56304
rect -10512 56270 -10478 56304
rect -10444 56270 -10410 56304
rect -10376 56270 -10342 56304
rect -10308 56270 -10274 56304
rect -10240 56270 -10206 56304
rect -10172 56270 -10138 56304
rect -10104 56270 -10070 56304
rect -10036 56270 -10002 56304
rect -9968 56270 -9934 56304
rect -9900 56270 -9866 56304
rect -9832 56270 -9798 56304
rect -9764 56270 -9730 56304
rect -9696 56270 -9662 56304
rect -9628 56270 -9594 56304
rect -9560 56270 -9526 56304
rect -9492 56270 -9458 56304
rect -9424 56270 -9390 56304
rect -9356 56270 -9322 56304
rect -9288 56270 -9254 56304
rect -9220 56270 -9186 56304
rect -9152 56270 -9118 56304
rect -9084 56270 -9050 56304
rect -9016 56270 -8982 56304
rect -8948 56270 -8914 56304
rect -8880 56270 -8846 56304
rect -8812 56270 -8778 56304
rect -8744 56270 -8710 56304
rect -8676 56270 -8642 56304
rect -8608 56270 -8574 56304
rect -8540 56270 -8506 56304
rect -8472 56270 -8438 56304
rect -8404 56270 -8370 56304
rect -8336 56270 -8302 56304
rect -8268 56270 -8234 56304
rect -8200 56270 -8166 56304
rect -8132 56270 -8098 56304
rect -8064 56270 -8030 56304
rect -7996 56270 -7962 56304
rect -7928 56270 -7894 56304
rect -7860 56270 -7826 56304
rect -7792 56270 -7758 56304
rect -7724 56270 -7690 56304
rect -7656 56270 -7622 56304
rect -7588 56270 -7554 56304
rect -7520 56270 -7486 56304
rect -7452 56270 -7418 56304
rect -7384 56270 -7350 56304
rect -7316 56270 -7282 56304
rect -7248 56270 -7173 56304
rect -3718 64088 -3684 64122
rect -3718 64020 -3684 64054
rect -3718 63952 -3684 63986
rect -3718 63884 -3684 63918
rect -3718 63816 -3684 63850
rect -3718 63748 -3684 63782
rect -3718 63680 -3684 63714
rect -3718 63612 -3684 63646
rect -3718 63544 -3684 63578
rect -3718 63476 -3684 63510
rect -3718 63408 -3684 63442
rect -3718 63340 -3684 63374
rect -3718 63272 -3684 63306
rect -3718 63204 -3684 63238
rect -3718 63136 -3684 63170
rect -3718 63068 -3684 63102
rect -3718 63000 -3684 63034
rect -3718 62932 -3684 62966
rect -3718 62864 -3684 62898
rect -3718 62796 -3684 62830
rect -3718 62728 -3684 62762
rect -3718 62660 -3684 62694
rect -3718 62592 -3684 62626
rect -3718 62524 -3684 62558
rect -3718 62456 -3684 62490
rect -3718 62388 -3684 62422
rect -3718 62320 -3684 62354
rect -3718 62252 -3684 62286
rect -3718 62184 -3684 62218
rect -3718 62116 -3684 62150
rect -3718 62048 -3684 62082
rect 59104 74772 59191 74806
rect 59225 74772 59259 74806
rect 59293 74772 59327 74806
rect 59361 74772 59395 74806
rect 59429 74772 59463 74806
rect 59497 74772 59531 74806
rect 59565 74772 59599 74806
rect 59633 74772 59667 74806
rect 59701 74772 59735 74806
rect 59769 74772 59803 74806
rect 59837 74772 59871 74806
rect 59905 74772 59939 74806
rect 59973 74772 60007 74806
rect 60041 74772 60075 74806
rect 60109 74772 60143 74806
rect 60177 74772 60211 74806
rect 60245 74772 60279 74806
rect 60313 74772 60347 74806
rect 60381 74772 60415 74806
rect 60449 74772 60483 74806
rect 60517 74772 60551 74806
rect 60585 74772 60619 74806
rect 60653 74772 60687 74806
rect 60721 74772 60755 74806
rect 60789 74772 60823 74806
rect 60857 74772 60891 74806
rect 60925 74772 60959 74806
rect 60993 74772 61027 74806
rect 61061 74772 61095 74806
rect 61129 74772 61163 74806
rect 61197 74772 61231 74806
rect 61265 74772 61299 74806
rect 61333 74772 61367 74806
rect 61401 74772 61435 74806
rect 61469 74772 61503 74806
rect 61537 74772 61571 74806
rect 61605 74772 61639 74806
rect 61673 74772 61707 74806
rect 61741 74772 61775 74806
rect 61809 74772 61843 74806
rect 61877 74772 61911 74806
rect 61945 74772 61979 74806
rect 62013 74772 62047 74806
rect 62081 74772 62115 74806
rect 62149 74772 62183 74806
rect 62217 74772 62251 74806
rect 62285 74772 62319 74806
rect 62353 74772 62387 74806
rect 62421 74772 62455 74806
rect 62489 74772 62523 74806
rect 62557 74772 62591 74806
rect 62625 74772 62659 74806
rect 62693 74772 62727 74806
rect 62761 74772 62795 74806
rect 62829 74772 62863 74806
rect 62897 74772 62931 74806
rect 62965 74772 62999 74806
rect 63033 74772 63067 74806
rect 63101 74772 63135 74806
rect 63169 74772 63203 74806
rect 63237 74772 63271 74806
rect 63305 74772 63339 74806
rect 63373 74772 63407 74806
rect 63441 74772 63475 74806
rect 63509 74772 63543 74806
rect 63577 74772 63611 74806
rect 63645 74772 63679 74806
rect 63713 74772 63747 74806
rect 63781 74772 63815 74806
rect 63849 74772 63883 74806
rect 63917 74772 63951 74806
rect 63985 74772 64019 74806
rect 64053 74772 64087 74806
rect 64121 74772 64155 74806
rect 64189 74772 64223 74806
rect 64257 74772 64291 74806
rect 64325 74772 64359 74806
rect 64393 74772 64427 74806
rect 64461 74772 64495 74806
rect 64529 74772 64563 74806
rect 64597 74772 64631 74806
rect 64665 74772 64699 74806
rect 64733 74772 64767 74806
rect 64801 74772 64835 74806
rect 64869 74772 64903 74806
rect 64937 74772 64971 74806
rect 65005 74772 65039 74806
rect 65073 74772 65107 74806
rect 65141 74772 65175 74806
rect 65209 74772 65243 74806
rect 65277 74772 65311 74806
rect 65345 74772 65379 74806
rect 65413 74772 65447 74806
rect 65481 74772 65515 74806
rect 65549 74772 65583 74806
rect 65617 74772 65651 74806
rect 65685 74772 65719 74806
rect 65753 74772 65787 74806
rect 65821 74772 65855 74806
rect 65889 74772 65923 74806
rect 65957 74772 65991 74806
rect 66025 74772 66059 74806
rect 66093 74772 66127 74806
rect 66161 74772 66195 74806
rect 66229 74772 66263 74806
rect 66297 74772 66331 74806
rect 66365 74772 66399 74806
rect 66433 74772 66467 74806
rect 66501 74772 66535 74806
rect 66569 74772 66603 74806
rect 66637 74772 66671 74806
rect 66705 74772 66739 74806
rect 66773 74772 66807 74806
rect 66841 74772 66875 74806
rect 66909 74772 66943 74806
rect 66977 74772 67011 74806
rect 67045 74772 67079 74806
rect 67113 74772 67147 74806
rect 67181 74772 67215 74806
rect 67249 74772 67283 74806
rect 67317 74772 67351 74806
rect 67385 74772 67419 74806
rect 67453 74772 67487 74806
rect 67521 74772 67555 74806
rect 67589 74772 67623 74806
rect 67657 74772 67691 74806
rect 67725 74772 67759 74806
rect 67793 74772 67827 74806
rect 67861 74772 67895 74806
rect 67929 74772 67963 74806
rect 67997 74772 68031 74806
rect 68065 74772 68099 74806
rect 68133 74772 68167 74806
rect 68201 74772 68235 74806
rect 68269 74772 68303 74806
rect 68337 74772 68371 74806
rect 68405 74772 68439 74806
rect 68473 74772 68507 74806
rect 68541 74772 68575 74806
rect 68609 74772 68643 74806
rect 68677 74772 68711 74806
rect 68745 74772 68779 74806
rect 68813 74772 68847 74806
rect 68881 74772 68915 74806
rect 68949 74772 68983 74806
rect 69017 74772 69051 74806
rect 69085 74772 69119 74806
rect 69153 74772 69187 74806
rect 69221 74772 69255 74806
rect 69289 74772 69323 74806
rect 69357 74772 69391 74806
rect 69425 74772 69459 74806
rect 69493 74772 69527 74806
rect 69561 74772 69595 74806
rect 69629 74772 69663 74806
rect 69697 74772 69731 74806
rect 69765 74772 69799 74806
rect 69833 74772 69867 74806
rect 69901 74772 69935 74806
rect 69969 74772 70003 74806
rect 70037 74772 70071 74806
rect 70105 74772 70139 74806
rect 70173 74772 70207 74806
rect 70241 74772 70275 74806
rect 70309 74772 70343 74806
rect 70377 74772 70411 74806
rect 70445 74772 70479 74806
rect 70513 74772 70547 74806
rect 70581 74772 70615 74806
rect 70649 74772 70683 74806
rect 70717 74772 70751 74806
rect 70785 74772 70872 74806
rect 59104 74745 59138 74772
rect 59104 74677 59138 74711
rect 59104 74609 59138 74643
rect 59104 74541 59138 74575
rect 59104 74473 59138 74507
rect 59104 74405 59138 74439
rect 59104 74337 59138 74371
rect 59104 74269 59138 74303
rect 59104 74201 59138 74235
rect 59104 74133 59138 74167
rect 59104 74065 59138 74099
rect 59104 73997 59138 74031
rect 59104 73929 59138 73963
rect 59104 73861 59138 73895
rect 59104 73793 59138 73827
rect 59104 73725 59138 73759
rect 59104 73657 59138 73691
rect 59104 73589 59138 73623
rect 59104 73521 59138 73555
rect 59104 73453 59138 73487
rect 59104 73385 59138 73419
rect 59104 73317 59138 73351
rect 59104 73249 59138 73283
rect 59104 73181 59138 73215
rect 59104 73113 59138 73147
rect 59104 73045 59138 73079
rect 59104 72977 59138 73011
rect 59104 72909 59138 72943
rect 59104 72841 59138 72875
rect 59104 72773 59138 72807
rect 59104 72705 59138 72739
rect 59104 72637 59138 72671
rect 59104 72569 59138 72603
rect 59104 72501 59138 72535
rect 59104 72433 59138 72467
rect 59104 72365 59138 72399
rect 59104 72297 59138 72331
rect 59104 72229 59138 72263
rect 59104 72161 59138 72195
rect 59104 72093 59138 72127
rect 59104 72025 59138 72059
rect 59104 71957 59138 71991
rect 59104 71889 59138 71923
rect 59104 71821 59138 71855
rect 59104 71753 59138 71787
rect 59104 71685 59138 71719
rect 59104 71617 59138 71651
rect 59104 71549 59138 71583
rect 59104 71481 59138 71515
rect 59104 71413 59138 71447
rect 59104 71345 59138 71379
rect 59104 71277 59138 71311
rect 59104 71209 59138 71243
rect 59104 71141 59138 71175
rect 59104 71073 59138 71107
rect 59104 71005 59138 71039
rect 59104 70937 59138 70971
rect 59104 70869 59138 70903
rect 59104 70801 59138 70835
rect 59104 70733 59138 70767
rect 59104 70665 59138 70699
rect 59104 70597 59138 70631
rect 59104 70529 59138 70563
rect 59104 70461 59138 70495
rect 59104 70393 59138 70427
rect 59104 70325 59138 70359
rect 59104 70257 59138 70291
rect 59104 70189 59138 70223
rect 59104 70121 59138 70155
rect 59104 70053 59138 70087
rect 59104 69985 59138 70019
rect 59104 69917 59138 69951
rect 59104 69849 59138 69883
rect 59104 69781 59138 69815
rect 59104 69713 59138 69747
rect 59104 69645 59138 69679
rect 59104 69577 59138 69611
rect 59104 69509 59138 69543
rect 59104 69441 59138 69475
rect 59104 69373 59138 69407
rect 59104 69305 59138 69339
rect 59104 69237 59138 69271
rect 59104 69169 59138 69203
rect 59104 69101 59138 69135
rect 59104 69033 59138 69067
rect 59104 68965 59138 68999
rect 59104 68897 59138 68931
rect 59104 68829 59138 68863
rect 59104 68761 59138 68795
rect 59104 68693 59138 68727
rect 59104 68625 59138 68659
rect 59104 68557 59138 68591
rect 59104 68489 59138 68523
rect 59104 68421 59138 68455
rect 59104 68353 59138 68387
rect 59104 68285 59138 68319
rect 59104 68217 59138 68251
rect 59104 68149 59138 68183
rect 59104 68081 59138 68115
rect 59104 68013 59138 68047
rect 59104 67945 59138 67979
rect 59104 67877 59138 67911
rect 59104 67809 59138 67843
rect 59104 67741 59138 67775
rect 59104 67673 59138 67707
rect 59104 67605 59138 67639
rect 59104 67537 59138 67571
rect 59104 67469 59138 67503
rect 59104 67401 59138 67435
rect 59104 67333 59138 67367
rect 59104 67265 59138 67299
rect 59104 67197 59138 67231
rect 59104 67129 59138 67163
rect 59104 67061 59138 67095
rect 59104 66993 59138 67027
rect 59104 66925 59138 66959
rect 59104 66857 59138 66891
rect 59104 66789 59138 66823
rect 59104 66721 59138 66755
rect 59104 66653 59138 66687
rect 59104 66585 59138 66619
rect 59104 66517 59138 66551
rect 59104 66449 59138 66483
rect 59104 66381 59138 66415
rect 59104 66313 59138 66347
rect 59104 66245 59138 66279
rect 59104 66177 59138 66211
rect 59104 66109 59138 66143
rect 59104 66041 59138 66075
rect 59104 65973 59138 66007
rect 59104 65905 59138 65939
rect 59104 65837 59138 65871
rect 59104 65769 59138 65803
rect 59104 65701 59138 65735
rect 59104 65633 59138 65667
rect 59104 65565 59138 65599
rect 59104 65497 59138 65531
rect 59104 65429 59138 65463
rect 59104 65361 59138 65395
rect 59104 65293 59138 65327
rect 59104 65225 59138 65259
rect 59104 65157 59138 65191
rect 59104 65089 59138 65123
rect 59104 65021 59138 65055
rect 59104 64953 59138 64987
rect 59104 64885 59138 64919
rect 59104 64817 59138 64851
rect 59104 64749 59138 64783
rect 59104 64681 59138 64715
rect 59104 64613 59138 64647
rect 59104 64545 59138 64579
rect 59104 64477 59138 64511
rect 59104 64409 59138 64443
rect 59104 64341 59138 64375
rect 59104 64273 59138 64307
rect 59104 64205 59138 64239
rect 59104 64137 59138 64171
rect 59104 64069 59138 64103
rect 59104 64001 59138 64035
rect 59104 63933 59138 63967
rect 59104 63865 59138 63899
rect 59104 63797 59138 63831
rect 59104 63729 59138 63763
rect 59104 63661 59138 63695
rect 59104 63593 59138 63627
rect 59104 63525 59138 63559
rect 59104 63457 59138 63491
rect 59104 63389 59138 63423
rect 59104 63321 59138 63355
rect 59104 63253 59138 63287
rect 59104 63185 59138 63219
rect 59104 63117 59138 63151
rect 59104 63049 59138 63083
rect 59104 62981 59138 63015
rect 59104 62913 59138 62947
rect 59104 62845 59138 62879
rect 59104 62777 59138 62811
rect 59104 62709 59138 62743
rect 59104 62641 59138 62675
rect 59104 62573 59138 62607
rect 59104 62505 59138 62539
rect 59104 62437 59138 62471
rect 59104 62369 59138 62403
rect 59104 62301 59138 62335
rect 59104 62233 59138 62267
rect 59104 62165 59138 62199
rect 59104 62097 59138 62131
rect -3718 61980 -3684 62014
rect -3718 61912 -3684 61946
rect -3718 61844 -3684 61878
rect -3718 61776 -3684 61810
rect -3718 61708 -3684 61742
rect -3718 61640 -3684 61674
rect -3718 61572 -3684 61606
rect -3718 61504 -3684 61538
rect -3718 61436 -3684 61470
rect -3718 61368 -3684 61402
rect -3718 61300 -3684 61334
rect -3718 61232 -3684 61266
rect -3718 61164 -3684 61198
rect -3718 61096 -3684 61130
rect -3718 61028 -3684 61062
rect -3718 60960 -3684 60994
rect -3718 60892 -3684 60926
rect -3718 60824 -3684 60858
rect -3718 60756 -3684 60790
rect -3718 60688 -3684 60722
rect -3718 60620 -3684 60654
rect -3718 60552 -3684 60586
rect -3718 60484 -3684 60518
rect -3718 60416 -3684 60450
rect -3718 60348 -3684 60382
rect -3718 60280 -3684 60314
rect -3718 60212 -3684 60246
rect -3718 60144 -3684 60178
rect -3718 60076 -3684 60110
rect -3718 60008 -3684 60042
rect -3718 59940 -3684 59974
rect -3718 59872 -3684 59906
rect -3718 59804 -3684 59838
rect -3718 59736 -3684 59770
rect -3718 59668 -3684 59702
rect -3718 59600 -3684 59634
rect -3718 59532 -3684 59566
rect -3718 59464 -3684 59498
rect -3718 59396 -3684 59430
rect -3718 59328 -3684 59362
rect -3718 59260 -3684 59294
rect -3718 59192 -3684 59226
rect -3718 59124 -3684 59158
rect -3718 59056 -3684 59090
rect -3718 58988 -3684 59022
rect -3718 58920 -3684 58954
rect -3718 58852 -3684 58886
rect -3718 58784 -3684 58818
rect -3718 58716 -3684 58750
rect -3718 58648 -3684 58682
rect -3718 58580 -3684 58614
rect -3718 58512 -3684 58546
rect -3718 58444 -3684 58478
rect -3718 58376 -3684 58410
rect 50456 62006 50530 62040
rect 50564 62006 50598 62040
rect 50632 62006 50666 62040
rect 50700 62006 50734 62040
rect 50768 62006 50802 62040
rect 50836 62006 50870 62040
rect 50904 62006 50938 62040
rect 50972 62006 51006 62040
rect 51040 62006 51074 62040
rect 51108 62006 51142 62040
rect 51176 62006 51210 62040
rect 51244 62006 51278 62040
rect 51312 62006 51346 62040
rect 51380 62006 51414 62040
rect 51448 62006 51482 62040
rect 51516 62006 51550 62040
rect 51584 62006 51618 62040
rect 51652 62006 51686 62040
rect 51720 62006 51754 62040
rect 51788 62006 51822 62040
rect 51856 62006 51890 62040
rect 51924 62006 51958 62040
rect 51992 62006 52026 62040
rect 52060 62006 52094 62040
rect 52128 62006 52162 62040
rect 52196 62006 52230 62040
rect 52264 62006 52298 62040
rect 52332 62006 52366 62040
rect 52400 62006 52434 62040
rect 52468 62006 52502 62040
rect 52536 62006 52570 62040
rect 52604 62006 52638 62040
rect 52672 62006 52706 62040
rect 52740 62006 52774 62040
rect 52808 62006 52842 62040
rect 52876 62006 52910 62040
rect 52944 62006 52978 62040
rect 53012 62006 53046 62040
rect 53080 62006 53114 62040
rect 53148 62006 53182 62040
rect 53216 62006 53250 62040
rect 53284 62006 53318 62040
rect 53352 62006 53386 62040
rect 53420 62006 53454 62040
rect 53488 62006 53522 62040
rect 53556 62006 53590 62040
rect 53624 62006 53658 62040
rect 53692 62006 53726 62040
rect 53760 62006 53794 62040
rect 53828 62006 53862 62040
rect 53896 62006 53930 62040
rect 53964 62006 53998 62040
rect 54032 62006 54066 62040
rect 54100 62006 54134 62040
rect 54168 62006 54202 62040
rect 54236 62006 54270 62040
rect 54304 62006 54338 62040
rect 54372 62006 54406 62040
rect 54440 62006 54474 62040
rect 54508 62006 54542 62040
rect 54576 62006 54610 62040
rect 54644 62006 54678 62040
rect 54712 62006 54746 62040
rect 54780 62006 54814 62040
rect 54848 62006 54882 62040
rect 54916 62006 54950 62040
rect 54984 62006 55018 62040
rect 55052 62006 55086 62040
rect 55120 62006 55154 62040
rect 55188 62006 55222 62040
rect 55256 62006 55290 62040
rect 55324 62006 55358 62040
rect 55392 62006 55426 62040
rect 55460 62006 55494 62040
rect 55528 62006 55562 62040
rect 55596 62006 55630 62040
rect 55664 62006 55698 62040
rect 55732 62006 55766 62040
rect 55800 62006 55834 62040
rect 55868 62006 55902 62040
rect 55936 62006 55970 62040
rect 56004 62006 56038 62040
rect 56072 62006 56106 62040
rect 56140 62006 56174 62040
rect 56208 62006 56242 62040
rect 56276 62006 56350 62040
rect 50456 61976 50490 62006
rect 50456 61908 50490 61942
rect 50456 61840 50490 61874
rect 50456 61772 50490 61806
rect 50456 61704 50490 61738
rect 50456 61636 50490 61670
rect 50456 61568 50490 61602
rect 50456 61500 50490 61534
rect 50456 61432 50490 61466
rect 50456 61364 50490 61398
rect 50456 61296 50490 61330
rect 50456 61228 50490 61262
rect 50456 61160 50490 61194
rect 50456 61092 50490 61126
rect 50456 61024 50490 61058
rect 50456 60956 50490 60990
rect 50456 60888 50490 60922
rect 50456 60820 50490 60854
rect 50456 60752 50490 60786
rect 50456 60684 50490 60718
rect 50456 60616 50490 60650
rect 50456 60548 50490 60582
rect 50456 60480 50490 60514
rect 50456 60412 50490 60446
rect 50456 60344 50490 60378
rect 50456 60276 50490 60310
rect 50456 60208 50490 60242
rect 50456 60140 50490 60174
rect 50456 60072 50490 60106
rect 50456 60004 50490 60038
rect 50456 59936 50490 59970
rect 50456 59868 50490 59902
rect 50456 59800 50490 59834
rect 50456 59732 50490 59766
rect 50456 59664 50490 59698
rect 50456 59596 50490 59630
rect 50456 59528 50490 59562
rect 50456 59460 50490 59494
rect 50456 59392 50490 59426
rect 50456 59324 50490 59358
rect 50456 59256 50490 59290
rect 50456 59188 50490 59222
rect 50456 59120 50490 59154
rect 50456 59052 50490 59086
rect 50456 58984 50490 59018
rect 50456 58916 50490 58950
rect 50456 58848 50490 58882
rect 50456 58780 50490 58814
rect 50456 58712 50490 58746
rect 50456 58644 50490 58678
rect 50456 58576 50490 58610
rect 50456 58508 50490 58542
rect 50456 58440 50490 58474
rect 50456 58376 50490 58406
rect 56316 61976 56350 62006
rect 56316 61908 56350 61942
rect 56316 61840 56350 61874
rect 56316 61772 56350 61806
rect 56316 61704 56350 61738
rect 56316 61636 56350 61670
rect 56316 61568 56350 61602
rect 56316 61500 56350 61534
rect 56316 61432 56350 61466
rect 56316 61364 56350 61398
rect 56316 61296 56350 61330
rect 56316 61228 56350 61262
rect 56316 61160 56350 61194
rect 56316 61092 56350 61126
rect 56316 61024 56350 61058
rect 56316 60956 56350 60990
rect 56316 60888 56350 60922
rect 56316 60820 56350 60854
rect 56316 60752 56350 60786
rect 56316 60684 56350 60718
rect 56316 60616 56350 60650
rect 56316 60548 56350 60582
rect 56316 60480 56350 60514
rect 56316 60412 56350 60446
rect 56316 60344 56350 60378
rect 56316 60276 56350 60310
rect 56316 60208 56350 60242
rect 56316 60140 56350 60174
rect 56316 60072 56350 60106
rect 56316 60004 56350 60038
rect 56316 59936 56350 59970
rect 56316 59868 56350 59902
rect 56316 59800 56350 59834
rect 56316 59732 56350 59766
rect 56316 59664 56350 59698
rect 56316 59596 56350 59630
rect 56316 59528 56350 59562
rect 56316 59460 56350 59494
rect 56316 59392 56350 59426
rect 56316 59324 56350 59358
rect 56316 59256 56350 59290
rect 56316 59188 56350 59222
rect 56316 59120 56350 59154
rect 56316 59052 56350 59086
rect 56316 58984 56350 59018
rect 56316 58916 56350 58950
rect 56316 58848 56350 58882
rect 56316 58780 56350 58814
rect 56316 58712 56350 58746
rect 56316 58644 56350 58678
rect 56316 58576 56350 58610
rect 56316 58508 56350 58542
rect 56316 58440 56350 58474
rect 56316 58376 56350 58406
rect 50456 58342 50530 58376
rect 50564 58342 50598 58376
rect 50632 58342 50666 58376
rect 50700 58342 50734 58376
rect 50768 58342 50802 58376
rect 50836 58342 50870 58376
rect 50904 58342 50938 58376
rect 50972 58342 51006 58376
rect 51040 58342 51074 58376
rect 51108 58342 51142 58376
rect 51176 58342 51210 58376
rect 51244 58342 51278 58376
rect 51312 58342 51346 58376
rect 51380 58342 51414 58376
rect 51448 58342 51482 58376
rect 51516 58342 51550 58376
rect 51584 58342 51618 58376
rect 51652 58342 51686 58376
rect 51720 58342 51754 58376
rect 51788 58342 51822 58376
rect 51856 58342 51890 58376
rect 51924 58342 51958 58376
rect 51992 58342 52026 58376
rect 52060 58342 52094 58376
rect 52128 58342 52162 58376
rect 52196 58342 52230 58376
rect 52264 58342 52298 58376
rect 52332 58342 52366 58376
rect 52400 58342 52434 58376
rect 52468 58342 52502 58376
rect 52536 58342 52570 58376
rect 52604 58342 52638 58376
rect 52672 58342 52706 58376
rect 52740 58342 52774 58376
rect 52808 58342 52842 58376
rect 52876 58342 52910 58376
rect 52944 58342 52978 58376
rect 53012 58342 53046 58376
rect 53080 58342 53114 58376
rect 53148 58342 53182 58376
rect 53216 58342 53250 58376
rect 53284 58342 53318 58376
rect 53352 58342 53386 58376
rect 53420 58342 53454 58376
rect 53488 58342 53522 58376
rect 53556 58342 53590 58376
rect 53624 58342 53658 58376
rect 53692 58342 53726 58376
rect 53760 58342 53794 58376
rect 53828 58342 53862 58376
rect 53896 58342 53930 58376
rect 53964 58342 53998 58376
rect 54032 58342 54066 58376
rect 54100 58342 54134 58376
rect 54168 58342 54202 58376
rect 54236 58342 54270 58376
rect 54304 58342 54338 58376
rect 54372 58342 54406 58376
rect 54440 58342 54474 58376
rect 54508 58342 54542 58376
rect 54576 58342 54610 58376
rect 54644 58342 54678 58376
rect 54712 58342 54746 58376
rect 54780 58342 54814 58376
rect 54848 58342 54882 58376
rect 54916 58342 54950 58376
rect 54984 58342 55018 58376
rect 55052 58342 55086 58376
rect 55120 58342 55154 58376
rect 55188 58342 55222 58376
rect 55256 58342 55290 58376
rect 55324 58342 55358 58376
rect 55392 58342 55426 58376
rect 55460 58342 55494 58376
rect 55528 58342 55562 58376
rect 55596 58342 55630 58376
rect 55664 58342 55698 58376
rect 55732 58342 55766 58376
rect 55800 58342 55834 58376
rect 55868 58342 55902 58376
rect 55936 58342 55970 58376
rect 56004 58342 56038 58376
rect 56072 58342 56106 58376
rect 56140 58342 56174 58376
rect 56208 58342 56242 58376
rect 56276 58342 56350 58376
rect 59104 62029 59138 62063
rect 59104 61961 59138 61995
rect 59104 61893 59138 61927
rect 59104 61825 59138 61859
rect 59104 61757 59138 61791
rect 59104 61689 59138 61723
rect 59104 61621 59138 61655
rect 59104 61553 59138 61587
rect 59104 61485 59138 61519
rect 59104 61417 59138 61451
rect 59104 61349 59138 61383
rect 59104 61281 59138 61315
rect 59104 61213 59138 61247
rect 59104 61145 59138 61179
rect 59104 61077 59138 61111
rect 59104 61009 59138 61043
rect 59104 60941 59138 60975
rect 59104 60873 59138 60907
rect 59104 60805 59138 60839
rect 59104 60737 59138 60771
rect 59104 60669 59138 60703
rect 59104 60601 59138 60635
rect 59104 60533 59138 60567
rect 59104 60465 59138 60499
rect 59104 60397 59138 60431
rect 59104 60329 59138 60363
rect 59104 60261 59138 60295
rect 59104 60193 59138 60227
rect 59104 60125 59138 60159
rect 59104 60057 59138 60091
rect 59104 59989 59138 60023
rect 59104 59921 59138 59955
rect 59104 59853 59138 59887
rect 59104 59785 59138 59819
rect 59104 59717 59138 59751
rect 59104 59649 59138 59683
rect 59104 59581 59138 59615
rect 59104 59513 59138 59547
rect 59104 59445 59138 59479
rect 59104 59377 59138 59411
rect 59104 59309 59138 59343
rect 59104 59241 59138 59275
rect 59104 59173 59138 59207
rect 59104 59105 59138 59139
rect 59104 59037 59138 59071
rect 59104 58969 59138 59003
rect 59104 58901 59138 58935
rect 59104 58833 59138 58867
rect 59104 58765 59138 58799
rect 59104 58697 59138 58731
rect 59104 58629 59138 58663
rect 59104 58561 59138 58595
rect 59104 58493 59138 58527
rect 59104 58425 59138 58459
rect 59104 58357 59138 58391
rect -3718 58308 -3684 58342
rect -3718 58240 -3684 58274
rect -3718 58172 -3684 58206
rect -3718 58104 -3684 58138
rect -3718 58036 -3684 58070
rect -3718 57968 -3684 58002
rect -3718 57900 -3684 57934
rect -3718 57832 -3684 57866
rect -3718 57764 -3684 57798
rect -3718 57696 -3684 57730
rect -3718 57628 -3684 57662
rect -3718 57560 -3684 57594
rect -3718 57492 -3684 57526
rect -3718 57424 -3684 57458
rect -3718 57356 -3684 57390
rect -3718 57288 -3684 57322
rect -3718 57220 -3684 57254
rect -3718 57152 -3684 57186
rect -3718 57084 -3684 57118
rect -3718 57016 -3684 57050
rect -3718 56948 -3684 56982
rect -3718 56880 -3684 56914
rect -3718 56812 -3684 56846
rect -3718 56744 -3684 56778
rect -3718 56676 -3684 56710
rect -3718 56608 -3684 56642
rect -3718 56540 -3684 56574
rect -3718 56472 -3684 56506
rect -3718 56404 -3684 56438
rect -3718 56336 -3684 56370
rect -10699 56245 -10665 56270
rect -10699 56177 -10665 56211
rect -10699 56109 -10665 56143
rect -10699 56041 -10665 56075
rect -10699 55973 -10665 56007
rect -10699 55905 -10665 55939
rect -10699 55837 -10665 55871
rect -10699 55769 -10665 55803
rect -10699 55701 -10665 55735
rect -10699 55633 -10665 55667
rect -10699 55565 -10665 55599
rect -10699 55497 -10665 55531
rect -10699 55429 -10665 55463
rect -10699 55361 -10665 55395
rect -10699 55293 -10665 55327
rect -10699 55225 -10665 55259
rect -10699 55157 -10665 55191
rect -10699 55089 -10665 55123
rect -10699 55021 -10665 55055
rect -10699 54953 -10665 54987
rect -10699 54885 -10665 54919
rect -10699 54817 -10665 54851
rect -10699 54749 -10665 54783
rect -10699 54681 -10665 54715
rect -10699 54613 -10665 54647
rect -10699 54545 -10665 54579
rect -10699 54477 -10665 54511
rect -10699 54409 -10665 54443
rect -10699 54341 -10665 54375
rect -10699 54273 -10665 54307
rect -10699 54205 -10665 54239
rect -10699 54137 -10665 54171
rect -10699 54069 -10665 54103
rect -10699 54001 -10665 54035
rect -10699 53933 -10665 53967
rect -10699 53865 -10665 53899
rect -10699 53797 -10665 53831
rect -10699 53729 -10665 53763
rect -10699 53661 -10665 53695
rect -10699 53593 -10665 53627
rect -10699 53525 -10665 53559
rect -10699 53457 -10665 53491
rect -10699 53389 -10665 53423
rect -10699 53321 -10665 53355
rect -10699 53253 -10665 53287
rect -10699 53185 -10665 53219
rect -10699 53117 -10665 53151
rect -10699 53049 -10665 53083
rect -10699 52981 -10665 53015
rect -10699 52913 -10665 52947
rect -10699 52845 -10665 52879
rect -10699 52777 -10665 52811
rect -10699 52709 -10665 52743
rect -10699 52641 -10665 52675
rect -10699 52573 -10665 52607
rect -10699 52505 -10665 52539
rect -10699 52437 -10665 52471
rect -10699 52369 -10665 52403
rect -10699 52301 -10665 52335
rect -10699 52233 -10665 52267
rect -10699 52165 -10665 52199
rect -10699 52097 -10665 52131
rect -10699 52029 -10665 52063
rect -10699 51961 -10665 51995
rect -10699 51893 -10665 51927
rect -10699 51825 -10665 51859
rect -10699 51757 -10665 51791
rect -10699 51689 -10665 51723
rect -10699 51621 -10665 51655
rect -10699 51553 -10665 51587
rect -10699 51485 -10665 51519
rect -10699 51417 -10665 51451
rect -10699 51349 -10665 51383
rect -10699 51281 -10665 51315
rect -10699 51213 -10665 51247
rect -10699 51145 -10665 51179
rect -10699 51077 -10665 51111
rect -10699 51009 -10665 51043
rect -10699 50941 -10665 50975
rect -10699 50873 -10665 50907
rect -10699 50805 -10665 50839
rect -10699 50737 -10665 50771
rect -10699 50669 -10665 50703
rect -10699 50601 -10665 50635
rect -10699 50533 -10665 50567
rect -10699 50465 -10665 50499
rect -10699 50397 -10665 50431
rect -10699 50329 -10665 50363
rect -10699 50261 -10665 50295
rect -10699 50193 -10665 50227
rect -10699 50125 -10665 50159
rect -10699 50057 -10665 50091
rect -10699 49989 -10665 50023
rect -10699 49921 -10665 49955
rect -10699 49853 -10665 49887
rect -10699 49785 -10665 49819
rect -10699 49717 -10665 49751
rect -10699 49649 -10665 49683
rect -10699 49581 -10665 49615
rect -10699 49513 -10665 49547
rect -10699 49445 -10665 49479
rect -10699 49377 -10665 49411
rect -10699 49309 -10665 49343
rect -10699 49241 -10665 49275
rect -10699 49173 -10665 49207
rect -10699 49105 -10665 49139
rect -10699 49037 -10665 49071
rect -10699 48969 -10665 49003
rect -10699 48901 -10665 48935
rect -10699 48833 -10665 48867
rect -10699 48765 -10665 48799
rect -10699 48697 -10665 48731
rect -10699 48629 -10665 48663
rect -10699 48561 -10665 48595
rect -10699 48493 -10665 48527
rect -10699 48425 -10665 48459
rect -10699 48357 -10665 48391
rect -10699 48289 -10665 48323
rect -10699 48221 -10665 48255
rect -10699 48153 -10665 48187
rect -10699 48085 -10665 48119
rect -10699 48017 -10665 48051
rect -10699 47949 -10665 47983
rect -10699 47881 -10665 47915
rect -10699 47813 -10665 47847
rect -10699 47745 -10665 47779
rect -10699 47677 -10665 47711
rect -10699 47609 -10665 47643
rect -10699 47541 -10665 47575
rect -10699 47473 -10665 47507
rect -10699 47405 -10665 47439
rect -10699 47337 -10665 47371
rect -10699 47269 -10665 47303
rect -10699 47201 -10665 47235
rect -10699 47133 -10665 47167
rect -10699 47065 -10665 47099
rect -10699 46997 -10665 47031
rect -10699 46929 -10665 46963
rect -10699 46861 -10665 46895
rect -10699 46793 -10665 46827
rect -10699 46725 -10665 46759
rect -10699 46657 -10665 46691
rect -10699 46589 -10665 46623
rect -10699 46521 -10665 46555
rect -10699 46453 -10665 46487
rect -10699 46385 -10665 46419
rect -10699 46317 -10665 46351
rect -10699 46249 -10665 46283
rect -10699 46181 -10665 46215
rect -10699 46113 -10665 46147
rect -10699 46045 -10665 46079
rect -10699 45977 -10665 46011
rect -10699 45909 -10665 45943
rect -10699 45841 -10665 45875
rect -10699 45773 -10665 45807
rect -10699 45705 -10665 45739
rect -10699 45637 -10665 45671
rect -10699 45569 -10665 45603
rect -10699 45501 -10665 45535
rect -10699 45433 -10665 45467
rect -10699 45365 -10665 45399
rect -10699 45297 -10665 45331
rect -10699 45229 -10665 45263
rect -10699 45161 -10665 45195
rect -10699 45093 -10665 45127
rect -10699 45025 -10665 45059
rect -10699 44957 -10665 44991
rect -10699 44889 -10665 44923
rect -10699 44821 -10665 44855
rect -10699 44753 -10665 44787
rect -10699 44685 -10665 44719
rect -10699 44617 -10665 44651
rect -10699 44549 -10665 44583
rect -10699 44481 -10665 44515
rect -10699 44413 -10665 44447
rect -10699 44345 -10665 44379
rect -10699 44280 -10665 44311
rect -3718 56268 -3684 56302
rect -3718 56200 -3684 56234
rect -3718 56132 -3684 56166
rect -3718 56064 -3684 56098
rect -3718 55996 -3684 56030
rect -3718 55928 -3684 55962
rect -3718 55860 -3684 55894
rect -3718 55792 -3684 55826
rect -3718 55724 -3684 55758
rect -3718 55656 -3684 55690
rect -3718 55588 -3684 55622
rect -3718 55520 -3684 55554
rect -3718 55452 -3684 55486
rect -3718 55384 -3684 55418
rect -3718 55316 -3684 55350
rect -3718 55248 -3684 55282
rect -3718 55180 -3684 55214
rect -3718 55112 -3684 55146
rect -3718 55044 -3684 55078
rect -3718 54976 -3684 55010
rect -3718 54908 -3684 54942
rect -3718 54840 -3684 54874
rect -3718 54772 -3684 54806
rect -3718 54704 -3684 54738
rect -3718 54636 -3684 54670
rect -3718 54568 -3684 54602
rect -3718 54500 -3684 54534
rect -3718 54432 -3684 54466
rect -3718 54364 -3684 54398
rect -3718 54296 -3684 54330
rect -3718 54228 -3684 54262
rect -3718 54160 -3684 54194
rect -3718 54092 -3684 54126
rect -3718 54024 -3684 54058
rect -3718 53956 -3684 53990
rect -3718 53888 -3684 53922
rect -3718 53820 -3684 53854
rect -3718 53752 -3684 53786
rect -3718 53684 -3684 53718
rect -3718 53616 -3684 53650
rect -3718 53548 -3684 53582
rect -3718 53480 -3684 53514
rect -3718 53412 -3684 53446
rect -3718 53344 -3684 53378
rect -3718 53276 -3684 53310
rect -3718 53208 -3684 53242
rect -3718 53140 -3684 53174
rect -3718 53072 -3684 53106
rect -3718 53004 -3684 53038
rect -3718 52936 -3684 52970
rect -3718 52868 -3684 52902
rect -3718 52800 -3684 52834
rect -3718 52732 -3684 52766
rect -3718 52664 -3684 52698
rect -3718 52596 -3684 52630
rect -3718 52528 -3684 52562
rect -3718 52460 -3684 52494
rect -3718 52392 -3684 52426
rect -3718 52324 -3684 52358
rect -3718 52256 -3684 52290
rect -3718 52188 -3684 52222
rect -3718 52120 -3684 52154
rect -3718 52052 -3684 52086
rect -3718 51984 -3684 52018
rect -3718 51916 -3684 51950
rect -3718 51848 -3684 51882
rect -3718 51780 -3684 51814
rect -3718 51712 -3684 51746
rect -3718 51644 -3684 51678
rect -3718 51576 -3684 51610
rect -3718 51508 -3684 51542
rect -3718 51440 -3684 51474
rect -3718 51372 -3684 51406
rect -3718 51304 -3684 51338
rect -3718 51236 -3684 51270
rect -3718 51168 -3684 51202
rect -3718 51100 -3684 51134
rect -3718 51032 -3684 51066
rect -3718 50964 -3684 50998
rect -3718 50896 -3684 50930
rect -3718 50828 -3684 50862
rect -3718 50760 -3684 50794
rect -3718 50692 -3684 50726
rect -3718 50624 -3684 50658
rect -3718 50556 -3684 50590
rect -3718 50488 -3684 50522
rect -3718 50420 -3684 50454
rect -3718 50352 -3684 50386
rect -3718 50284 -3684 50318
rect -3718 50216 -3684 50250
rect -3718 50148 -3684 50182
rect -3718 50080 -3684 50114
rect -3718 50012 -3684 50046
rect -3718 49944 -3684 49978
rect -3718 49876 -3684 49910
rect -3718 49808 -3684 49842
rect -3718 49740 -3684 49774
rect -3718 49672 -3684 49706
rect -3718 49604 -3684 49638
rect -3718 49536 -3684 49570
rect -3718 49468 -3684 49502
rect -3718 49400 -3684 49434
rect -3718 49332 -3684 49366
rect -3718 49264 -3684 49298
rect -3718 49196 -3684 49230
rect -3718 49128 -3684 49162
rect -3718 49060 -3684 49094
rect -3718 48992 -3684 49026
rect -3718 48924 -3684 48958
rect -3718 48856 -3684 48890
rect -3718 48788 -3684 48822
rect -3718 48720 -3684 48754
rect -3718 48652 -3684 48686
rect -3718 48584 -3684 48618
rect -3718 48516 -3684 48550
rect -3718 48448 -3684 48482
rect -3718 48380 -3684 48414
rect -3718 48312 -3684 48346
rect -3718 48244 -3684 48278
rect -3718 48176 -3684 48210
rect -3718 48108 -3684 48142
rect -3718 48040 -3684 48074
rect -3718 47972 -3684 48006
rect -3718 47904 -3684 47938
rect -3718 47836 -3684 47870
rect -3718 47768 -3684 47802
rect -3718 47700 -3684 47734
rect -3718 47632 -3684 47666
rect -3718 47564 -3684 47598
rect -3718 47496 -3684 47530
rect -3718 47428 -3684 47462
rect -3718 47360 -3684 47394
rect -3718 47292 -3684 47326
rect -3718 47224 -3684 47258
rect -3718 47156 -3684 47190
rect -3718 47088 -3684 47122
rect -3718 47020 -3684 47054
rect -3718 46952 -3684 46986
rect -3718 46884 -3684 46918
rect -3718 46816 -3684 46850
rect -3718 46748 -3684 46782
rect -3718 46680 -3684 46714
rect -3718 46612 -3684 46646
rect -3718 46544 -3684 46578
rect -3718 46476 -3684 46510
rect -3718 46408 -3684 46442
rect -3718 46340 -3684 46374
rect -3718 46272 -3684 46306
rect -3718 46204 -3684 46238
rect -3718 46136 -3684 46170
rect -3718 46068 -3684 46102
rect -3718 46000 -3684 46034
rect -3718 45932 -3684 45966
rect -3718 45864 -3684 45898
rect 59104 58289 59138 58323
rect 59104 58221 59138 58255
rect 59104 58153 59138 58187
rect 59104 58085 59138 58119
rect 59104 58017 59138 58051
rect 59104 57949 59138 57983
rect 59104 57881 59138 57915
rect 59104 57813 59138 57847
rect 59104 57745 59138 57779
rect 59104 57677 59138 57711
rect 59104 57609 59138 57643
rect 59104 57541 59138 57575
rect 59104 57473 59138 57507
rect 59104 57405 59138 57439
rect 59104 57337 59138 57371
rect 59104 57269 59138 57303
rect 59104 57201 59138 57235
rect 59104 57133 59138 57167
rect 59104 57065 59138 57099
rect 59104 56997 59138 57031
rect 59104 56929 59138 56963
rect 59104 56861 59138 56895
rect 59104 56793 59138 56827
rect 59104 56725 59138 56759
rect 59104 56657 59138 56691
rect 59104 56589 59138 56623
rect 59104 56521 59138 56555
rect 59104 56453 59138 56487
rect 59104 56385 59138 56419
rect 59104 56317 59138 56351
rect 59104 56249 59138 56283
rect 59104 56181 59138 56215
rect 59104 56113 59138 56147
rect 59104 56045 59138 56079
rect 59104 55977 59138 56011
rect 59104 55909 59138 55943
rect 59104 55841 59138 55875
rect 59104 55773 59138 55807
rect 59104 55705 59138 55739
rect 59104 55637 59138 55671
rect 59104 55569 59138 55603
rect 59104 55501 59138 55535
rect 59104 55433 59138 55467
rect 59104 55365 59138 55399
rect 59104 55297 59138 55331
rect 59104 55229 59138 55263
rect 59104 55161 59138 55195
rect 59104 55093 59138 55127
rect 59104 55025 59138 55059
rect 59104 54957 59138 54991
rect 59104 54889 59138 54923
rect 59104 54821 59138 54855
rect 59104 54753 59138 54787
rect 59104 54685 59138 54719
rect 59104 54617 59138 54651
rect 59104 54549 59138 54583
rect 59104 54481 59138 54515
rect 59104 54413 59138 54447
rect 59104 54345 59138 54379
rect 59104 54277 59138 54311
rect 59104 54209 59138 54243
rect 59104 54141 59138 54175
rect 59104 54073 59138 54107
rect 59104 54005 59138 54039
rect 59104 53937 59138 53971
rect 59104 53869 59138 53903
rect 59104 53801 59138 53835
rect 59104 53733 59138 53767
rect 59104 53665 59138 53699
rect 59104 53597 59138 53631
rect 59104 53529 59138 53563
rect 59104 53461 59138 53495
rect 59104 53393 59138 53427
rect 59104 53325 59138 53359
rect 59104 53257 59138 53291
rect 59104 53189 59138 53223
rect 59104 53121 59138 53155
rect 59104 53053 59138 53087
rect 59104 52985 59138 53019
rect 59104 52917 59138 52951
rect 59104 52849 59138 52883
rect 59104 52781 59138 52815
rect 59104 52713 59138 52747
rect 59104 52645 59138 52679
rect 59104 52577 59138 52611
rect 59104 52509 59138 52543
rect 59104 52441 59138 52475
rect 59104 52373 59138 52407
rect 59104 52305 59138 52339
rect 59104 52237 59138 52271
rect 59104 52169 59138 52203
rect 59104 52101 59138 52135
rect 59104 52033 59138 52067
rect 59104 51965 59138 51999
rect 59104 51897 59138 51931
rect 59104 51829 59138 51863
rect 59104 51761 59138 51795
rect 59104 51693 59138 51727
rect 59104 51625 59138 51659
rect 59104 51557 59138 51591
rect 59104 51489 59138 51523
rect 59104 51421 59138 51455
rect 59104 51353 59138 51387
rect 59104 51285 59138 51319
rect 59104 51217 59138 51251
rect 59104 51149 59138 51183
rect 59104 51081 59138 51115
rect 59104 51013 59138 51047
rect 59104 50945 59138 50979
rect 59104 50877 59138 50911
rect 59104 50809 59138 50843
rect 59104 50741 59138 50775
rect 59104 50673 59138 50707
rect 59104 50605 59138 50639
rect 59104 50537 59138 50571
rect 59104 50469 59138 50503
rect 59104 50401 59138 50435
rect 59104 50333 59138 50367
rect 59104 50265 59138 50299
rect 59104 50197 59138 50231
rect 59104 50129 59138 50163
rect 59104 50061 59138 50095
rect 59104 49993 59138 50027
rect 59104 49925 59138 49959
rect 59104 49857 59138 49891
rect 59104 49789 59138 49823
rect 59104 49721 59138 49755
rect 59104 49653 59138 49687
rect 59104 49585 59138 49619
rect 59104 49517 59138 49551
rect 59104 49449 59138 49483
rect 59104 49381 59138 49415
rect 59104 49313 59138 49347
rect 59104 49245 59138 49279
rect 59104 49177 59138 49211
rect 59104 49109 59138 49143
rect 59104 49041 59138 49075
rect 59104 48973 59138 49007
rect 59104 48905 59138 48939
rect 59104 48837 59138 48871
rect 59104 48769 59138 48803
rect 59104 48701 59138 48735
rect 59104 48633 59138 48667
rect 59104 48565 59138 48599
rect 59104 48497 59138 48531
rect 59104 48429 59138 48463
rect 59104 48361 59138 48395
rect 59104 48293 59138 48327
rect 59104 48225 59138 48259
rect 59104 48157 59138 48191
rect 59104 48089 59138 48123
rect 59104 48021 59138 48055
rect 59104 47953 59138 47987
rect 59104 47885 59138 47919
rect 59104 47817 59138 47851
rect 59104 47749 59138 47783
rect 59104 47681 59138 47715
rect 59104 47613 59138 47647
rect 59104 47545 59138 47579
rect 59104 47477 59138 47511
rect 59104 47409 59138 47443
rect 59104 47341 59138 47375
rect 59104 47273 59138 47307
rect 59104 47205 59138 47239
rect 59104 47137 59138 47171
rect 59104 47069 59138 47103
rect 59104 47001 59138 47035
rect 59104 46933 59138 46967
rect 59104 46865 59138 46899
rect 59104 46797 59138 46831
rect 59104 46729 59138 46763
rect 59104 46661 59138 46695
rect 59104 46593 59138 46627
rect 59104 46525 59138 46559
rect 59104 46457 59138 46491
rect 59104 46389 59138 46423
rect 59104 46321 59138 46355
rect 59104 46253 59138 46287
rect 59104 46185 59138 46219
rect 59104 46117 59138 46151
rect 59104 46049 59138 46083
rect 59104 45981 59138 46015
rect 59104 45920 59138 45947
rect 70838 74745 70872 74772
rect 70838 74677 70872 74711
rect 70838 74609 70872 74643
rect 70838 74541 70872 74575
rect 70838 74473 70872 74507
rect 70838 74405 70872 74439
rect 70838 74337 70872 74371
rect 70838 74269 70872 74303
rect 70838 74201 70872 74235
rect 70838 74133 70872 74167
rect 70838 74065 70872 74099
rect 70838 73997 70872 74031
rect 70838 73929 70872 73963
rect 70838 73861 70872 73895
rect 70838 73793 70872 73827
rect 70838 73725 70872 73759
rect 70838 73657 70872 73691
rect 70838 73589 70872 73623
rect 70838 73521 70872 73555
rect 70838 73453 70872 73487
rect 70838 73385 70872 73419
rect 70838 73317 70872 73351
rect 70838 73249 70872 73283
rect 70838 73181 70872 73215
rect 70838 73113 70872 73147
rect 70838 73045 70872 73079
rect 70838 72977 70872 73011
rect 70838 72909 70872 72943
rect 70838 72841 70872 72875
rect 70838 72773 70872 72807
rect 70838 72705 70872 72739
rect 70838 72637 70872 72671
rect 70838 72569 70872 72603
rect 70838 72501 70872 72535
rect 70838 72433 70872 72467
rect 70838 72365 70872 72399
rect 70838 72297 70872 72331
rect 70838 72229 70872 72263
rect 70838 72161 70872 72195
rect 70838 72093 70872 72127
rect 70838 72025 70872 72059
rect 70838 71957 70872 71991
rect 70838 71889 70872 71923
rect 70838 71821 70872 71855
rect 70838 71753 70872 71787
rect 70838 71685 70872 71719
rect 70838 71617 70872 71651
rect 70838 71549 70872 71583
rect 70838 71481 70872 71515
rect 70838 71413 70872 71447
rect 70838 71345 70872 71379
rect 70838 71277 70872 71311
rect 70838 71209 70872 71243
rect 70838 71141 70872 71175
rect 70838 71073 70872 71107
rect 70838 71005 70872 71039
rect 70838 70937 70872 70971
rect 70838 70869 70872 70903
rect 70838 70801 70872 70835
rect 70838 70733 70872 70767
rect 70838 70665 70872 70699
rect 70838 70597 70872 70631
rect 70838 70529 70872 70563
rect 70838 70461 70872 70495
rect 70838 70393 70872 70427
rect 70838 70325 70872 70359
rect 70838 70257 70872 70291
rect 70838 70189 70872 70223
rect 70838 70121 70872 70155
rect 70838 70053 70872 70087
rect 70838 69985 70872 70019
rect 70838 69917 70872 69951
rect 70838 69849 70872 69883
rect 70838 69781 70872 69815
rect 70838 69713 70872 69747
rect 70838 69645 70872 69679
rect 70838 69577 70872 69611
rect 70838 69509 70872 69543
rect 70838 69441 70872 69475
rect 70838 69373 70872 69407
rect 70838 69305 70872 69339
rect 70838 69237 70872 69271
rect 70838 69169 70872 69203
rect 70838 69101 70872 69135
rect 70838 69033 70872 69067
rect 70838 68965 70872 68999
rect 70838 68897 70872 68931
rect 70838 68829 70872 68863
rect 70838 68761 70872 68795
rect 70838 68693 70872 68727
rect 70838 68625 70872 68659
rect 70838 68557 70872 68591
rect 70838 68489 70872 68523
rect 70838 68421 70872 68455
rect 70838 68353 70872 68387
rect 70838 68285 70872 68319
rect 70838 68217 70872 68251
rect 70838 68149 70872 68183
rect 70838 68081 70872 68115
rect 70838 68013 70872 68047
rect 70838 67945 70872 67979
rect 70838 67877 70872 67911
rect 70838 67809 70872 67843
rect 70838 67741 70872 67775
rect 70838 67673 70872 67707
rect 70838 67605 70872 67639
rect 70838 67537 70872 67571
rect 70838 67469 70872 67503
rect 70838 67401 70872 67435
rect 70838 67333 70872 67367
rect 70838 67265 70872 67299
rect 70838 67197 70872 67231
rect 70838 67129 70872 67163
rect 70838 67061 70872 67095
rect 70838 66993 70872 67027
rect 70838 66925 70872 66959
rect 70838 66857 70872 66891
rect 70838 66789 70872 66823
rect 70838 66721 70872 66755
rect 70838 66653 70872 66687
rect 70838 66585 70872 66619
rect 70838 66517 70872 66551
rect 70838 66449 70872 66483
rect 70838 66381 70872 66415
rect 70838 66313 70872 66347
rect 70838 66245 70872 66279
rect 70838 66177 70872 66211
rect 70838 66109 70872 66143
rect 70838 66041 70872 66075
rect 70838 65973 70872 66007
rect 70838 65905 70872 65939
rect 70838 65837 70872 65871
rect 70838 65769 70872 65803
rect 70838 65701 70872 65735
rect 70838 65633 70872 65667
rect 70838 65565 70872 65599
rect 70838 65497 70872 65531
rect 70838 65429 70872 65463
rect 70838 65361 70872 65395
rect 70838 65293 70872 65327
rect 70838 65225 70872 65259
rect 70838 65157 70872 65191
rect 70838 65089 70872 65123
rect 70838 65021 70872 65055
rect 70838 64953 70872 64987
rect 70838 64885 70872 64919
rect 70838 64817 70872 64851
rect 70838 64749 70872 64783
rect 70838 64681 70872 64715
rect 70838 64613 70872 64647
rect 70838 64545 70872 64579
rect 70838 64477 70872 64511
rect 70838 64409 70872 64443
rect 70838 64341 70872 64375
rect 70838 64273 70872 64307
rect 70838 64205 70872 64239
rect 70838 64137 70872 64171
rect 70838 64069 70872 64103
rect 70838 64001 70872 64035
rect 70838 63933 70872 63967
rect 70838 63865 70872 63899
rect 70838 63797 70872 63831
rect 70838 63729 70872 63763
rect 70838 63661 70872 63695
rect 70838 63593 70872 63627
rect 70838 63525 70872 63559
rect 70838 63457 70872 63491
rect 70838 63389 70872 63423
rect 70838 63321 70872 63355
rect 70838 63253 70872 63287
rect 70838 63185 70872 63219
rect 70838 63117 70872 63151
rect 70838 63049 70872 63083
rect 70838 62981 70872 63015
rect 70838 62913 70872 62947
rect 70838 62845 70872 62879
rect 70838 62777 70872 62811
rect 70838 62709 70872 62743
rect 70838 62641 70872 62675
rect 70838 62573 70872 62607
rect 70838 62505 70872 62539
rect 70838 62437 70872 62471
rect 70838 62369 70872 62403
rect 70838 62301 70872 62335
rect 70838 62233 70872 62267
rect 70838 62165 70872 62199
rect 70838 62097 70872 62131
rect 70838 62029 70872 62063
rect 70838 61961 70872 61995
rect 70838 61893 70872 61927
rect 70838 61825 70872 61859
rect 70838 61757 70872 61791
rect 70838 61689 70872 61723
rect 70838 61621 70872 61655
rect 70838 61553 70872 61587
rect 70838 61485 70872 61519
rect 70838 61417 70872 61451
rect 70838 61349 70872 61383
rect 70838 61281 70872 61315
rect 70838 61213 70872 61247
rect 70838 61145 70872 61179
rect 70838 61077 70872 61111
rect 70838 61009 70872 61043
rect 70838 60941 70872 60975
rect 70838 60873 70872 60907
rect 70838 60805 70872 60839
rect 70838 60737 70872 60771
rect 70838 60669 70872 60703
rect 70838 60601 70872 60635
rect 70838 60533 70872 60567
rect 70838 60465 70872 60499
rect 70838 60397 70872 60431
rect 70838 60329 70872 60363
rect 70838 60261 70872 60295
rect 70838 60193 70872 60227
rect 70838 60125 70872 60159
rect 70838 60057 70872 60091
rect 70838 59989 70872 60023
rect 70838 59921 70872 59955
rect 70838 59853 70872 59887
rect 70838 59785 70872 59819
rect 70838 59717 70872 59751
rect 70838 59649 70872 59683
rect 70838 59581 70872 59615
rect 70838 59513 70872 59547
rect 70838 59445 70872 59479
rect 70838 59377 70872 59411
rect 70838 59309 70872 59343
rect 70838 59241 70872 59275
rect 70838 59173 70872 59207
rect 70838 59105 70872 59139
rect 70838 59037 70872 59071
rect 70838 58969 70872 59003
rect 70838 58901 70872 58935
rect 70838 58833 70872 58867
rect 70838 58765 70872 58799
rect 70838 58697 70872 58731
rect 70838 58629 70872 58663
rect 70838 58561 70872 58595
rect 70838 58493 70872 58527
rect 70838 58425 70872 58459
rect 70838 58357 70872 58391
rect 70838 58289 70872 58323
rect 70838 58221 70872 58255
rect 70838 58153 70872 58187
rect 70838 58085 70872 58119
rect 70838 58017 70872 58051
rect 70838 57949 70872 57983
rect 70838 57881 70872 57915
rect 70838 57813 70872 57847
rect 70838 57745 70872 57779
rect 70838 57677 70872 57711
rect 70838 57609 70872 57643
rect 70838 57541 70872 57575
rect 70838 57473 70872 57507
rect 70838 57405 70872 57439
rect 70838 57337 70872 57371
rect 70838 57269 70872 57303
rect 70838 57201 70872 57235
rect 70838 57133 70872 57167
rect 70838 57065 70872 57099
rect 70838 56997 70872 57031
rect 70838 56929 70872 56963
rect 70838 56861 70872 56895
rect 70838 56793 70872 56827
rect 70838 56725 70872 56759
rect 70838 56657 70872 56691
rect 70838 56589 70872 56623
rect 70838 56521 70872 56555
rect 70838 56453 70872 56487
rect 70838 56385 70872 56419
rect 70838 56317 70872 56351
rect 70838 56249 70872 56283
rect 70838 56181 70872 56215
rect 70838 56113 70872 56147
rect 70838 56045 70872 56079
rect 70838 55977 70872 56011
rect 70838 55909 70872 55943
rect 70838 55841 70872 55875
rect 70838 55773 70872 55807
rect 70838 55705 70872 55739
rect 70838 55637 70872 55671
rect 70838 55569 70872 55603
rect 70838 55501 70872 55535
rect 70838 55433 70872 55467
rect 70838 55365 70872 55399
rect 70838 55297 70872 55331
rect 70838 55229 70872 55263
rect 70838 55161 70872 55195
rect 70838 55093 70872 55127
rect 70838 55025 70872 55059
rect 70838 54957 70872 54991
rect 70838 54889 70872 54923
rect 70838 54821 70872 54855
rect 70838 54753 70872 54787
rect 70838 54685 70872 54719
rect 70838 54617 70872 54651
rect 70838 54549 70872 54583
rect 70838 54481 70872 54515
rect 70838 54413 70872 54447
rect 70838 54345 70872 54379
rect 70838 54277 70872 54311
rect 70838 54209 70872 54243
rect 70838 54141 70872 54175
rect 70838 54073 70872 54107
rect 70838 54005 70872 54039
rect 70838 53937 70872 53971
rect 70838 53869 70872 53903
rect 70838 53801 70872 53835
rect 70838 53733 70872 53767
rect 70838 53665 70872 53699
rect 70838 53597 70872 53631
rect 70838 53529 70872 53563
rect 70838 53461 70872 53495
rect 70838 53393 70872 53427
rect 70838 53325 70872 53359
rect 70838 53257 70872 53291
rect 70838 53189 70872 53223
rect 70838 53121 70872 53155
rect 70838 53053 70872 53087
rect 70838 52985 70872 53019
rect 70838 52917 70872 52951
rect 70838 52849 70872 52883
rect 70838 52781 70872 52815
rect 70838 52713 70872 52747
rect 70838 52645 70872 52679
rect 70838 52577 70872 52611
rect 70838 52509 70872 52543
rect 70838 52441 70872 52475
rect 70838 52373 70872 52407
rect 70838 52305 70872 52339
rect 70838 52237 70872 52271
rect 70838 52169 70872 52203
rect 70838 52101 70872 52135
rect 70838 52033 70872 52067
rect 70838 51965 70872 51999
rect 70838 51897 70872 51931
rect 70838 51829 70872 51863
rect 70838 51761 70872 51795
rect 70838 51693 70872 51727
rect 70838 51625 70872 51659
rect 70838 51557 70872 51591
rect 70838 51489 70872 51523
rect 70838 51421 70872 51455
rect 70838 51353 70872 51387
rect 70838 51285 70872 51319
rect 70838 51217 70872 51251
rect 70838 51149 70872 51183
rect 70838 51081 70872 51115
rect 70838 51013 70872 51047
rect 70838 50945 70872 50979
rect 70838 50877 70872 50911
rect 70838 50809 70872 50843
rect 70838 50741 70872 50775
rect 70838 50673 70872 50707
rect 70838 50605 70872 50639
rect 70838 50537 70872 50571
rect 70838 50469 70872 50503
rect 70838 50401 70872 50435
rect 70838 50333 70872 50367
rect 70838 50265 70872 50299
rect 70838 50197 70872 50231
rect 70838 50129 70872 50163
rect 70838 50061 70872 50095
rect 70838 49993 70872 50027
rect 70838 49925 70872 49959
rect 70838 49857 70872 49891
rect 70838 49789 70872 49823
rect 70838 49721 70872 49755
rect 70838 49653 70872 49687
rect 70838 49585 70872 49619
rect 70838 49517 70872 49551
rect 70838 49449 70872 49483
rect 70838 49381 70872 49415
rect 70838 49313 70872 49347
rect 70838 49245 70872 49279
rect 70838 49177 70872 49211
rect 70838 49109 70872 49143
rect 70838 49041 70872 49075
rect 70838 48973 70872 49007
rect 70838 48905 70872 48939
rect 70838 48837 70872 48871
rect 70838 48769 70872 48803
rect 70838 48701 70872 48735
rect 70838 48633 70872 48667
rect 70838 48565 70872 48599
rect 70838 48497 70872 48531
rect 70838 48429 70872 48463
rect 70838 48361 70872 48395
rect 70838 48293 70872 48327
rect 70838 48225 70872 48259
rect 70838 48157 70872 48191
rect 70838 48089 70872 48123
rect 70838 48021 70872 48055
rect 70838 47953 70872 47987
rect 70838 47885 70872 47919
rect 70838 47817 70872 47851
rect 70838 47749 70872 47783
rect 70838 47681 70872 47715
rect 70838 47613 70872 47647
rect 70838 47545 70872 47579
rect 70838 47477 70872 47511
rect 70838 47409 70872 47443
rect 70838 47341 70872 47375
rect 70838 47273 70872 47307
rect 70838 47205 70872 47239
rect 70838 47137 70872 47171
rect 70838 47069 70872 47103
rect 70838 47001 70872 47035
rect 70838 46933 70872 46967
rect 70838 46865 70872 46899
rect 70838 46797 70872 46831
rect 70838 46729 70872 46763
rect 70838 46661 70872 46695
rect 70838 46593 70872 46627
rect 70838 46525 70872 46559
rect 70838 46457 70872 46491
rect 70838 46389 70872 46423
rect 70838 46321 70872 46355
rect 70838 46253 70872 46287
rect 70838 46185 70872 46219
rect 70838 46117 70872 46151
rect 70838 46049 70872 46083
rect 70838 45981 70872 46015
rect 70838 45920 70872 45947
rect 59104 45886 59191 45920
rect 59225 45886 59259 45920
rect 59293 45886 59327 45920
rect 59361 45886 59395 45920
rect 59429 45886 59463 45920
rect 59497 45886 59531 45920
rect 59565 45886 59599 45920
rect 59633 45886 59667 45920
rect 59701 45886 59735 45920
rect 59769 45886 59803 45920
rect 59837 45886 59871 45920
rect 59905 45886 59939 45920
rect 59973 45886 60007 45920
rect 60041 45886 60075 45920
rect 60109 45886 60143 45920
rect 60177 45886 60211 45920
rect 60245 45886 60279 45920
rect 60313 45886 60347 45920
rect 60381 45886 60415 45920
rect 60449 45886 60483 45920
rect 60517 45886 60551 45920
rect 60585 45886 60619 45920
rect 60653 45886 60687 45920
rect 60721 45886 60755 45920
rect 60789 45886 60823 45920
rect 60857 45886 60891 45920
rect 60925 45886 60959 45920
rect 60993 45886 61027 45920
rect 61061 45886 61095 45920
rect 61129 45886 61163 45920
rect 61197 45886 61231 45920
rect 61265 45886 61299 45920
rect 61333 45886 61367 45920
rect 61401 45886 61435 45920
rect 61469 45886 61503 45920
rect 61537 45886 61571 45920
rect 61605 45886 61639 45920
rect 61673 45886 61707 45920
rect 61741 45886 61775 45920
rect 61809 45886 61843 45920
rect 61877 45886 61911 45920
rect 61945 45886 61979 45920
rect 62013 45886 62047 45920
rect 62081 45886 62115 45920
rect 62149 45886 62183 45920
rect 62217 45886 62251 45920
rect 62285 45886 62319 45920
rect 62353 45886 62387 45920
rect 62421 45886 62455 45920
rect 62489 45886 62523 45920
rect 62557 45886 62591 45920
rect 62625 45886 62659 45920
rect 62693 45886 62727 45920
rect 62761 45886 62795 45920
rect 62829 45886 62863 45920
rect 62897 45886 62931 45920
rect 62965 45886 62999 45920
rect 63033 45886 63067 45920
rect 63101 45886 63135 45920
rect 63169 45886 63203 45920
rect 63237 45886 63271 45920
rect 63305 45886 63339 45920
rect 63373 45886 63407 45920
rect 63441 45886 63475 45920
rect 63509 45886 63543 45920
rect 63577 45886 63611 45920
rect 63645 45886 63679 45920
rect 63713 45886 63747 45920
rect 63781 45886 63815 45920
rect 63849 45886 63883 45920
rect 63917 45886 63951 45920
rect 63985 45886 64019 45920
rect 64053 45886 64087 45920
rect 64121 45886 64155 45920
rect 64189 45886 64223 45920
rect 64257 45886 64291 45920
rect 64325 45886 64359 45920
rect 64393 45886 64427 45920
rect 64461 45886 64495 45920
rect 64529 45886 64563 45920
rect 64597 45886 64631 45920
rect 64665 45886 64699 45920
rect 64733 45886 64767 45920
rect 64801 45886 64835 45920
rect 64869 45886 64903 45920
rect 64937 45886 64971 45920
rect 65005 45886 65039 45920
rect 65073 45886 65107 45920
rect 65141 45886 65175 45920
rect 65209 45886 65243 45920
rect 65277 45886 65311 45920
rect 65345 45886 65379 45920
rect 65413 45886 65447 45920
rect 65481 45886 65515 45920
rect 65549 45886 65583 45920
rect 65617 45886 65651 45920
rect 65685 45886 65719 45920
rect 65753 45886 65787 45920
rect 65821 45886 65855 45920
rect 65889 45886 65923 45920
rect 65957 45886 65991 45920
rect 66025 45886 66059 45920
rect 66093 45886 66127 45920
rect 66161 45886 66195 45920
rect 66229 45886 66263 45920
rect 66297 45886 66331 45920
rect 66365 45886 66399 45920
rect 66433 45886 66467 45920
rect 66501 45886 66535 45920
rect 66569 45886 66603 45920
rect 66637 45886 66671 45920
rect 66705 45886 66739 45920
rect 66773 45886 66807 45920
rect 66841 45886 66875 45920
rect 66909 45886 66943 45920
rect 66977 45886 67011 45920
rect 67045 45886 67079 45920
rect 67113 45886 67147 45920
rect 67181 45886 67215 45920
rect 67249 45886 67283 45920
rect 67317 45886 67351 45920
rect 67385 45886 67419 45920
rect 67453 45886 67487 45920
rect 67521 45886 67555 45920
rect 67589 45886 67623 45920
rect 67657 45886 67691 45920
rect 67725 45886 67759 45920
rect 67793 45886 67827 45920
rect 67861 45886 67895 45920
rect 67929 45886 67963 45920
rect 67997 45886 68031 45920
rect 68065 45886 68099 45920
rect 68133 45886 68167 45920
rect 68201 45886 68235 45920
rect 68269 45886 68303 45920
rect 68337 45886 68371 45920
rect 68405 45886 68439 45920
rect 68473 45886 68507 45920
rect 68541 45886 68575 45920
rect 68609 45886 68643 45920
rect 68677 45886 68711 45920
rect 68745 45886 68779 45920
rect 68813 45886 68847 45920
rect 68881 45886 68915 45920
rect 68949 45886 68983 45920
rect 69017 45886 69051 45920
rect 69085 45886 69119 45920
rect 69153 45886 69187 45920
rect 69221 45886 69255 45920
rect 69289 45886 69323 45920
rect 69357 45886 69391 45920
rect 69425 45886 69459 45920
rect 69493 45886 69527 45920
rect 69561 45886 69595 45920
rect 69629 45886 69663 45920
rect 69697 45886 69731 45920
rect 69765 45886 69799 45920
rect 69833 45886 69867 45920
rect 69901 45886 69935 45920
rect 69969 45886 70003 45920
rect 70037 45886 70071 45920
rect 70105 45886 70139 45920
rect 70173 45886 70207 45920
rect 70241 45886 70275 45920
rect 70309 45886 70343 45920
rect 70377 45886 70411 45920
rect 70445 45886 70479 45920
rect 70513 45886 70547 45920
rect 70581 45886 70615 45920
rect 70649 45886 70683 45920
rect 70717 45886 70751 45920
rect 70785 45886 70872 45920
rect -3718 45796 -3684 45830
rect -3718 45728 -3684 45762
rect -3718 45660 -3684 45694
rect -3718 45592 -3684 45626
rect -3718 45524 -3684 45558
rect -3718 45456 -3684 45490
rect -3718 45388 -3684 45422
rect -3718 45320 -3684 45354
rect -3718 45252 -3684 45286
rect -3718 45184 -3684 45218
rect -3718 45116 -3684 45150
rect -3718 45048 -3684 45082
rect -3718 44980 -3684 45014
rect -3718 44912 -3684 44946
rect -3718 44844 -3684 44878
rect -3718 44776 -3684 44810
rect -3718 44708 -3684 44742
rect -3718 44640 -3684 44674
rect -3718 44572 -3684 44606
rect -3718 44504 -3684 44538
rect -3718 44436 -3684 44470
rect -3718 44368 -3684 44402
rect -3718 44280 -3684 44334
rect -10699 44246 -10609 44280
rect -10575 44246 -10541 44280
rect -10507 44246 -10473 44280
rect -10439 44246 -10405 44280
rect -10371 44246 -10337 44280
rect -10303 44246 -10269 44280
rect -10235 44246 -10201 44280
rect -10167 44246 -10133 44280
rect -10099 44246 -10065 44280
rect -10031 44246 -9997 44280
rect -9963 44246 -9929 44280
rect -9895 44246 -9861 44280
rect -9827 44246 -9793 44280
rect -9759 44246 -9725 44280
rect -9691 44246 -9657 44280
rect -9623 44246 -9589 44280
rect -9555 44246 -9521 44280
rect -9487 44246 -9453 44280
rect -9419 44246 -9385 44280
rect -9351 44246 -9317 44280
rect -9283 44246 -9249 44280
rect -9215 44246 -9181 44280
rect -9147 44246 -9113 44280
rect -9079 44246 -9045 44280
rect -9011 44246 -8977 44280
rect -8943 44246 -8909 44280
rect -8875 44246 -8841 44280
rect -8807 44246 -8773 44280
rect -8739 44246 -8705 44280
rect -8671 44246 -8637 44280
rect -8603 44246 -8569 44280
rect -8535 44246 -8501 44280
rect -8467 44246 -8433 44280
rect -8399 44246 -8365 44280
rect -8331 44246 -8297 44280
rect -8263 44246 -8229 44280
rect -8195 44246 -8161 44280
rect -8127 44246 -8093 44280
rect -8059 44246 -8025 44280
rect -7991 44246 -7957 44280
rect -7923 44246 -7889 44280
rect -7855 44246 -7821 44280
rect -7787 44246 -7753 44280
rect -7719 44246 -7685 44280
rect -7651 44246 -7617 44280
rect -7583 44246 -7549 44280
rect -7515 44246 -7481 44280
rect -7447 44246 -7413 44280
rect -7379 44246 -7345 44280
rect -7311 44246 -7277 44280
rect -7243 44246 -7209 44280
rect -7175 44246 -7141 44280
rect -7107 44246 -7073 44280
rect -7039 44246 -7005 44280
rect -6971 44246 -6937 44280
rect -6903 44246 -6869 44280
rect -6835 44246 -6801 44280
rect -6767 44246 -6733 44280
rect -6699 44246 -6665 44280
rect -6631 44246 -6597 44280
rect -6563 44246 -6529 44280
rect -6495 44246 -6461 44280
rect -6427 44246 -6393 44280
rect -6359 44246 -6325 44280
rect -6291 44246 -6257 44280
rect -6223 44246 -6189 44280
rect -6155 44246 -6121 44280
rect -6087 44246 -6053 44280
rect -6019 44246 -5985 44280
rect -5951 44246 -5917 44280
rect -5883 44246 -5849 44280
rect -5815 44246 -5781 44280
rect -5747 44246 -5713 44280
rect -5679 44246 -5645 44280
rect -5611 44246 -5577 44280
rect -5543 44246 -5509 44280
rect -5475 44246 -5441 44280
rect -5407 44246 -5373 44280
rect -5339 44246 -5305 44280
rect -5271 44246 -5237 44280
rect -5203 44246 -5169 44280
rect -5135 44246 -5101 44280
rect -5067 44246 -5033 44280
rect -4999 44246 -4965 44280
rect -4931 44246 -4897 44280
rect -4863 44246 -4829 44280
rect -4795 44246 -4761 44280
rect -4727 44246 -4693 44280
rect -4659 44246 -4625 44280
rect -4591 44246 -4557 44280
rect -4523 44246 -4489 44280
rect -4455 44246 -4421 44280
rect -4387 44246 -4353 44280
rect -4319 44246 -4285 44280
rect -4251 44246 -4217 44280
rect -4183 44246 -4149 44280
rect -4115 44246 -4081 44280
rect -4047 44246 -4013 44280
rect -3979 44246 -3945 44280
rect -3911 44246 -3877 44280
rect -3843 44246 -3809 44280
rect -3775 44246 -3684 44280
rect -2396 19487 -2318 19521
rect -2284 19487 -2250 19521
rect -2216 19487 -2182 19521
rect -2148 19487 -2114 19521
rect -2080 19487 -2046 19521
rect -2012 19487 -1978 19521
rect -1944 19487 -1910 19521
rect -1876 19487 -1842 19521
rect -1808 19487 -1774 19521
rect -1740 19487 -1706 19521
rect -1672 19487 -1638 19521
rect -1604 19487 -1570 19521
rect -1536 19487 -1502 19521
rect -1468 19487 -1434 19521
rect -1400 19487 -1366 19521
rect -1332 19487 -1298 19521
rect -1264 19487 -1230 19521
rect -1196 19487 -1162 19521
rect -1128 19487 -1094 19521
rect -1060 19487 -1026 19521
rect -992 19487 -958 19521
rect -924 19487 -890 19521
rect -856 19487 -822 19521
rect -788 19487 -754 19521
rect -720 19487 -686 19521
rect -652 19487 -618 19521
rect -584 19487 -550 19521
rect -516 19487 -482 19521
rect -448 19487 -414 19521
rect -380 19487 -346 19521
rect -312 19487 -278 19521
rect -244 19487 -210 19521
rect -176 19487 -142 19521
rect -108 19487 -74 19521
rect -40 19487 -6 19521
rect 28 19487 62 19521
rect 96 19487 130 19521
rect 164 19487 198 19521
rect 232 19487 266 19521
rect 300 19487 334 19521
rect 368 19487 402 19521
rect 436 19487 470 19521
rect 504 19487 538 19521
rect 572 19487 606 19521
rect 640 19487 674 19521
rect 708 19487 742 19521
rect 776 19487 810 19521
rect 844 19487 878 19521
rect 912 19487 946 19521
rect 980 19487 1014 19521
rect 1048 19487 1082 19521
rect 1116 19487 1150 19521
rect 1184 19487 1218 19521
rect 1252 19487 1286 19521
rect 1320 19487 1354 19521
rect 1388 19487 1422 19521
rect 1456 19487 1490 19521
rect 1524 19487 1558 19521
rect 1592 19487 1626 19521
rect 1660 19487 1694 19521
rect 1728 19487 1762 19521
rect 1796 19487 1830 19521
rect 1864 19487 1898 19521
rect 1932 19487 1966 19521
rect 2000 19487 2034 19521
rect 2068 19487 2102 19521
rect 2136 19487 2170 19521
rect 2204 19487 2238 19521
rect 2272 19487 2306 19521
rect 2340 19487 2374 19521
rect 2408 19487 2442 19521
rect 2476 19487 2510 19521
rect 2544 19487 2578 19521
rect 2612 19487 2646 19521
rect 2680 19487 2714 19521
rect 2748 19487 2782 19521
rect 2816 19487 2850 19521
rect 2884 19487 2918 19521
rect 2952 19487 2986 19521
rect 3020 19487 3054 19521
rect 3088 19487 3122 19521
rect 3156 19487 3190 19521
rect 3224 19487 3258 19521
rect 3292 19487 3326 19521
rect 3360 19487 3394 19521
rect 3428 19487 3462 19521
rect 3496 19487 3530 19521
rect 3564 19487 3598 19521
rect 3632 19487 3666 19521
rect 3700 19487 3734 19521
rect 3768 19487 3802 19521
rect 3836 19487 3870 19521
rect 3904 19487 3938 19521
rect 3972 19487 4006 19521
rect 4040 19487 4074 19521
rect 4108 19487 4142 19521
rect 4176 19487 4210 19521
rect 4244 19487 4278 19521
rect 4312 19487 4346 19521
rect 4380 19487 4414 19521
rect 4448 19487 4482 19521
rect 4516 19487 4550 19521
rect 4584 19487 4618 19521
rect 4652 19487 4686 19521
rect 4720 19487 4754 19521
rect 4788 19487 4822 19521
rect 4856 19487 4890 19521
rect 4924 19487 4958 19521
rect 4992 19487 5026 19521
rect 5060 19487 5094 19521
rect 5128 19487 5162 19521
rect 5196 19487 5230 19521
rect 5264 19487 5298 19521
rect 5332 19487 5366 19521
rect 5400 19487 5434 19521
rect 5468 19487 5502 19521
rect 5536 19487 5570 19521
rect 5604 19487 5638 19521
rect 5672 19487 5706 19521
rect 5740 19487 5774 19521
rect 5808 19487 5842 19521
rect 5876 19487 5910 19521
rect 5944 19487 5978 19521
rect 6012 19487 6046 19521
rect 6080 19487 6114 19521
rect 6148 19487 6182 19521
rect 6216 19487 6250 19521
rect 6284 19487 6318 19521
rect 6352 19487 6386 19521
rect 6420 19487 6454 19521
rect 6488 19487 6522 19521
rect 6556 19487 6590 19521
rect 6624 19487 6658 19521
rect 6692 19487 6726 19521
rect 6760 19487 6794 19521
rect 6828 19487 6862 19521
rect 6896 19487 6930 19521
rect 6964 19487 6998 19521
rect 7032 19487 7066 19521
rect 7100 19487 7134 19521
rect 7168 19487 7202 19521
rect 7236 19487 7270 19521
rect 7304 19487 7338 19521
rect 7372 19487 7406 19521
rect 7440 19487 7474 19521
rect 7508 19487 7542 19521
rect 7576 19487 7610 19521
rect 7644 19487 7678 19521
rect 7712 19487 7746 19521
rect 7780 19487 7814 19521
rect 7848 19487 7882 19521
rect 7916 19487 7950 19521
rect 7984 19487 8018 19521
rect 8052 19487 8086 19521
rect 8120 19487 8154 19521
rect 8188 19487 8222 19521
rect 8256 19487 8290 19521
rect 8324 19487 8358 19521
rect 8392 19487 8426 19521
rect 8460 19487 8494 19521
rect 8528 19487 8562 19521
rect 8596 19487 8630 19521
rect 8664 19487 8698 19521
rect 8732 19487 8766 19521
rect 8800 19487 8834 19521
rect 8868 19487 8902 19521
rect 8936 19487 8970 19521
rect 9004 19487 9038 19521
rect 9072 19487 9106 19521
rect 9140 19487 9174 19521
rect 9208 19487 9242 19521
rect 9276 19487 9310 19521
rect 9344 19487 9378 19521
rect 9412 19487 9446 19521
rect 9480 19487 9514 19521
rect 9548 19487 9582 19521
rect 9616 19487 9650 19521
rect 9684 19487 9718 19521
rect 9752 19487 9786 19521
rect 9820 19487 9854 19521
rect 9888 19487 9922 19521
rect 9956 19487 9990 19521
rect 10024 19487 10058 19521
rect 10092 19487 10126 19521
rect 10160 19487 10194 19521
rect 10228 19487 10262 19521
rect 10296 19487 10330 19521
rect 10364 19487 10398 19521
rect 10432 19487 10466 19521
rect 10500 19487 10534 19521
rect 10568 19487 10602 19521
rect 10636 19487 10670 19521
rect 10704 19487 10738 19521
rect 10772 19487 10806 19521
rect 10840 19487 10874 19521
rect 10908 19487 10942 19521
rect 10976 19487 11010 19521
rect 11044 19487 11078 19521
rect 11112 19487 11146 19521
rect 11180 19487 11214 19521
rect 11248 19487 11282 19521
rect 11316 19487 11350 19521
rect 11384 19487 11418 19521
rect 11452 19487 11486 19521
rect 11520 19487 11554 19521
rect 11588 19487 11622 19521
rect 11656 19487 11690 19521
rect 11724 19487 11758 19521
rect 11792 19487 11826 19521
rect 11860 19487 11894 19521
rect 11928 19487 11962 19521
rect 11996 19487 12030 19521
rect 12064 19487 12098 19521
rect 12132 19487 12166 19521
rect 12200 19487 12234 19521
rect 12268 19487 12302 19521
rect 12336 19487 12370 19521
rect 12404 19487 12438 19521
rect 12472 19487 12506 19521
rect 12540 19487 12574 19521
rect 12608 19487 12642 19521
rect 12676 19487 12710 19521
rect 12744 19487 12778 19521
rect 12812 19487 12846 19521
rect 12880 19487 12914 19521
rect 12948 19487 12982 19521
rect 13016 19487 13050 19521
rect 13084 19487 13118 19521
rect 13152 19487 13186 19521
rect 13220 19487 13254 19521
rect 13288 19487 13322 19521
rect 13356 19487 13390 19521
rect 13424 19487 13458 19521
rect 13492 19487 13526 19521
rect 13560 19487 13594 19521
rect 13628 19487 13662 19521
rect 13696 19487 13730 19521
rect 13764 19487 13798 19521
rect 13832 19487 13866 19521
rect 13900 19487 13934 19521
rect 13968 19487 14002 19521
rect 14036 19487 14070 19521
rect 14104 19487 14138 19521
rect 14172 19487 14206 19521
rect 14240 19487 14274 19521
rect 14308 19487 14342 19521
rect 14376 19487 14410 19521
rect 14444 19487 14478 19521
rect 14512 19487 14546 19521
rect 14580 19487 14614 19521
rect 14648 19487 14682 19521
rect 14716 19487 14750 19521
rect 14784 19487 14818 19521
rect 14852 19487 14886 19521
rect 14920 19487 14954 19521
rect 14988 19487 15022 19521
rect 15056 19487 15090 19521
rect 15124 19487 15158 19521
rect 15192 19487 15226 19521
rect 15260 19487 15294 19521
rect 15328 19487 15362 19521
rect 15396 19487 15430 19521
rect 15464 19487 15498 19521
rect 15532 19487 15566 19521
rect 15600 19487 15634 19521
rect 15668 19487 15702 19521
rect 15736 19487 15770 19521
rect 15804 19487 15838 19521
rect 15872 19487 15906 19521
rect 15940 19487 15974 19521
rect 16008 19487 16042 19521
rect 16076 19487 16110 19521
rect 16144 19487 16178 19521
rect 16212 19487 16246 19521
rect 16280 19487 16314 19521
rect 16348 19487 16382 19521
rect 16416 19487 16450 19521
rect 16484 19487 16518 19521
rect 16552 19487 16586 19521
rect 16620 19487 16654 19521
rect 16688 19487 16722 19521
rect 16756 19487 16790 19521
rect 16824 19487 16858 19521
rect 16892 19487 16926 19521
rect 16960 19487 16994 19521
rect 17028 19487 17062 19521
rect 17096 19487 17130 19521
rect 17164 19487 17198 19521
rect 17232 19487 17266 19521
rect 17300 19487 17334 19521
rect 17368 19487 17402 19521
rect 17436 19487 17470 19521
rect 17504 19487 17538 19521
rect 17572 19487 17606 19521
rect 17640 19487 17674 19521
rect 17708 19487 17742 19521
rect 17776 19487 17810 19521
rect 17844 19487 17878 19521
rect 17912 19487 17946 19521
rect 17980 19487 18014 19521
rect 18048 19487 18082 19521
rect 18116 19487 18150 19521
rect 18184 19487 18218 19521
rect 18252 19487 18286 19521
rect 18320 19487 18354 19521
rect 18388 19487 18422 19521
rect 18456 19487 18490 19521
rect 18524 19487 18558 19521
rect 18592 19487 18626 19521
rect 18660 19487 18694 19521
rect 18728 19487 18762 19521
rect 18796 19487 18830 19521
rect 18864 19487 18898 19521
rect 18932 19487 18966 19521
rect 19000 19487 19034 19521
rect 19068 19487 19102 19521
rect 19136 19487 19170 19521
rect 19204 19487 19238 19521
rect 19272 19487 19306 19521
rect 19340 19487 19374 19521
rect 19408 19487 19442 19521
rect 19476 19487 19510 19521
rect 19544 19487 19578 19521
rect 19612 19487 19646 19521
rect 19680 19487 19714 19521
rect 19748 19487 19782 19521
rect 19816 19487 19850 19521
rect 19884 19487 19918 19521
rect 19952 19487 19986 19521
rect 20020 19487 20054 19521
rect 20088 19487 20122 19521
rect 20156 19487 20190 19521
rect 20224 19487 20258 19521
rect 20292 19487 20326 19521
rect 20360 19487 20394 19521
rect 20428 19487 20462 19521
rect 20496 19487 20530 19521
rect 20564 19487 20598 19521
rect 20632 19487 20666 19521
rect 20700 19487 20734 19521
rect 20768 19487 20802 19521
rect 20836 19487 20870 19521
rect 20904 19487 20938 19521
rect 20972 19487 21006 19521
rect 21040 19487 21074 19521
rect 21108 19487 21142 19521
rect 21176 19487 21210 19521
rect 21244 19487 21278 19521
rect 21312 19487 21346 19521
rect 21380 19487 21414 19521
rect 21448 19487 21482 19521
rect 21516 19487 21550 19521
rect 21584 19487 21618 19521
rect 21652 19487 21686 19521
rect 21720 19487 21754 19521
rect 21788 19487 21822 19521
rect 21856 19487 21890 19521
rect 21924 19487 21958 19521
rect 21992 19487 22026 19521
rect 22060 19487 22094 19521
rect 22128 19487 22162 19521
rect 22196 19487 22230 19521
rect 22264 19487 22298 19521
rect 22332 19487 22366 19521
rect 22400 19487 22434 19521
rect 22468 19487 22502 19521
rect 22536 19487 22570 19521
rect 22604 19487 22638 19521
rect 22672 19487 22706 19521
rect 22740 19487 22774 19521
rect 22808 19487 22842 19521
rect 22876 19487 22910 19521
rect 22944 19487 22978 19521
rect 23012 19487 23046 19521
rect 23080 19487 23114 19521
rect 23148 19487 23182 19521
rect 23216 19487 23250 19521
rect 23284 19487 23318 19521
rect 23352 19487 23386 19521
rect 23420 19487 23454 19521
rect 23488 19487 23522 19521
rect 23556 19487 23590 19521
rect 23624 19487 23658 19521
rect 23692 19487 23726 19521
rect 23760 19487 23794 19521
rect 23828 19487 23862 19521
rect 23896 19487 23930 19521
rect 23964 19487 23998 19521
rect 24032 19487 24066 19521
rect 24100 19487 24134 19521
rect 24168 19487 24202 19521
rect 24236 19487 24270 19521
rect 24304 19487 24338 19521
rect 24372 19487 24406 19521
rect 24440 19487 24474 19521
rect 24508 19487 24542 19521
rect 24576 19487 24610 19521
rect 24644 19487 24678 19521
rect 24712 19487 24746 19521
rect 24780 19487 24814 19521
rect 24848 19487 24882 19521
rect 24916 19487 24950 19521
rect 24984 19487 25018 19521
rect 25052 19487 25086 19521
rect 25120 19487 25154 19521
rect 25188 19487 25222 19521
rect 25256 19487 25290 19521
rect 25324 19487 25358 19521
rect 25392 19487 25426 19521
rect 25460 19487 25494 19521
rect 25528 19487 25562 19521
rect 25596 19487 25630 19521
rect 25664 19487 25698 19521
rect 25732 19487 25766 19521
rect 25800 19487 25834 19521
rect 25868 19487 25902 19521
rect 25936 19487 25970 19521
rect 26004 19487 26038 19521
rect 26072 19487 26106 19521
rect 26140 19487 26174 19521
rect 26208 19487 26242 19521
rect 26276 19487 26310 19521
rect 26344 19487 26378 19521
rect 26412 19487 26446 19521
rect 26480 19487 26514 19521
rect 26548 19487 26582 19521
rect 26616 19487 26650 19521
rect 26684 19487 26718 19521
rect 26752 19487 26786 19521
rect 26820 19487 26854 19521
rect 26888 19487 26922 19521
rect 26956 19487 26990 19521
rect 27024 19487 27058 19521
rect 27092 19487 27126 19521
rect 27160 19487 27194 19521
rect 27228 19487 27262 19521
rect 27296 19487 27330 19521
rect 27364 19487 27398 19521
rect 27432 19487 27466 19521
rect 27500 19487 27534 19521
rect 27568 19487 27602 19521
rect 27636 19487 27670 19521
rect 27704 19487 27738 19521
rect 27772 19487 27806 19521
rect 27840 19487 27874 19521
rect 27908 19487 27942 19521
rect 27976 19487 28010 19521
rect 28044 19487 28078 19521
rect 28112 19487 28146 19521
rect 28180 19487 28214 19521
rect 28248 19487 28282 19521
rect 28316 19487 28350 19521
rect 28384 19487 28418 19521
rect 28452 19487 28486 19521
rect 28520 19487 28554 19521
rect 28588 19487 28622 19521
rect 28656 19487 28690 19521
rect 28724 19487 28758 19521
rect 28792 19487 28826 19521
rect 28860 19487 28894 19521
rect 28928 19487 28962 19521
rect 28996 19487 29030 19521
rect 29064 19487 29098 19521
rect 29132 19487 29166 19521
rect 29200 19487 29234 19521
rect 29268 19487 29302 19521
rect 29336 19487 29370 19521
rect 29404 19487 29438 19521
rect 29472 19487 29506 19521
rect 29540 19487 29574 19521
rect 29608 19487 29642 19521
rect 29676 19487 29710 19521
rect 29744 19487 29778 19521
rect 29812 19487 29846 19521
rect 29880 19487 29914 19521
rect 29948 19487 29982 19521
rect 30016 19487 30050 19521
rect 30084 19487 30118 19521
rect 30152 19487 30186 19521
rect 30220 19487 30254 19521
rect 30288 19487 30322 19521
rect 30356 19487 30390 19521
rect 30424 19487 30458 19521
rect 30492 19487 30526 19521
rect 30560 19487 30594 19521
rect 30628 19487 30662 19521
rect 30696 19487 30730 19521
rect 30764 19487 30798 19521
rect 30832 19487 30866 19521
rect 30900 19487 30934 19521
rect 30968 19487 31002 19521
rect 31036 19487 31070 19521
rect 31104 19487 31138 19521
rect 31172 19487 31206 19521
rect 31240 19487 31274 19521
rect 31308 19487 31342 19521
rect 31376 19487 31410 19521
rect 31444 19487 31478 19521
rect 31512 19487 31546 19521
rect 31580 19487 31614 19521
rect 31648 19487 31682 19521
rect 31716 19487 31750 19521
rect 31784 19487 31818 19521
rect 31852 19487 31886 19521
rect 31920 19487 31954 19521
rect 31988 19487 32022 19521
rect 32056 19487 32090 19521
rect 32124 19487 32158 19521
rect 32192 19487 32226 19521
rect 32260 19487 32294 19521
rect 32328 19487 32362 19521
rect 32396 19487 32430 19521
rect 32464 19487 32498 19521
rect 32532 19487 32566 19521
rect 32600 19487 32634 19521
rect 32668 19487 32702 19521
rect 32736 19487 32770 19521
rect 32804 19487 32838 19521
rect 32872 19487 32906 19521
rect 32940 19487 32974 19521
rect 33008 19487 33042 19521
rect 33076 19487 33110 19521
rect 33144 19487 33178 19521
rect 33212 19487 33246 19521
rect 33280 19487 33314 19521
rect 33348 19487 33382 19521
rect 33416 19487 33450 19521
rect 33484 19487 33518 19521
rect 33552 19487 33586 19521
rect 33620 19487 33654 19521
rect 33688 19487 33722 19521
rect 33756 19487 33790 19521
rect 33824 19487 33858 19521
rect 33892 19487 33926 19521
rect 33960 19487 33994 19521
rect 34028 19487 34062 19521
rect 34096 19487 34130 19521
rect 34164 19487 34198 19521
rect 34232 19487 34266 19521
rect 34300 19487 34334 19521
rect 34368 19487 34402 19521
rect 34436 19487 34470 19521
rect 34504 19487 34538 19521
rect 34572 19487 34606 19521
rect 34640 19487 34674 19521
rect 34708 19487 34742 19521
rect 34776 19487 34810 19521
rect 34844 19487 34878 19521
rect 34912 19487 34946 19521
rect 34980 19487 35014 19521
rect 35048 19487 35082 19521
rect 35116 19487 35150 19521
rect 35184 19487 35218 19521
rect 35252 19487 35286 19521
rect 35320 19487 35354 19521
rect 35388 19487 35422 19521
rect 35456 19487 35490 19521
rect 35524 19487 35558 19521
rect 35592 19487 35626 19521
rect 35660 19487 35694 19521
rect 35728 19487 35762 19521
rect 35796 19487 35830 19521
rect 35864 19487 35898 19521
rect 35932 19487 35966 19521
rect 36000 19487 36034 19521
rect 36068 19487 36102 19521
rect 36136 19487 36170 19521
rect 36204 19487 36238 19521
rect 36272 19487 36306 19521
rect 36340 19487 36374 19521
rect 36408 19487 36442 19521
rect 36476 19487 36510 19521
rect 36544 19487 36578 19521
rect 36612 19487 36646 19521
rect 36680 19487 36714 19521
rect 36748 19487 36782 19521
rect 36816 19487 36850 19521
rect 36884 19487 36918 19521
rect 36952 19487 36986 19521
rect 37020 19487 37054 19521
rect 37088 19487 37122 19521
rect 37156 19487 37190 19521
rect 37224 19487 37258 19521
rect 37292 19487 37326 19521
rect 37360 19487 37394 19521
rect 37428 19487 37462 19521
rect 37496 19487 37530 19521
rect 37564 19487 37598 19521
rect 37632 19487 37666 19521
rect 37700 19487 37734 19521
rect 37768 19487 37802 19521
rect 37836 19487 37870 19521
rect 37904 19487 37938 19521
rect 37972 19487 38006 19521
rect 38040 19487 38074 19521
rect 38108 19487 38142 19521
rect 38176 19487 38210 19521
rect 38244 19487 38278 19521
rect 38312 19487 38346 19521
rect 38380 19487 38414 19521
rect 38448 19487 38482 19521
rect 38516 19487 38550 19521
rect 38584 19487 38618 19521
rect 38652 19487 38686 19521
rect 38720 19487 38754 19521
rect 38788 19487 38822 19521
rect 38856 19487 38890 19521
rect 38924 19487 38958 19521
rect 38992 19487 39026 19521
rect 39060 19487 39094 19521
rect 39128 19487 39162 19521
rect 39196 19487 39230 19521
rect 39264 19487 39298 19521
rect 39332 19487 39366 19521
rect 39400 19487 39434 19521
rect 39468 19487 39502 19521
rect 39536 19487 39570 19521
rect 39604 19487 39638 19521
rect 39672 19487 39706 19521
rect 39740 19487 39774 19521
rect 39808 19487 39842 19521
rect 39876 19487 39910 19521
rect 39944 19487 39978 19521
rect 40012 19487 40046 19521
rect 40080 19487 40114 19521
rect 40148 19487 40182 19521
rect 40216 19487 40250 19521
rect 40284 19487 40318 19521
rect 40352 19487 40386 19521
rect 40420 19487 40454 19521
rect 40488 19487 40522 19521
rect 40556 19487 40590 19521
rect 40624 19487 40658 19521
rect 40692 19487 40726 19521
rect 40760 19487 40794 19521
rect 40828 19487 40862 19521
rect 40896 19487 40930 19521
rect 40964 19487 40998 19521
rect 41032 19487 41066 19521
rect 41100 19487 41134 19521
rect 41168 19487 41202 19521
rect 41236 19487 41270 19521
rect 41304 19487 41338 19521
rect 41372 19487 41406 19521
rect 41440 19487 41474 19521
rect 41508 19487 41542 19521
rect 41576 19487 41610 19521
rect 41644 19487 41678 19521
rect 41712 19487 41746 19521
rect 41780 19487 41814 19521
rect 41848 19487 41882 19521
rect 41916 19487 41950 19521
rect 41984 19487 42018 19521
rect 42052 19487 42086 19521
rect 42120 19487 42154 19521
rect 42188 19487 42222 19521
rect 42256 19487 42290 19521
rect 42324 19487 42358 19521
rect 42392 19487 42426 19521
rect 42460 19487 42494 19521
rect 42528 19487 42562 19521
rect 42596 19487 42630 19521
rect 42664 19487 42698 19521
rect 42732 19487 42766 19521
rect 42800 19487 42834 19521
rect 42868 19487 42902 19521
rect 42936 19487 42970 19521
rect 43004 19487 43038 19521
rect 43072 19487 43106 19521
rect 43140 19487 43174 19521
rect 43208 19487 43242 19521
rect 43276 19487 43310 19521
rect 43344 19487 43378 19521
rect 43412 19487 43446 19521
rect 43480 19487 43514 19521
rect 43548 19487 43582 19521
rect 43616 19487 43650 19521
rect 43684 19487 43718 19521
rect 43752 19487 43786 19521
rect 43820 19487 43854 19521
rect 43888 19487 43922 19521
rect 43956 19487 43990 19521
rect 44024 19487 44058 19521
rect 44092 19487 44126 19521
rect 44160 19487 44194 19521
rect 44228 19487 44262 19521
rect 44296 19487 44330 19521
rect 44364 19487 44398 19521
rect 44432 19487 44466 19521
rect 44500 19487 44534 19521
rect 44568 19487 44602 19521
rect 44636 19487 44670 19521
rect 44704 19487 44738 19521
rect 44772 19487 44806 19521
rect 44840 19487 44874 19521
rect 44908 19487 44942 19521
rect 44976 19487 45010 19521
rect 45044 19487 45078 19521
rect 45112 19487 45146 19521
rect 45180 19487 45214 19521
rect 45248 19487 45282 19521
rect 45316 19487 45350 19521
rect 45384 19487 45418 19521
rect 45452 19487 45486 19521
rect 45520 19487 45554 19521
rect 45588 19487 45622 19521
rect 45656 19487 45690 19521
rect 45724 19487 45758 19521
rect 45792 19487 45826 19521
rect 45860 19487 45894 19521
rect 45928 19487 45962 19521
rect 45996 19487 46030 19521
rect 46064 19487 46098 19521
rect 46132 19487 46166 19521
rect 46200 19487 46234 19521
rect 46268 19487 46302 19521
rect 46336 19487 46370 19521
rect 46404 19487 46438 19521
rect 46472 19487 46506 19521
rect 46540 19487 46574 19521
rect 46608 19487 46642 19521
rect 46676 19487 46710 19521
rect 46744 19487 46778 19521
rect 46812 19487 46846 19521
rect 46880 19487 46914 19521
rect 46948 19487 46982 19521
rect 47016 19487 47050 19521
rect 47084 19487 47118 19521
rect 47152 19487 47230 19521
rect -2396 19434 -2362 19487
rect -2396 19366 -2362 19400
rect -2396 19298 -2362 19332
rect -2396 19230 -2362 19264
rect -2396 19162 -2362 19196
rect -2396 19094 -2362 19128
rect -2396 19026 -2362 19060
rect -2396 18958 -2362 18992
rect -2396 18890 -2362 18924
rect -2396 18822 -2362 18856
rect -2396 18754 -2362 18788
rect -2396 18686 -2362 18720
rect -2396 18618 -2362 18652
rect -2396 18550 -2362 18584
rect -2396 18482 -2362 18516
rect -2396 18414 -2362 18448
rect -2396 18346 -2362 18380
rect -2396 18278 -2362 18312
rect -2396 18210 -2362 18244
rect -2396 18142 -2362 18176
rect -2396 18074 -2362 18108
rect -2396 18006 -2362 18040
rect -2396 17938 -2362 17972
rect -2396 17870 -2362 17904
rect -2396 17802 -2362 17836
rect -2396 17734 -2362 17768
rect -2396 17666 -2362 17700
rect -2396 17598 -2362 17632
rect -2396 17530 -2362 17564
rect -2396 17462 -2362 17496
rect -2396 17394 -2362 17428
rect -2396 17326 -2362 17360
rect -2396 17258 -2362 17292
rect -2396 17190 -2362 17224
rect -2396 17122 -2362 17156
rect -2396 17054 -2362 17088
rect -2396 16986 -2362 17020
rect -2396 16918 -2362 16952
rect -2396 16850 -2362 16884
rect -2396 16782 -2362 16816
rect -2396 16714 -2362 16748
rect -2396 16646 -2362 16680
rect -2396 16578 -2362 16612
rect -2396 16510 -2362 16544
rect -2396 16442 -2362 16476
rect -2396 16374 -2362 16408
rect -2396 16306 -2362 16340
rect -2396 16238 -2362 16272
rect -2396 16170 -2362 16204
rect -2396 16102 -2362 16136
rect -2396 16034 -2362 16068
rect -2396 15966 -2362 16000
rect -2396 15898 -2362 15932
rect -2396 15830 -2362 15864
rect -2396 15762 -2362 15796
rect -2396 15694 -2362 15728
rect -2396 15626 -2362 15660
rect -2396 15558 -2362 15592
rect -2396 15490 -2362 15524
rect -2396 15422 -2362 15456
rect -2396 15354 -2362 15388
rect -2396 15286 -2362 15320
rect -2396 15218 -2362 15252
rect -2396 15150 -2362 15184
rect -2396 15082 -2362 15116
rect -2396 15014 -2362 15048
rect -2396 14946 -2362 14980
rect -2396 14878 -2362 14912
rect -2396 14810 -2362 14844
rect -2396 14742 -2362 14776
rect -2396 14674 -2362 14708
rect -2396 14606 -2362 14640
rect -2396 14538 -2362 14572
rect -2396 14470 -2362 14504
rect -2396 14402 -2362 14436
rect -2396 14334 -2362 14368
rect -2396 14266 -2362 14300
rect -2396 14198 -2362 14232
rect -2396 14130 -2362 14164
rect -2396 14062 -2362 14096
rect -2396 13994 -2362 14028
rect -2396 13926 -2362 13960
rect -2396 13858 -2362 13892
rect -2396 13790 -2362 13824
rect -2396 13722 -2362 13756
rect -2396 13654 -2362 13688
rect -2396 13586 -2362 13620
rect -2396 13518 -2362 13552
rect -2396 13450 -2362 13484
rect -2396 13382 -2362 13416
rect -2396 13314 -2362 13348
rect -2396 13246 -2362 13280
rect -2396 13178 -2362 13212
rect -2396 13110 -2362 13144
rect -2396 13042 -2362 13076
rect -2396 12974 -2362 13008
rect -2396 12906 -2362 12940
rect -2396 12838 -2362 12872
rect -2396 12770 -2362 12804
rect -2396 12702 -2362 12736
rect -2396 12634 -2362 12668
rect -2396 12566 -2362 12600
rect -2396 12498 -2362 12532
rect -2396 12430 -2362 12464
rect -2396 12362 -2362 12396
rect -2396 12294 -2362 12328
rect -2396 12226 -2362 12260
rect -2396 12158 -2362 12192
rect -2396 12090 -2362 12124
rect -2396 12022 -2362 12056
rect -2396 11954 -2362 11988
rect -2396 11886 -2362 11920
rect -2396 11818 -2362 11852
rect -2396 11750 -2362 11784
rect -2396 11682 -2362 11716
rect -2396 11614 -2362 11648
rect -2396 11546 -2362 11580
rect -2396 11478 -2362 11512
rect -2396 11410 -2362 11444
rect -2396 11342 -2362 11376
rect -2396 11274 -2362 11308
rect -2396 11206 -2362 11240
rect -2396 11138 -2362 11172
rect -2396 11070 -2362 11104
rect -2396 11002 -2362 11036
rect -2396 10934 -2362 10968
rect -2396 10866 -2362 10900
rect -2396 10798 -2362 10832
rect -2396 10730 -2362 10764
rect -2396 10662 -2362 10696
rect -2396 10594 -2362 10628
rect -2396 10526 -2362 10560
rect -2396 10458 -2362 10492
rect -2396 10390 -2362 10424
rect -2396 10322 -2362 10356
rect -2396 10254 -2362 10288
rect -2396 10186 -2362 10220
rect -2396 10118 -2362 10152
rect -2396 10050 -2362 10084
rect -2396 9982 -2362 10016
rect -2396 9914 -2362 9948
rect -2396 9846 -2362 9880
rect -2396 9778 -2362 9812
rect -2396 9710 -2362 9744
rect -2396 9642 -2362 9676
rect -2396 9574 -2362 9608
rect -2396 9506 -2362 9540
rect -2396 9438 -2362 9472
rect -2396 9370 -2362 9404
rect -2396 9302 -2362 9336
rect -2396 9234 -2362 9268
rect -2396 9166 -2362 9200
rect -2396 9098 -2362 9132
rect -2396 9030 -2362 9064
rect -2396 8962 -2362 8996
rect -2396 8894 -2362 8928
rect -2396 8826 -2362 8860
rect -2396 8758 -2362 8792
rect -2396 8690 -2362 8724
rect -2396 8622 -2362 8656
rect -2396 8554 -2362 8588
rect -2396 8486 -2362 8520
rect -2396 8418 -2362 8452
rect -2396 8350 -2362 8384
rect -2396 8282 -2362 8316
rect -2396 8214 -2362 8248
rect -2396 8146 -2362 8180
rect -2396 8078 -2362 8112
rect -2396 8010 -2362 8044
rect -2396 7942 -2362 7976
rect -2396 7874 -2362 7908
rect -2396 7806 -2362 7840
rect -2396 7738 -2362 7772
rect -2396 7670 -2362 7704
rect -2396 7602 -2362 7636
rect -2396 7534 -2362 7568
rect -2396 7466 -2362 7500
rect -2396 7398 -2362 7432
rect -2396 7330 -2362 7364
rect -2396 7262 -2362 7296
rect -2396 7194 -2362 7228
rect -2396 7126 -2362 7160
rect -2396 7058 -2362 7092
rect -2396 6990 -2362 7024
rect -2396 6922 -2362 6956
rect -2396 6854 -2362 6888
rect -2396 6786 -2362 6820
rect -2396 6718 -2362 6752
rect -2396 6650 -2362 6684
rect -2396 6582 -2362 6616
rect -2396 6514 -2362 6548
rect -2396 6446 -2362 6480
rect -2396 6378 -2362 6412
rect -2396 6310 -2362 6344
rect -2396 6242 -2362 6276
rect -2396 6174 -2362 6208
rect -2396 6106 -2362 6140
rect -2396 6038 -2362 6072
rect -2396 5970 -2362 6004
rect -2396 5902 -2362 5936
rect -2396 5834 -2362 5868
rect -2396 5766 -2362 5800
rect -2396 5698 -2362 5732
rect -2396 5630 -2362 5664
rect -2396 5562 -2362 5596
rect -2396 5494 -2362 5528
rect -2396 5426 -2362 5460
rect -2396 5358 -2362 5392
rect -2396 5290 -2362 5324
rect -2396 5222 -2362 5256
rect -2396 5154 -2362 5188
rect -2396 5086 -2362 5120
rect -2396 5018 -2362 5052
rect -2396 4950 -2362 4984
rect -2396 4882 -2362 4916
rect -2396 4814 -2362 4848
rect -2396 4746 -2362 4780
rect -2396 4678 -2362 4712
rect -2396 4610 -2362 4644
rect -2396 4542 -2362 4576
rect -2396 4474 -2362 4508
rect -2396 4406 -2362 4440
rect -2396 4338 -2362 4372
rect -2396 4270 -2362 4304
rect -2396 4202 -2362 4236
rect -2396 4134 -2362 4168
rect -2396 4066 -2362 4100
rect -2396 3998 -2362 4032
rect -2396 3930 -2362 3964
rect -2396 3862 -2362 3896
rect -2396 3794 -2362 3828
rect -2396 3726 -2362 3760
rect -2396 3640 -2362 3692
rect 47196 19434 47230 19487
rect 47196 19366 47230 19400
rect 47196 19298 47230 19332
rect 47196 19230 47230 19264
rect 47196 19162 47230 19196
rect 47196 19094 47230 19128
rect 47196 19026 47230 19060
rect 47196 18958 47230 18992
rect 47196 18890 47230 18924
rect 47196 18822 47230 18856
rect 47196 18754 47230 18788
rect 47196 18686 47230 18720
rect 47196 18618 47230 18652
rect 47196 18550 47230 18584
rect 47196 18482 47230 18516
rect 47196 18414 47230 18448
rect 47196 18346 47230 18380
rect 47196 18278 47230 18312
rect 47196 18210 47230 18244
rect 47196 18142 47230 18176
rect 47196 18074 47230 18108
rect 47196 18006 47230 18040
rect 47196 17938 47230 17972
rect 47196 17870 47230 17904
rect 47196 17802 47230 17836
rect 47196 17734 47230 17768
rect 47196 17666 47230 17700
rect 47196 17598 47230 17632
rect 47196 17530 47230 17564
rect 47196 17462 47230 17496
rect 47196 17394 47230 17428
rect 47196 17326 47230 17360
rect 47196 17258 47230 17292
rect 47196 17190 47230 17224
rect 47196 17122 47230 17156
rect 47196 17054 47230 17088
rect 47196 16986 47230 17020
rect 47196 16918 47230 16952
rect 47196 16850 47230 16884
rect 47196 16782 47230 16816
rect 47196 16714 47230 16748
rect 47196 16646 47230 16680
rect 47196 16578 47230 16612
rect 47196 16510 47230 16544
rect 47196 16442 47230 16476
rect 47196 16374 47230 16408
rect 47196 16306 47230 16340
rect 47196 16238 47230 16272
rect 47196 16170 47230 16204
rect 47196 16102 47230 16136
rect 47196 16034 47230 16068
rect 47196 15966 47230 16000
rect 47196 15898 47230 15932
rect 47196 15830 47230 15864
rect 47196 15762 47230 15796
rect 47196 15694 47230 15728
rect 47196 15626 47230 15660
rect 47196 15558 47230 15592
rect 47196 15490 47230 15524
rect 47196 15422 47230 15456
rect 47196 15354 47230 15388
rect 47196 15286 47230 15320
rect 47196 15218 47230 15252
rect 47196 15150 47230 15184
rect 47196 15082 47230 15116
rect 47196 15014 47230 15048
rect 47196 14946 47230 14980
rect 47196 14878 47230 14912
rect 47196 14810 47230 14844
rect 47196 14742 47230 14776
rect 47196 14674 47230 14708
rect 47196 14606 47230 14640
rect 47196 14538 47230 14572
rect 47196 14470 47230 14504
rect 47196 14402 47230 14436
rect 47196 14334 47230 14368
rect 47196 14266 47230 14300
rect 47196 14198 47230 14232
rect 47196 14130 47230 14164
rect 47196 14062 47230 14096
rect 47196 13994 47230 14028
rect 47196 13926 47230 13960
rect 47196 13858 47230 13892
rect 47196 13790 47230 13824
rect 47196 13722 47230 13756
rect 47196 13654 47230 13688
rect 47196 13586 47230 13620
rect 47196 13518 47230 13552
rect 47196 13450 47230 13484
rect 47196 13382 47230 13416
rect 47196 13314 47230 13348
rect 47196 13246 47230 13280
rect 47196 13178 47230 13212
rect 47196 13110 47230 13144
rect 47196 13042 47230 13076
rect 47196 12974 47230 13008
rect 47196 12906 47230 12940
rect 47196 12838 47230 12872
rect 47196 12770 47230 12804
rect 47196 12702 47230 12736
rect 47196 12634 47230 12668
rect 47196 12566 47230 12600
rect 47196 12498 47230 12532
rect 47196 12430 47230 12464
rect 47196 12362 47230 12396
rect 47196 12294 47230 12328
rect 47196 12226 47230 12260
rect 47196 12158 47230 12192
rect 47196 12090 47230 12124
rect 47196 12022 47230 12056
rect 47196 11954 47230 11988
rect 47196 11886 47230 11920
rect 47196 11818 47230 11852
rect 47196 11750 47230 11784
rect 47196 11682 47230 11716
rect 47196 11614 47230 11648
rect 47196 11546 47230 11580
rect 47196 11478 47230 11512
rect 47196 11410 47230 11444
rect 47196 11342 47230 11376
rect 47196 11274 47230 11308
rect 47196 11206 47230 11240
rect 47196 11138 47230 11172
rect 47196 11070 47230 11104
rect 47196 11002 47230 11036
rect 47196 10934 47230 10968
rect 47196 10866 47230 10900
rect 47196 10798 47230 10832
rect 47196 10730 47230 10764
rect 47196 10662 47230 10696
rect 47196 10594 47230 10628
rect 47196 10526 47230 10560
rect 47196 10458 47230 10492
rect 47196 10390 47230 10424
rect 47196 10322 47230 10356
rect 47196 10254 47230 10288
rect 47196 10186 47230 10220
rect 47196 10118 47230 10152
rect 47196 10050 47230 10084
rect 47196 9982 47230 10016
rect 47196 9914 47230 9948
rect 47196 9846 47230 9880
rect 47196 9778 47230 9812
rect 47196 9710 47230 9744
rect 47196 9642 47230 9676
rect 47196 9574 47230 9608
rect 47196 9506 47230 9540
rect 47196 9438 47230 9472
rect 47196 9370 47230 9404
rect 47196 9302 47230 9336
rect 47196 9234 47230 9268
rect 47196 9166 47230 9200
rect 47196 9098 47230 9132
rect 47196 9030 47230 9064
rect 47196 8962 47230 8996
rect 47196 8894 47230 8928
rect 47196 8826 47230 8860
rect 47196 8758 47230 8792
rect 47196 8690 47230 8724
rect 47196 8622 47230 8656
rect 47196 8554 47230 8588
rect 47196 8486 47230 8520
rect 47196 8418 47230 8452
rect 47196 8350 47230 8384
rect 47196 8282 47230 8316
rect 47196 8214 47230 8248
rect 47196 8146 47230 8180
rect 47196 8078 47230 8112
rect 47196 8010 47230 8044
rect 47196 7942 47230 7976
rect 47196 7874 47230 7908
rect 47196 7806 47230 7840
rect 47196 7738 47230 7772
rect 47196 7670 47230 7704
rect 47196 7602 47230 7636
rect 47196 7534 47230 7568
rect 47196 7466 47230 7500
rect 47196 7398 47230 7432
rect 47196 7330 47230 7364
rect 47196 7262 47230 7296
rect 47196 7194 47230 7228
rect 47196 7126 47230 7160
rect 47196 7058 47230 7092
rect 47196 6990 47230 7024
rect 47196 6922 47230 6956
rect 47196 6854 47230 6888
rect 47196 6786 47230 6820
rect 47196 6718 47230 6752
rect 47196 6650 47230 6684
rect 47196 6582 47230 6616
rect 47196 6514 47230 6548
rect 47196 6446 47230 6480
rect 47196 6378 47230 6412
rect 47196 6310 47230 6344
rect 47196 6242 47230 6276
rect 47196 6174 47230 6208
rect 47196 6106 47230 6140
rect 47196 6038 47230 6072
rect 47196 5970 47230 6004
rect 47196 5902 47230 5936
rect 47196 5834 47230 5868
rect 47196 5766 47230 5800
rect 47196 5698 47230 5732
rect 47196 5630 47230 5664
rect 47196 5562 47230 5596
rect 47196 5494 47230 5528
rect 47196 5426 47230 5460
rect 47196 5358 47230 5392
rect 47196 5290 47230 5324
rect 47196 5222 47230 5256
rect 47196 5154 47230 5188
rect 47196 5086 47230 5120
rect 47196 5018 47230 5052
rect 47196 4950 47230 4984
rect 47196 4882 47230 4916
rect 47196 4814 47230 4848
rect 47196 4746 47230 4780
rect 47196 4678 47230 4712
rect 47196 4610 47230 4644
rect 47196 4542 47230 4576
rect 47196 4474 47230 4508
rect 47196 4406 47230 4440
rect 47196 4338 47230 4372
rect 47196 4270 47230 4304
rect 47196 4202 47230 4236
rect 47196 4134 47230 4168
rect 47196 4066 47230 4100
rect 47196 3998 47230 4032
rect 47196 3930 47230 3964
rect 47196 3862 47230 3896
rect 47196 3794 47230 3828
rect 47196 3726 47230 3760
rect 47196 3640 47230 3692
rect -2396 3606 -2318 3640
rect -2284 3606 -2250 3640
rect -2216 3606 -2182 3640
rect -2148 3606 -2114 3640
rect -2080 3606 -2046 3640
rect -2012 3606 -1978 3640
rect -1944 3606 -1910 3640
rect -1876 3606 -1842 3640
rect -1808 3606 -1774 3640
rect -1740 3606 -1706 3640
rect -1672 3606 -1638 3640
rect -1604 3606 -1570 3640
rect -1536 3606 -1502 3640
rect -1468 3606 -1434 3640
rect -1400 3606 -1366 3640
rect -1332 3606 -1298 3640
rect -1264 3606 -1230 3640
rect -1196 3606 -1162 3640
rect -1128 3606 -1094 3640
rect -1060 3606 -1026 3640
rect -992 3606 -958 3640
rect -924 3606 -890 3640
rect -856 3606 -822 3640
rect -788 3606 -754 3640
rect -720 3606 -686 3640
rect -652 3606 -618 3640
rect -584 3606 -550 3640
rect -516 3606 -482 3640
rect -448 3606 -414 3640
rect -380 3606 -346 3640
rect -312 3606 -278 3640
rect -244 3606 -210 3640
rect -176 3606 -142 3640
rect -108 3606 -74 3640
rect -40 3606 -6 3640
rect 28 3606 62 3640
rect 96 3606 130 3640
rect 164 3606 198 3640
rect 232 3606 266 3640
rect 300 3606 334 3640
rect 368 3606 402 3640
rect 436 3606 470 3640
rect 504 3606 538 3640
rect 572 3606 606 3640
rect 640 3606 674 3640
rect 708 3606 742 3640
rect 776 3606 810 3640
rect 844 3606 878 3640
rect 912 3606 946 3640
rect 980 3606 1014 3640
rect 1048 3606 1082 3640
rect 1116 3606 1150 3640
rect 1184 3606 1218 3640
rect 1252 3606 1286 3640
rect 1320 3606 1354 3640
rect 1388 3606 1422 3640
rect 1456 3606 1490 3640
rect 1524 3606 1558 3640
rect 1592 3606 1626 3640
rect 1660 3606 1694 3640
rect 1728 3606 1762 3640
rect 1796 3606 1830 3640
rect 1864 3606 1898 3640
rect 1932 3606 1966 3640
rect 2000 3606 2034 3640
rect 2068 3606 2102 3640
rect 2136 3606 2170 3640
rect 2204 3606 2238 3640
rect 2272 3606 2306 3640
rect 2340 3606 2374 3640
rect 2408 3606 2442 3640
rect 2476 3606 2510 3640
rect 2544 3606 2578 3640
rect 2612 3606 2646 3640
rect 2680 3606 2714 3640
rect 2748 3606 2782 3640
rect 2816 3606 2850 3640
rect 2884 3606 2918 3640
rect 2952 3606 2986 3640
rect 3020 3606 3054 3640
rect 3088 3606 3122 3640
rect 3156 3606 3190 3640
rect 3224 3606 3258 3640
rect 3292 3606 3326 3640
rect 3360 3606 3394 3640
rect 3428 3606 3462 3640
rect 3496 3606 3530 3640
rect 3564 3606 3598 3640
rect 3632 3606 3666 3640
rect 3700 3606 3734 3640
rect 3768 3606 3802 3640
rect 3836 3606 3870 3640
rect 3904 3606 3938 3640
rect 3972 3606 4006 3640
rect 4040 3606 4074 3640
rect 4108 3606 4142 3640
rect 4176 3606 4210 3640
rect 4244 3606 4278 3640
rect 4312 3606 4346 3640
rect 4380 3606 4414 3640
rect 4448 3606 4482 3640
rect 4516 3606 4550 3640
rect 4584 3606 4618 3640
rect 4652 3606 4686 3640
rect 4720 3606 4754 3640
rect 4788 3606 4822 3640
rect 4856 3606 4890 3640
rect 4924 3606 4958 3640
rect 4992 3606 5026 3640
rect 5060 3606 5094 3640
rect 5128 3606 5162 3640
rect 5196 3606 5230 3640
rect 5264 3606 5298 3640
rect 5332 3606 5366 3640
rect 5400 3606 5434 3640
rect 5468 3606 5502 3640
rect 5536 3606 5570 3640
rect 5604 3606 5638 3640
rect 5672 3606 5706 3640
rect 5740 3606 5774 3640
rect 5808 3606 5842 3640
rect 5876 3606 5910 3640
rect 5944 3606 5978 3640
rect 6012 3606 6046 3640
rect 6080 3606 6114 3640
rect 6148 3606 6182 3640
rect 6216 3606 6250 3640
rect 6284 3606 6318 3640
rect 6352 3606 6386 3640
rect 6420 3606 6454 3640
rect 6488 3606 6522 3640
rect 6556 3606 6590 3640
rect 6624 3606 6658 3640
rect 6692 3606 6726 3640
rect 6760 3606 6794 3640
rect 6828 3606 6862 3640
rect 6896 3606 6930 3640
rect 6964 3606 6998 3640
rect 7032 3606 7066 3640
rect 7100 3606 7134 3640
rect 7168 3606 7202 3640
rect 7236 3606 7270 3640
rect 7304 3606 7338 3640
rect 7372 3606 7406 3640
rect 7440 3606 7474 3640
rect 7508 3606 7542 3640
rect 7576 3606 7610 3640
rect 7644 3606 7678 3640
rect 7712 3606 7746 3640
rect 7780 3606 7814 3640
rect 7848 3606 7882 3640
rect 7916 3606 7950 3640
rect 7984 3606 8018 3640
rect 8052 3606 8086 3640
rect 8120 3606 8154 3640
rect 8188 3606 8222 3640
rect 8256 3606 8290 3640
rect 8324 3606 8358 3640
rect 8392 3606 8426 3640
rect 8460 3606 8494 3640
rect 8528 3606 8562 3640
rect 8596 3606 8630 3640
rect 8664 3606 8698 3640
rect 8732 3606 8766 3640
rect 8800 3606 8834 3640
rect 8868 3606 8902 3640
rect 8936 3606 8970 3640
rect 9004 3606 9038 3640
rect 9072 3606 9106 3640
rect 9140 3606 9174 3640
rect 9208 3606 9242 3640
rect 9276 3606 9310 3640
rect 9344 3606 9378 3640
rect 9412 3606 9446 3640
rect 9480 3606 9514 3640
rect 9548 3606 9582 3640
rect 9616 3606 9650 3640
rect 9684 3606 9718 3640
rect 9752 3606 9786 3640
rect 9820 3606 9854 3640
rect 9888 3606 9922 3640
rect 9956 3606 9990 3640
rect 10024 3606 10058 3640
rect 10092 3606 10126 3640
rect 10160 3606 10194 3640
rect 10228 3606 10262 3640
rect 10296 3606 10330 3640
rect 10364 3606 10398 3640
rect 10432 3606 10466 3640
rect 10500 3606 10534 3640
rect 10568 3606 10602 3640
rect 10636 3606 10670 3640
rect 10704 3606 10738 3640
rect 10772 3606 10806 3640
rect 10840 3606 10874 3640
rect 10908 3606 10942 3640
rect 10976 3606 11010 3640
rect 11044 3606 11078 3640
rect 11112 3606 11146 3640
rect 11180 3606 11214 3640
rect 11248 3606 11282 3640
rect 11316 3606 11350 3640
rect 11384 3606 11418 3640
rect 11452 3606 11486 3640
rect 11520 3606 11554 3640
rect 11588 3606 11622 3640
rect 11656 3606 11690 3640
rect 11724 3606 11758 3640
rect 11792 3606 11826 3640
rect 11860 3606 11894 3640
rect 11928 3606 11962 3640
rect 11996 3606 12030 3640
rect 12064 3606 12098 3640
rect 12132 3606 12166 3640
rect 12200 3606 12234 3640
rect 12268 3606 12302 3640
rect 12336 3606 12370 3640
rect 12404 3606 12438 3640
rect 12472 3606 12506 3640
rect 12540 3606 12574 3640
rect 12608 3606 12642 3640
rect 12676 3606 12710 3640
rect 12744 3606 12778 3640
rect 12812 3606 12846 3640
rect 12880 3606 12914 3640
rect 12948 3606 12982 3640
rect 13016 3606 13050 3640
rect 13084 3606 13118 3640
rect 13152 3606 13186 3640
rect 13220 3606 13254 3640
rect 13288 3606 13322 3640
rect 13356 3606 13390 3640
rect 13424 3606 13458 3640
rect 13492 3606 13526 3640
rect 13560 3606 13594 3640
rect 13628 3606 13662 3640
rect 13696 3606 13730 3640
rect 13764 3606 13798 3640
rect 13832 3606 13866 3640
rect 13900 3606 13934 3640
rect 13968 3606 14002 3640
rect 14036 3606 14070 3640
rect 14104 3606 14138 3640
rect 14172 3606 14206 3640
rect 14240 3606 14274 3640
rect 14308 3606 14342 3640
rect 14376 3606 14410 3640
rect 14444 3606 14478 3640
rect 14512 3606 14546 3640
rect 14580 3606 14614 3640
rect 14648 3606 14682 3640
rect 14716 3606 14750 3640
rect 14784 3606 14818 3640
rect 14852 3606 14886 3640
rect 14920 3606 14954 3640
rect 14988 3606 15022 3640
rect 15056 3606 15090 3640
rect 15124 3606 15158 3640
rect 15192 3606 15226 3640
rect 15260 3606 15294 3640
rect 15328 3606 15362 3640
rect 15396 3606 15430 3640
rect 15464 3606 15498 3640
rect 15532 3606 15566 3640
rect 15600 3606 15634 3640
rect 15668 3606 15702 3640
rect 15736 3606 15770 3640
rect 15804 3606 15838 3640
rect 15872 3606 15906 3640
rect 15940 3606 15974 3640
rect 16008 3606 16042 3640
rect 16076 3606 16110 3640
rect 16144 3606 16178 3640
rect 16212 3606 16246 3640
rect 16280 3606 16314 3640
rect 16348 3606 16382 3640
rect 16416 3606 16450 3640
rect 16484 3606 16518 3640
rect 16552 3606 16586 3640
rect 16620 3606 16654 3640
rect 16688 3606 16722 3640
rect 16756 3606 16790 3640
rect 16824 3606 16858 3640
rect 16892 3606 16926 3640
rect 16960 3606 16994 3640
rect 17028 3606 17062 3640
rect 17096 3606 17130 3640
rect 17164 3606 17198 3640
rect 17232 3606 17266 3640
rect 17300 3606 17334 3640
rect 17368 3606 17402 3640
rect 17436 3606 17470 3640
rect 17504 3606 17538 3640
rect 17572 3606 17606 3640
rect 17640 3606 17674 3640
rect 17708 3606 17742 3640
rect 17776 3606 17810 3640
rect 17844 3606 17878 3640
rect 17912 3606 17946 3640
rect 17980 3606 18014 3640
rect 18048 3606 18082 3640
rect 18116 3606 18150 3640
rect 18184 3606 18218 3640
rect 18252 3606 18286 3640
rect 18320 3606 18354 3640
rect 18388 3606 18422 3640
rect 18456 3606 18490 3640
rect 18524 3606 18558 3640
rect 18592 3606 18626 3640
rect 18660 3606 18694 3640
rect 18728 3606 18762 3640
rect 18796 3606 18830 3640
rect 18864 3606 18898 3640
rect 18932 3606 18966 3640
rect 19000 3606 19034 3640
rect 19068 3606 19102 3640
rect 19136 3606 19170 3640
rect 19204 3606 19238 3640
rect 19272 3606 19306 3640
rect 19340 3606 19374 3640
rect 19408 3606 19442 3640
rect 19476 3606 19510 3640
rect 19544 3606 19578 3640
rect 19612 3606 19646 3640
rect 19680 3606 19714 3640
rect 19748 3606 19782 3640
rect 19816 3606 19850 3640
rect 19884 3606 19918 3640
rect 19952 3606 19986 3640
rect 20020 3606 20054 3640
rect 20088 3606 20122 3640
rect 20156 3606 20190 3640
rect 20224 3606 20258 3640
rect 20292 3606 20326 3640
rect 20360 3606 20394 3640
rect 20428 3606 20462 3640
rect 20496 3606 20530 3640
rect 20564 3606 20598 3640
rect 20632 3606 20666 3640
rect 20700 3606 20734 3640
rect 20768 3606 20802 3640
rect 20836 3606 20870 3640
rect 20904 3606 20938 3640
rect 20972 3606 21006 3640
rect 21040 3606 21074 3640
rect 21108 3606 21142 3640
rect 21176 3606 21210 3640
rect 21244 3606 21278 3640
rect 21312 3606 21346 3640
rect 21380 3606 21414 3640
rect 21448 3606 21482 3640
rect 21516 3606 21550 3640
rect 21584 3606 21618 3640
rect 21652 3606 21686 3640
rect 21720 3606 21754 3640
rect 21788 3606 21822 3640
rect 21856 3606 21890 3640
rect 21924 3606 21958 3640
rect 21992 3606 22026 3640
rect 22060 3606 22094 3640
rect 22128 3606 22162 3640
rect 22196 3606 22230 3640
rect 22264 3606 22298 3640
rect 22332 3606 22366 3640
rect 22400 3606 22434 3640
rect 22468 3606 22502 3640
rect 22536 3606 22570 3640
rect 22604 3606 22638 3640
rect 22672 3606 22706 3640
rect 22740 3606 22774 3640
rect 22808 3606 22842 3640
rect 22876 3606 22910 3640
rect 22944 3606 22978 3640
rect 23012 3606 23046 3640
rect 23080 3606 23114 3640
rect 23148 3606 23182 3640
rect 23216 3606 23250 3640
rect 23284 3606 23318 3640
rect 23352 3606 23386 3640
rect 23420 3606 23454 3640
rect 23488 3606 23522 3640
rect 23556 3606 23590 3640
rect 23624 3606 23658 3640
rect 23692 3606 23726 3640
rect 23760 3606 23794 3640
rect 23828 3606 23862 3640
rect 23896 3606 23930 3640
rect 23964 3606 23998 3640
rect 24032 3606 24066 3640
rect 24100 3606 24134 3640
rect 24168 3606 24202 3640
rect 24236 3606 24270 3640
rect 24304 3606 24338 3640
rect 24372 3606 24406 3640
rect 24440 3606 24474 3640
rect 24508 3606 24542 3640
rect 24576 3606 24610 3640
rect 24644 3606 24678 3640
rect 24712 3606 24746 3640
rect 24780 3606 24814 3640
rect 24848 3606 24882 3640
rect 24916 3606 24950 3640
rect 24984 3606 25018 3640
rect 25052 3606 25086 3640
rect 25120 3606 25154 3640
rect 25188 3606 25222 3640
rect 25256 3606 25290 3640
rect 25324 3606 25358 3640
rect 25392 3606 25426 3640
rect 25460 3606 25494 3640
rect 25528 3606 25562 3640
rect 25596 3606 25630 3640
rect 25664 3606 25698 3640
rect 25732 3606 25766 3640
rect 25800 3606 25834 3640
rect 25868 3606 25902 3640
rect 25936 3606 25970 3640
rect 26004 3606 26038 3640
rect 26072 3606 26106 3640
rect 26140 3606 26174 3640
rect 26208 3606 26242 3640
rect 26276 3606 26310 3640
rect 26344 3606 26378 3640
rect 26412 3606 26446 3640
rect 26480 3606 26514 3640
rect 26548 3606 26582 3640
rect 26616 3606 26650 3640
rect 26684 3606 26718 3640
rect 26752 3606 26786 3640
rect 26820 3606 26854 3640
rect 26888 3606 26922 3640
rect 26956 3606 26990 3640
rect 27024 3606 27058 3640
rect 27092 3606 27126 3640
rect 27160 3606 27194 3640
rect 27228 3606 27262 3640
rect 27296 3606 27330 3640
rect 27364 3606 27398 3640
rect 27432 3606 27466 3640
rect 27500 3606 27534 3640
rect 27568 3606 27602 3640
rect 27636 3606 27670 3640
rect 27704 3606 27738 3640
rect 27772 3606 27806 3640
rect 27840 3606 27874 3640
rect 27908 3606 27942 3640
rect 27976 3606 28010 3640
rect 28044 3606 28078 3640
rect 28112 3606 28146 3640
rect 28180 3606 28214 3640
rect 28248 3606 28282 3640
rect 28316 3606 28350 3640
rect 28384 3606 28418 3640
rect 28452 3606 28486 3640
rect 28520 3606 28554 3640
rect 28588 3606 28622 3640
rect 28656 3606 28690 3640
rect 28724 3606 28758 3640
rect 28792 3606 28826 3640
rect 28860 3606 28894 3640
rect 28928 3606 28962 3640
rect 28996 3606 29030 3640
rect 29064 3606 29098 3640
rect 29132 3606 29166 3640
rect 29200 3606 29234 3640
rect 29268 3606 29302 3640
rect 29336 3606 29370 3640
rect 29404 3606 29438 3640
rect 29472 3606 29506 3640
rect 29540 3606 29574 3640
rect 29608 3606 29642 3640
rect 29676 3606 29710 3640
rect 29744 3606 29778 3640
rect 29812 3606 29846 3640
rect 29880 3606 29914 3640
rect 29948 3606 29982 3640
rect 30016 3606 30050 3640
rect 30084 3606 30118 3640
rect 30152 3606 30186 3640
rect 30220 3606 30254 3640
rect 30288 3606 30322 3640
rect 30356 3606 30390 3640
rect 30424 3606 30458 3640
rect 30492 3606 30526 3640
rect 30560 3606 30594 3640
rect 30628 3606 30662 3640
rect 30696 3606 30730 3640
rect 30764 3606 30798 3640
rect 30832 3606 30866 3640
rect 30900 3606 30934 3640
rect 30968 3606 31002 3640
rect 31036 3606 31070 3640
rect 31104 3606 31138 3640
rect 31172 3606 31206 3640
rect 31240 3606 31274 3640
rect 31308 3606 31342 3640
rect 31376 3606 31410 3640
rect 31444 3606 31478 3640
rect 31512 3606 31546 3640
rect 31580 3606 31614 3640
rect 31648 3606 31682 3640
rect 31716 3606 31750 3640
rect 31784 3606 31818 3640
rect 31852 3606 31886 3640
rect 31920 3606 31954 3640
rect 31988 3606 32022 3640
rect 32056 3606 32090 3640
rect 32124 3606 32158 3640
rect 32192 3606 32226 3640
rect 32260 3606 32294 3640
rect 32328 3606 32362 3640
rect 32396 3606 32430 3640
rect 32464 3606 32498 3640
rect 32532 3606 32566 3640
rect 32600 3606 32634 3640
rect 32668 3606 32702 3640
rect 32736 3606 32770 3640
rect 32804 3606 32838 3640
rect 32872 3606 32906 3640
rect 32940 3606 32974 3640
rect 33008 3606 33042 3640
rect 33076 3606 33110 3640
rect 33144 3606 33178 3640
rect 33212 3606 33246 3640
rect 33280 3606 33314 3640
rect 33348 3606 33382 3640
rect 33416 3606 33450 3640
rect 33484 3606 33518 3640
rect 33552 3606 33586 3640
rect 33620 3606 33654 3640
rect 33688 3606 33722 3640
rect 33756 3606 33790 3640
rect 33824 3606 33858 3640
rect 33892 3606 33926 3640
rect 33960 3606 33994 3640
rect 34028 3606 34062 3640
rect 34096 3606 34130 3640
rect 34164 3606 34198 3640
rect 34232 3606 34266 3640
rect 34300 3606 34334 3640
rect 34368 3606 34402 3640
rect 34436 3606 34470 3640
rect 34504 3606 34538 3640
rect 34572 3606 34606 3640
rect 34640 3606 34674 3640
rect 34708 3606 34742 3640
rect 34776 3606 34810 3640
rect 34844 3606 34878 3640
rect 34912 3606 34946 3640
rect 34980 3606 35014 3640
rect 35048 3606 35082 3640
rect 35116 3606 35150 3640
rect 35184 3606 35218 3640
rect 35252 3606 35286 3640
rect 35320 3606 35354 3640
rect 35388 3606 35422 3640
rect 35456 3606 35490 3640
rect 35524 3606 35558 3640
rect 35592 3606 35626 3640
rect 35660 3606 35694 3640
rect 35728 3606 35762 3640
rect 35796 3606 35830 3640
rect 35864 3606 35898 3640
rect 35932 3606 35966 3640
rect 36000 3606 36034 3640
rect 36068 3606 36102 3640
rect 36136 3606 36170 3640
rect 36204 3606 36238 3640
rect 36272 3606 36306 3640
rect 36340 3606 36374 3640
rect 36408 3606 36442 3640
rect 36476 3606 36510 3640
rect 36544 3606 36578 3640
rect 36612 3606 36646 3640
rect 36680 3606 36714 3640
rect 36748 3606 36782 3640
rect 36816 3606 36850 3640
rect 36884 3606 36918 3640
rect 36952 3606 36986 3640
rect 37020 3606 37054 3640
rect 37088 3606 37122 3640
rect 37156 3606 37190 3640
rect 37224 3606 37258 3640
rect 37292 3606 37326 3640
rect 37360 3606 37394 3640
rect 37428 3606 37462 3640
rect 37496 3606 37530 3640
rect 37564 3606 37598 3640
rect 37632 3606 37666 3640
rect 37700 3606 37734 3640
rect 37768 3606 37802 3640
rect 37836 3606 37870 3640
rect 37904 3606 37938 3640
rect 37972 3606 38006 3640
rect 38040 3606 38074 3640
rect 38108 3606 38142 3640
rect 38176 3606 38210 3640
rect 38244 3606 38278 3640
rect 38312 3606 38346 3640
rect 38380 3606 38414 3640
rect 38448 3606 38482 3640
rect 38516 3606 38550 3640
rect 38584 3606 38618 3640
rect 38652 3606 38686 3640
rect 38720 3606 38754 3640
rect 38788 3606 38822 3640
rect 38856 3606 38890 3640
rect 38924 3606 38958 3640
rect 38992 3606 39026 3640
rect 39060 3606 39094 3640
rect 39128 3606 39162 3640
rect 39196 3606 39230 3640
rect 39264 3606 39298 3640
rect 39332 3606 39366 3640
rect 39400 3606 39434 3640
rect 39468 3606 39502 3640
rect 39536 3606 39570 3640
rect 39604 3606 39638 3640
rect 39672 3606 39706 3640
rect 39740 3606 39774 3640
rect 39808 3606 39842 3640
rect 39876 3606 39910 3640
rect 39944 3606 39978 3640
rect 40012 3606 40046 3640
rect 40080 3606 40114 3640
rect 40148 3606 40182 3640
rect 40216 3606 40250 3640
rect 40284 3606 40318 3640
rect 40352 3606 40386 3640
rect 40420 3606 40454 3640
rect 40488 3606 40522 3640
rect 40556 3606 40590 3640
rect 40624 3606 40658 3640
rect 40692 3606 40726 3640
rect 40760 3606 40794 3640
rect 40828 3606 40862 3640
rect 40896 3606 40930 3640
rect 40964 3606 40998 3640
rect 41032 3606 41066 3640
rect 41100 3606 41134 3640
rect 41168 3606 41202 3640
rect 41236 3606 41270 3640
rect 41304 3606 41338 3640
rect 41372 3606 41406 3640
rect 41440 3606 41474 3640
rect 41508 3606 41542 3640
rect 41576 3606 41610 3640
rect 41644 3606 41678 3640
rect 41712 3606 41746 3640
rect 41780 3606 41814 3640
rect 41848 3606 41882 3640
rect 41916 3606 41950 3640
rect 41984 3606 42018 3640
rect 42052 3606 42086 3640
rect 42120 3606 42154 3640
rect 42188 3606 42222 3640
rect 42256 3606 42290 3640
rect 42324 3606 42358 3640
rect 42392 3606 42426 3640
rect 42460 3606 42494 3640
rect 42528 3606 42562 3640
rect 42596 3606 42630 3640
rect 42664 3606 42698 3640
rect 42732 3606 42766 3640
rect 42800 3606 42834 3640
rect 42868 3606 42902 3640
rect 42936 3606 42970 3640
rect 43004 3606 43038 3640
rect 43072 3606 43106 3640
rect 43140 3606 43174 3640
rect 43208 3606 43242 3640
rect 43276 3606 43310 3640
rect 43344 3606 43378 3640
rect 43412 3606 43446 3640
rect 43480 3606 43514 3640
rect 43548 3606 43582 3640
rect 43616 3606 43650 3640
rect 43684 3606 43718 3640
rect 43752 3606 43786 3640
rect 43820 3606 43854 3640
rect 43888 3606 43922 3640
rect 43956 3606 43990 3640
rect 44024 3606 44058 3640
rect 44092 3606 44126 3640
rect 44160 3606 44194 3640
rect 44228 3606 44262 3640
rect 44296 3606 44330 3640
rect 44364 3606 44398 3640
rect 44432 3606 44466 3640
rect 44500 3606 44534 3640
rect 44568 3606 44602 3640
rect 44636 3606 44670 3640
rect 44704 3606 44738 3640
rect 44772 3606 44806 3640
rect 44840 3606 44874 3640
rect 44908 3606 44942 3640
rect 44976 3606 45010 3640
rect 45044 3606 45078 3640
rect 45112 3606 45146 3640
rect 45180 3606 45214 3640
rect 45248 3606 45282 3640
rect 45316 3606 45350 3640
rect 45384 3606 45418 3640
rect 45452 3606 45486 3640
rect 45520 3606 45554 3640
rect 45588 3606 45622 3640
rect 45656 3606 45690 3640
rect 45724 3606 45758 3640
rect 45792 3606 45826 3640
rect 45860 3606 45894 3640
rect 45928 3606 45962 3640
rect 45996 3606 46030 3640
rect 46064 3606 46098 3640
rect 46132 3606 46166 3640
rect 46200 3606 46234 3640
rect 46268 3606 46302 3640
rect 46336 3606 46370 3640
rect 46404 3606 46438 3640
rect 46472 3606 46506 3640
rect 46540 3606 46574 3640
rect 46608 3606 46642 3640
rect 46676 3606 46710 3640
rect 46744 3606 46778 3640
rect 46812 3606 46846 3640
rect 46880 3606 46914 3640
rect 46948 3606 46982 3640
rect 47016 3606 47050 3640
rect 47084 3606 47118 3640
rect 47152 3606 47230 3640
<< metal1 >>
rect -11103 122091 71105 122097
rect -11103 121847 61093 122091
rect 61465 121847 67093 122091
rect 67465 121847 71105 122091
rect -11103 121841 71105 121847
rect -11103 121579 71105 121585
rect -11103 121527 -10558 121579
rect -10506 121527 -3878 121579
rect -3826 121527 50511 121579
rect 50563 121527 56043 121579
rect 56095 121527 71105 121579
rect -11103 121515 71105 121527
rect -11103 121463 -10558 121515
rect -10506 121463 -3878 121515
rect -3826 121463 50511 121515
rect 50563 121463 56043 121515
rect 56095 121463 71105 121515
rect -11103 121451 71105 121463
rect -11103 121399 -10558 121451
rect -10506 121399 -3878 121451
rect -3826 121399 50511 121451
rect 50563 121399 56043 121451
rect 56095 121399 71105 121451
rect -11103 121387 71105 121399
rect -11103 121335 -10558 121387
rect -10506 121335 -3878 121387
rect -3826 121335 50511 121387
rect 50563 121335 56043 121387
rect 56095 121335 71105 121387
rect -11103 121329 71105 121335
rect -11103 121066 71105 121072
rect -11103 120822 46789 121066
rect 46905 120822 71105 121066
rect -11103 120816 71105 120822
rect -2083 115221 -1943 120816
rect -1333 120537 70157 120561
rect -1333 120485 70093 120537
rect 70145 120485 70157 120537
rect -1333 120461 70157 120485
rect -1333 118607 -1233 120461
rect 3469 120337 69005 120361
rect 3469 120285 68941 120337
rect 68993 120285 69005 120337
rect 3469 120261 69005 120285
rect 3469 118690 3569 120261
rect 8271 120137 67853 120161
rect 8271 120085 67789 120137
rect 67841 120085 67853 120137
rect 8271 120061 67853 120085
rect 8271 118659 8371 120061
rect 13073 119937 66701 119961
rect 13073 119885 66637 119937
rect 66689 119885 66701 119937
rect 13073 119861 66701 119885
rect 13073 118671 13173 119861
rect 17875 119737 65549 119761
rect 17875 119685 65485 119737
rect 65537 119685 65549 119737
rect 17875 119661 65549 119685
rect 17875 118665 17975 119661
rect 22677 119537 64397 119561
rect 22677 119485 64333 119537
rect 64385 119485 64397 119537
rect 22677 119461 64397 119485
rect 22677 118632 22777 119461
rect 27479 119337 63245 119361
rect 27479 119285 63181 119337
rect 63233 119285 63245 119337
rect 27479 119261 63245 119285
rect 27479 118674 27579 119261
rect 32281 119137 62093 119161
rect 32281 119085 62029 119137
rect 62081 119085 62093 119137
rect 32281 119061 62093 119085
rect 32281 118632 32381 119061
rect 37083 118937 60941 118961
rect 37083 118885 60877 118937
rect 60929 118885 60941 118937
rect 37083 118861 60941 118885
rect 37083 118613 37183 118861
rect 41885 118737 59789 118761
rect 41885 118685 59725 118737
rect 59777 118685 59789 118737
rect 41885 118661 59789 118685
rect -2093 115209 -1933 115221
rect -2093 115093 -2071 115209
rect -1955 115093 -1933 115209
rect -2093 115081 -1933 115093
rect -10590 76099 -10474 76121
rect -10590 76047 -10558 76099
rect -10506 76047 -10474 76099
rect -10590 76025 -10474 76047
rect -4251 67457 -4241 67509
rect -4189 67457 -4179 67509
rect 614 61885 50056 61900
rect 614 61819 644 61885
rect -4692 61577 644 61819
rect 44472 61833 49994 61885
rect 50046 61833 50056 61885
rect 44472 61821 50056 61833
rect 44472 61769 49994 61821
rect 50046 61769 50056 61821
rect 44472 61757 50056 61769
rect 44472 61705 49994 61757
rect 50046 61705 50056 61757
rect 44472 61693 50056 61705
rect 44472 61641 49994 61693
rect 50046 61641 50056 61693
rect 44472 61629 50056 61641
rect 44472 61577 49994 61629
rect 50046 61577 50056 61629
rect -4692 61563 50056 61577
rect -3739 61429 49335 61435
rect -3739 61377 -3723 61429
rect -3671 61377 49267 61429
rect 49319 61377 49335 61429
rect -3739 61371 49335 61377
rect -4576 60656 50787 60678
rect -4576 60604 -4544 60656
rect -4492 60604 50703 60656
rect 50755 60604 50787 60656
rect -4576 60582 50787 60604
rect 50367 60347 50377 60399
rect 50429 60390 50439 60399
rect 50429 60356 50623 60390
rect 50429 60347 50439 60356
rect 49984 60282 49994 60334
rect 50046 60316 50056 60334
rect 50046 60282 50737 60316
rect 49984 60048 49994 60100
rect 50046 60066 50538 60100
rect 50046 60048 50056 60066
rect 55955 59899 58409 59939
rect 58397 59887 58409 59899
rect 58461 59887 58473 59939
rect 58525 59887 58537 59939
rect -3911 59852 50595 59874
rect -3911 59800 -3879 59852
rect -3827 59800 50511 59852
rect 50563 59800 50595 59852
rect -3911 59778 50595 59800
rect 58637 59727 58649 59779
rect 58701 59727 58713 59779
rect 58765 59727 58777 59779
rect 55964 59687 58777 59727
rect 55930 59608 58777 59648
rect 58637 59556 58649 59608
rect 58701 59556 58713 59608
rect 58765 59556 58777 59608
rect -3739 59013 49336 59019
rect -3739 58961 -3723 59013
rect -3671 58961 49268 59013
rect 49320 58961 49336 59013
rect -3739 58955 49336 58961
rect -4704 58812 50056 58827
rect -4704 58571 644 58812
rect 614 58504 644 58571
rect 44472 58760 49994 58812
rect 50046 58760 50056 58812
rect 44472 58748 50056 58760
rect 44472 58696 49994 58748
rect 50046 58696 50056 58748
rect 44472 58684 50056 58696
rect 44472 58632 49994 58684
rect 50046 58632 50056 58684
rect 44472 58620 50056 58632
rect 44472 58568 49994 58620
rect 50046 58568 50056 58620
rect 44472 58556 50056 58568
rect 44472 58504 49994 58556
rect 50046 58504 50056 58556
rect 614 58490 50056 58504
rect -4251 52881 -4241 52933
rect -4189 52881 -4179 52933
rect -4576 44343 -4460 44365
rect -4576 44291 -4544 44343
rect -4492 44291 -4460 44343
rect -4576 44269 -4460 44291
rect -10590 44073 -3206 44075
rect -10590 43957 -3334 44073
rect -3218 43957 -3206 44073
rect -10590 43955 -3206 43957
rect -10590 43833 -2212 43835
rect -10590 43717 -2350 43833
rect -2234 43717 -2212 43833
rect -10590 43715 -2212 43717
rect -10590 43593 -3339 43595
rect -10590 43477 -3467 43593
rect -3351 43477 -3339 43593
rect -10590 43475 -3339 43477
rect -1813 5497 -1653 5509
rect -1813 5381 -1791 5497
rect -1675 5381 -1653 5497
rect -1813 5369 -1653 5381
rect -1803 -432 -1663 5369
rect -1332 -76 -1232 1737
rect 3470 124 3570 1737
rect 8272 324 8372 1698
rect 13074 524 13174 1688
rect 17876 724 17976 1748
rect 22678 924 22778 1743
rect 27480 1124 27580 1798
rect 41886 1700 59789 1724
rect 32282 1324 32382 1700
rect 37084 1524 37184 1680
rect 41886 1648 59725 1700
rect 59777 1648 59789 1700
rect 41886 1624 59789 1648
rect 37084 1500 60941 1524
rect 37084 1448 60877 1500
rect 60929 1448 60941 1500
rect 37084 1424 60941 1448
rect 32282 1300 62093 1324
rect 32282 1248 62029 1300
rect 62081 1248 62093 1300
rect 32282 1224 62093 1248
rect 27480 1100 63245 1124
rect 27480 1048 63181 1100
rect 63233 1048 63245 1100
rect 27480 1024 63245 1048
rect 22678 900 64397 924
rect 22678 848 64333 900
rect 64385 848 64397 900
rect 22678 824 64397 848
rect 17876 700 65549 724
rect 17876 648 65485 700
rect 65537 648 65549 700
rect 17876 624 65549 648
rect 13074 500 66701 524
rect 13074 448 66637 500
rect 66689 448 66701 500
rect 13074 424 66701 448
rect 8272 300 67853 324
rect 8272 248 67789 300
rect 67841 248 67853 300
rect 8272 224 67853 248
rect 3470 100 69005 124
rect 3470 48 68941 100
rect 68993 48 69005 100
rect 3470 24 69005 48
rect -1332 -100 70157 -76
rect -1332 -152 70093 -100
rect 70145 -152 70157 -100
rect -1332 -176 70157 -152
rect -11102 -438 71106 -432
rect -11102 -682 46509 -438
rect 46625 -682 71106 -438
rect -11102 -688 71106 -682
rect -11102 -950 71106 -944
rect -11102 -1002 -4544 -950
rect -4492 -1002 50703 -950
rect 50755 -1002 55851 -950
rect 55903 -1002 71106 -950
rect -11102 -1014 71106 -1002
rect -11102 -1066 -4544 -1014
rect -4492 -1066 50703 -1014
rect 50755 -1066 55851 -1014
rect 55903 -1066 71106 -1014
rect -11102 -1078 71106 -1066
rect -11102 -1130 -4544 -1078
rect -4492 -1130 50703 -1078
rect 50755 -1130 55851 -1078
rect 55903 -1130 71106 -1078
rect -11102 -1142 71106 -1130
rect -11102 -1194 -4544 -1142
rect -4492 -1194 50703 -1142
rect 50755 -1194 55851 -1142
rect 55903 -1194 71106 -1142
rect -11102 -1200 71106 -1194
rect -11102 -1463 71106 -1457
rect -11102 -1707 64093 -1463
rect 64465 -1707 71106 -1463
rect -11102 -1713 71106 -1707
<< via1 >>
rect 61093 121847 61465 122091
rect 67093 121847 67465 122091
rect -10558 121527 -10506 121579
rect -3878 121527 -3826 121579
rect 50511 121527 50563 121579
rect 56043 121527 56095 121579
rect -10558 121463 -10506 121515
rect -3878 121463 -3826 121515
rect 50511 121463 50563 121515
rect 56043 121463 56095 121515
rect -10558 121399 -10506 121451
rect -3878 121399 -3826 121451
rect 50511 121399 50563 121451
rect 56043 121399 56095 121451
rect -10558 121335 -10506 121387
rect -3878 121335 -3826 121387
rect 50511 121335 50563 121387
rect 56043 121335 56095 121387
rect 46789 120822 46905 121066
rect 70093 120485 70145 120537
rect 68941 120285 68993 120337
rect 67789 120085 67841 120137
rect 66637 119885 66689 119937
rect 65485 119685 65537 119737
rect 64333 119485 64385 119537
rect 63181 119285 63233 119337
rect 62029 119085 62081 119137
rect 60877 118885 60929 118937
rect 59725 118685 59777 118737
rect -2071 115093 -1955 115209
rect -10558 76047 -10506 76099
rect -4241 67457 -4189 67509
rect 644 61577 44472 61885
rect 49994 61833 50046 61885
rect 49994 61769 50046 61821
rect 49994 61705 50046 61757
rect 49994 61641 50046 61693
rect 49994 61577 50046 61629
rect -3723 61377 -3671 61429
rect 49267 61377 49319 61429
rect -4544 60604 -4492 60656
rect 50703 60604 50755 60656
rect 50377 60347 50429 60399
rect 49994 60282 50046 60334
rect 49994 60048 50046 60100
rect 58409 59887 58461 59939
rect 58473 59887 58525 59939
rect -3879 59800 -3827 59852
rect 50511 59800 50563 59852
rect 58649 59727 58701 59779
rect 58713 59727 58765 59779
rect 58649 59556 58701 59608
rect 58713 59556 58765 59608
rect -3723 58961 -3671 59013
rect 49268 58961 49320 59013
rect 644 58504 44472 58812
rect 49994 58760 50046 58812
rect 49994 58696 50046 58748
rect 49994 58632 50046 58684
rect 49994 58568 50046 58620
rect 49994 58504 50046 58556
rect -4241 52881 -4189 52933
rect -4544 44291 -4492 44343
rect -3334 43957 -3218 44073
rect -2350 43717 -2234 43833
rect -3467 43477 -3351 43593
rect -1791 5381 -1675 5497
rect 59725 1648 59777 1700
rect 60877 1448 60929 1500
rect 62029 1248 62081 1300
rect 63181 1048 63233 1100
rect 64333 848 64385 900
rect 65485 648 65537 700
rect 66637 448 66689 500
rect 67789 248 67841 300
rect 68941 48 68993 100
rect 70093 -152 70145 -100
rect 46509 -682 46625 -438
rect -4544 -1002 -4492 -950
rect 50703 -1002 50755 -950
rect 55851 -1002 55903 -950
rect -4544 -1066 -4492 -1014
rect 50703 -1066 50755 -1014
rect 55851 -1066 55903 -1014
rect -4544 -1130 -4492 -1078
rect 50703 -1130 50755 -1078
rect 55851 -1130 55903 -1078
rect -4544 -1194 -4492 -1142
rect 50703 -1194 50755 -1142
rect 55851 -1194 55903 -1142
rect 64093 -1707 64465 -1463
<< metal2 >>
rect 61079 122091 61479 122107
rect 61079 122077 61093 122091
rect 61465 122077 61479 122091
rect 61079 121861 61091 122077
rect 61467 121861 61479 122077
rect 61079 121847 61093 121861
rect 61465 121847 61479 121861
rect 61079 121831 61479 121847
rect 67079 122091 67479 122107
rect 67079 122077 67093 122091
rect 67465 122077 67479 122091
rect 67079 121861 67091 122077
rect 67467 121861 67479 122077
rect 67079 121847 67093 121861
rect 67465 121847 67479 121861
rect 67079 121831 67479 121847
rect -10580 121579 -10484 121595
rect -10580 121527 -10558 121579
rect -10506 121527 -10484 121579
rect -10580 121515 -10484 121527
rect -10580 121463 -10558 121515
rect -10506 121463 -10484 121515
rect -10580 121451 -10484 121463
rect -10580 121399 -10558 121451
rect -10506 121399 -10484 121451
rect -10580 121387 -10484 121399
rect -10580 121335 -10558 121387
rect -10506 121335 -10484 121387
rect -10580 76099 -10484 121335
rect -3901 121579 -3803 121595
rect -3901 121565 -3878 121579
rect -3826 121565 -3803 121579
rect -3901 121509 -3880 121565
rect -3824 121509 -3803 121565
rect -3901 121485 -3878 121509
rect -3826 121485 -3803 121509
rect -3901 121429 -3880 121485
rect -3824 121429 -3803 121485
rect -3901 121405 -3878 121429
rect -3826 121405 -3803 121429
rect -3901 121349 -3880 121405
rect -3824 121349 -3803 121405
rect -3901 121335 -3878 121349
rect -3826 121335 -3803 121349
rect -3901 121319 -3803 121335
rect 50489 121579 50585 121595
rect 50489 121527 50511 121579
rect 50563 121527 50585 121579
rect 50489 121515 50585 121527
rect 50489 121463 50511 121515
rect 50563 121463 50585 121515
rect 50489 121451 50585 121463
rect 50489 121399 50511 121451
rect 50563 121399 50585 121451
rect 50489 121387 50585 121399
rect 50489 121335 50511 121387
rect 50563 121335 50585 121387
rect 46777 121066 46917 121082
rect 46777 121052 46789 121066
rect 46905 121052 46917 121066
rect 46777 120836 46779 121052
rect 46915 120836 46917 121052
rect 46777 120822 46789 120836
rect 46905 120822 46917 120836
rect 46777 120806 46917 120822
rect -2083 115209 -1943 115231
rect -2083 115093 -2071 115209
rect -1955 115093 -1943 115209
rect -2083 115071 -1943 115093
rect 46777 115219 46917 115231
rect 46777 115083 46779 115219
rect 46915 115083 46917 115219
rect 46777 115071 46917 115083
rect -10580 76047 -10558 76099
rect -10506 76047 -10484 76099
rect -10580 76015 -10484 76047
rect 49261 72059 49325 72101
rect 49261 72003 49265 72059
rect 49321 72003 49325 72059
rect 49097 69099 49217 69141
rect 49097 69043 49129 69099
rect 49185 69043 49217 69099
rect 49097 69001 49217 69043
rect 48897 67619 49017 67661
rect 48897 67563 48929 67619
rect 48985 67563 49017 67619
rect -4241 67509 -4189 67519
rect -3729 67511 -3665 67525
rect 48897 67521 49017 67563
rect -3729 67509 -3725 67511
rect -4189 67457 -3725 67509
rect -4241 67447 -4189 67457
rect -3729 67455 -3725 67457
rect -3669 67509 -3665 67511
rect -3669 67457 -3621 67509
rect -3669 67455 -3665 67457
rect -3729 67441 -3665 67455
rect 48697 66139 48817 66181
rect 48697 66083 48729 66139
rect 48785 66083 48817 66139
rect 48697 66041 48817 66083
rect 48497 64659 48617 64701
rect 48497 64603 48529 64659
rect 48585 64603 48617 64659
rect 48497 64561 48617 64603
rect 48297 63179 48417 63221
rect 48297 63123 48329 63179
rect 48385 63123 48417 63179
rect 48297 63081 48417 63123
rect 48097 62579 48217 62621
rect 48097 62523 48129 62579
rect 48185 62523 48217 62579
rect 48097 62481 48217 62523
rect 624 61885 44492 61910
rect 624 61577 644 61885
rect 44472 61577 44492 61885
rect 624 61553 44492 61577
rect -3729 61431 -3665 61445
rect -3729 61375 -3725 61431
rect -3669 61375 -3665 61431
rect -3729 61361 -3665 61375
rect 49261 61429 49325 72003
rect 49261 61377 49267 61429
rect 49319 61377 49325 61429
rect 49261 61361 49325 61377
rect 49994 61885 50046 61910
rect 49994 61821 50046 61833
rect 49994 61757 50046 61769
rect 50489 61753 50585 121335
rect 56021 121579 56117 121595
rect 56021 121527 56043 121579
rect 56095 121527 56117 121579
rect 56021 121515 56117 121527
rect 56021 121463 56043 121515
rect 56095 121463 56117 121515
rect 56021 121451 56117 121463
rect 56021 121399 56043 121451
rect 56095 121399 56117 121451
rect 56021 121387 56117 121399
rect 56021 121335 56043 121387
rect 56095 121335 56117 121387
rect 56021 61765 56117 121335
rect 70091 120537 70147 120571
rect 70091 120485 70093 120537
rect 70145 120485 70147 120537
rect 68939 120337 68995 120371
rect 68939 120285 68941 120337
rect 68993 120285 68995 120337
rect 67787 120137 67843 120171
rect 67787 120085 67789 120137
rect 67841 120085 67843 120137
rect 66635 119937 66691 119971
rect 66635 119885 66637 119937
rect 66689 119885 66691 119937
rect 65483 119737 65539 119771
rect 65483 119685 65485 119737
rect 65537 119685 65539 119737
rect 64331 119537 64387 119571
rect 64331 119485 64333 119537
rect 64385 119485 64387 119537
rect 63179 119337 63235 119371
rect 63179 119285 63181 119337
rect 63233 119285 63235 119337
rect 62027 119137 62083 119171
rect 62027 119085 62029 119137
rect 62081 119085 62083 119137
rect 60875 118937 60931 118971
rect 60875 118885 60877 118937
rect 60929 118885 60931 118937
rect 59723 118737 59779 118771
rect 59723 118685 59725 118737
rect 59777 118685 59779 118737
rect 59723 74724 59779 118685
rect 60875 74579 60931 118885
rect 62027 74727 62083 119085
rect 63179 74697 63235 119285
rect 64331 74694 64387 119485
rect 65483 74727 65539 119685
rect 66635 74707 66691 119885
rect 67787 74718 67843 120085
rect 68939 74701 68995 120285
rect 70091 74726 70147 120485
rect 58647 70579 58767 70621
rect 58647 70523 58679 70579
rect 58735 70523 58767 70579
rect 49994 61693 50046 61705
rect 49994 61629 50046 61641
rect -4566 60658 -4470 60688
rect -4566 60602 -4546 60658
rect -4490 60602 -4470 60658
rect -4566 60572 -4470 60602
rect 49994 60334 50046 61577
rect 50681 60656 50777 60688
rect 50681 60604 50703 60656
rect 50755 60604 50777 60656
rect 50681 60572 50777 60604
rect 49994 60272 50046 60282
rect 50377 60399 50429 60409
rect 50377 60234 50429 60347
rect -3280 60220 -3216 60234
rect -3280 60164 -3276 60220
rect -3220 60164 -3216 60220
rect -3901 59854 -3805 59884
rect -3901 59798 -3881 59854
rect -3825 59798 -3805 59854
rect -3901 59768 -3805 59798
rect -3729 59015 -3665 59029
rect -3729 58959 -3725 59015
rect -3669 58959 -3665 59015
rect -3729 58945 -3665 58959
rect -4241 52933 -4189 52943
rect -3729 52935 -3665 52949
rect -3729 52933 -3725 52935
rect -4189 52881 -3725 52933
rect -4241 52871 -4189 52881
rect -3729 52879 -3725 52881
rect -3669 52879 -3665 52935
rect -3729 52865 -3665 52879
rect -4566 44343 -4470 44375
rect -4566 44291 -4544 44343
rect -4492 44291 -4470 44343
rect -4566 -950 -4470 44291
rect -3280 44085 -3216 60164
rect 50365 60220 50429 60234
rect 50365 60164 50369 60220
rect 50425 60164 50429 60220
rect 50365 60150 50429 60164
rect 49994 60100 50046 60110
rect 49262 59013 49326 59029
rect 49262 58961 49268 59013
rect 49320 58961 49326 59013
rect 624 58812 44492 58837
rect 624 58504 644 58812
rect 44472 58504 44492 58812
rect 624 58480 44492 58504
rect 47898 58219 48018 58261
rect 47898 58163 47930 58219
rect 47986 58163 48018 58219
rect 47898 58121 48018 58163
rect 47698 57859 47818 57901
rect 47698 57803 47730 57859
rect 47786 57803 47818 57859
rect 47698 57761 47818 57803
rect 47498 57259 47618 57301
rect 47498 57203 47530 57259
rect 47586 57203 47618 57259
rect 47498 57161 47618 57203
rect 47298 55779 47418 55821
rect 47298 55723 47330 55779
rect 47386 55723 47418 55779
rect 47298 55681 47418 55723
rect 49262 48379 49326 58961
rect 49994 58812 50046 60048
rect 49994 58748 50046 58760
rect 49994 58684 50046 58696
rect 49994 58620 50046 58632
rect 49994 58556 50046 58568
rect 49994 58480 50046 58504
rect 50377 51381 50429 60150
rect 58407 59939 58527 59949
rect 58407 59887 58409 59939
rect 58461 59887 58473 59939
rect 58525 59887 58527 59939
rect 50489 59852 50585 59884
rect 50489 59800 50511 59852
rect 50563 59800 50585 59852
rect 50489 59768 50585 59800
rect 50375 51339 50431 51381
rect 50375 51241 50431 51283
rect 49262 48323 49266 48379
rect 49322 48323 49326 48379
rect 49262 48281 49326 48323
rect 49686 49859 49806 49901
rect 49686 49803 49718 49859
rect 49774 49803 49806 49859
rect -3336 44073 -3216 44085
rect -3336 43957 -3334 44073
rect -3218 43957 -3216 44073
rect -3336 43945 -3216 43957
rect -2362 43833 -2222 43845
rect -2362 43717 -2350 43833
rect -2234 43717 -2222 43833
rect -2362 43705 -2222 43717
rect -3469 43593 -3349 43605
rect -3469 43477 -3467 43593
rect -3351 43477 -3349 43593
rect -3469 43465 -3349 43477
rect -1803 5497 -1663 5519
rect -1803 5381 -1791 5497
rect -1675 5381 -1663 5497
rect -1803 5359 -1663 5381
rect 46497 5507 46638 5520
rect 46497 5371 46499 5507
rect 46635 5371 46638 5507
rect 46497 5359 46638 5371
rect -3469 -240 -3349 -230
rect 49686 -240 49806 49803
rect -3469 -272 49806 -240
rect -3469 -328 -3437 -272
rect -3381 -328 49806 -272
rect -3469 -360 49806 -328
rect -3469 -370 -3349 -360
rect 46497 -438 46638 -422
rect 46497 -452 46509 -438
rect 46625 -452 46638 -438
rect 46497 -668 46499 -452
rect 46635 -668 46638 -452
rect 46497 -682 46509 -668
rect 46625 -682 46638 -668
rect 46497 -698 46638 -682
rect -4566 -1002 -4544 -950
rect -4492 -1002 -4470 -950
rect -4566 -1014 -4470 -1002
rect -4566 -1066 -4544 -1014
rect -4492 -1066 -4470 -1014
rect -4566 -1078 -4470 -1066
rect -4566 -1130 -4544 -1078
rect -4492 -1130 -4470 -1078
rect -4566 -1142 -4470 -1130
rect -4566 -1194 -4544 -1142
rect -4492 -1194 -4470 -1142
rect -4566 -1210 -4470 -1194
rect 50681 -950 50777 59494
rect 50681 -1002 50703 -950
rect 50755 -1002 50777 -950
rect 50681 -1014 50777 -1002
rect 50681 -1066 50703 -1014
rect 50755 -1066 50777 -1014
rect 50681 -1078 50777 -1066
rect 50681 -1130 50703 -1078
rect 50755 -1130 50777 -1078
rect 50681 -1142 50777 -1130
rect 50681 -1194 50703 -1142
rect 50755 -1194 50777 -1142
rect 50681 -1210 50777 -1194
rect 55829 -950 55925 58910
rect 58407 52819 58527 59887
rect 58647 59779 58767 70523
rect 59127 62579 59247 62621
rect 59127 62523 59159 62579
rect 59215 62523 59247 62579
rect 59127 61699 59247 62523
rect 59127 61643 59159 61699
rect 59215 61643 59247 61699
rect 59127 61601 59247 61643
rect 58647 59727 58649 59779
rect 58701 59727 58713 59779
rect 58765 59727 58767 59779
rect 58647 59687 58767 59727
rect 58887 60219 59007 60261
rect 58887 60163 58919 60219
rect 58975 60163 59007 60219
rect 58647 59608 58767 59648
rect 58647 59556 58649 59608
rect 58701 59556 58713 59608
rect 58765 59556 58767 59608
rect 58647 54299 58767 59556
rect 58887 58219 59007 60163
rect 58887 58163 58919 58219
rect 58975 58163 59007 58219
rect 58887 58121 59007 58163
rect 59127 58739 59247 58781
rect 59127 58683 59159 58739
rect 59215 58683 59247 58739
rect 59127 57859 59247 58683
rect 59127 57803 59159 57859
rect 59215 57803 59247 57859
rect 59127 57761 59247 57803
rect 58647 54243 58679 54299
rect 58735 54243 58767 54299
rect 58647 54201 58767 54243
rect 58407 52763 58439 52819
rect 58495 52763 58527 52819
rect 58407 52721 58527 52763
rect 59723 1700 59779 46402
rect 59723 1648 59725 1700
rect 59777 1648 59779 1700
rect 59723 1614 59779 1648
rect 60875 1500 60931 46402
rect 60875 1448 60877 1500
rect 60929 1448 60931 1500
rect 60875 1414 60931 1448
rect 62027 1300 62083 46402
rect 62027 1248 62029 1300
rect 62081 1248 62083 1300
rect 62027 1214 62083 1248
rect 63179 1100 63235 46402
rect 63179 1048 63181 1100
rect 63233 1048 63235 1100
rect 63179 1014 63235 1048
rect 64331 900 64387 46402
rect 64331 848 64333 900
rect 64385 848 64387 900
rect 64331 814 64387 848
rect 65483 700 65539 46402
rect 65483 648 65485 700
rect 65537 648 65539 700
rect 65483 614 65539 648
rect 66635 500 66691 46402
rect 66635 448 66637 500
rect 66689 448 66691 500
rect 66635 414 66691 448
rect 67787 300 67843 46402
rect 67787 248 67789 300
rect 67841 248 67843 300
rect 67787 214 67843 248
rect 68939 100 68995 46402
rect 68939 48 68941 100
rect 68993 48 68995 100
rect 68939 14 68995 48
rect 70091 -100 70147 46402
rect 70091 -152 70093 -100
rect 70145 -152 70147 -100
rect 70091 -186 70147 -152
rect 55829 -1002 55851 -950
rect 55903 -1002 55925 -950
rect 55829 -1014 55925 -1002
rect 55829 -1066 55851 -1014
rect 55903 -1066 55925 -1014
rect 55829 -1078 55925 -1066
rect 55829 -1130 55851 -1078
rect 55903 -1130 55925 -1078
rect 55829 -1142 55925 -1130
rect 55829 -1194 55851 -1142
rect 55903 -1194 55925 -1142
rect 55829 -1210 55925 -1194
rect 64079 -1463 64479 -1447
rect 64079 -1477 64093 -1463
rect 64465 -1477 64479 -1463
rect 64079 -1693 64091 -1477
rect 64467 -1693 64479 -1477
rect 64079 -1707 64093 -1693
rect 64465 -1707 64479 -1693
rect 64079 -1723 64479 -1707
<< via2 >>
rect 61091 121861 61093 122077
rect 61093 121861 61465 122077
rect 61465 121861 61467 122077
rect 67091 121861 67093 122077
rect 67093 121861 67465 122077
rect 67465 121861 67467 122077
rect -3880 121527 -3878 121565
rect -3878 121527 -3826 121565
rect -3826 121527 -3824 121565
rect -3880 121515 -3824 121527
rect -3880 121509 -3878 121515
rect -3878 121509 -3826 121515
rect -3826 121509 -3824 121515
rect -3880 121463 -3878 121485
rect -3878 121463 -3826 121485
rect -3826 121463 -3824 121485
rect -3880 121451 -3824 121463
rect -3880 121429 -3878 121451
rect -3878 121429 -3826 121451
rect -3826 121429 -3824 121451
rect -3880 121399 -3878 121405
rect -3878 121399 -3826 121405
rect -3826 121399 -3824 121405
rect -3880 121387 -3824 121399
rect -3880 121349 -3878 121387
rect -3878 121349 -3826 121387
rect -3826 121349 -3824 121387
rect 46779 120836 46789 121052
rect 46789 120836 46905 121052
rect 46905 120836 46915 121052
rect 46779 115083 46915 115219
rect 49265 72003 49321 72059
rect 49129 69043 49185 69099
rect 48929 67563 48985 67619
rect -3725 67455 -3669 67511
rect 48729 66083 48785 66139
rect 48529 64603 48585 64659
rect 48329 63123 48385 63179
rect 48129 62523 48185 62579
rect 650 61583 44466 61879
rect -3725 61429 -3669 61431
rect -3725 61377 -3723 61429
rect -3723 61377 -3671 61429
rect -3671 61377 -3669 61429
rect -3725 61375 -3669 61377
rect 58679 70523 58735 70579
rect -4546 60656 -4490 60658
rect -4546 60604 -4544 60656
rect -4544 60604 -4492 60656
rect -4492 60604 -4490 60656
rect -4546 60602 -4490 60604
rect -3276 60164 -3220 60220
rect -3881 59852 -3825 59854
rect -3881 59800 -3879 59852
rect -3879 59800 -3827 59852
rect -3827 59800 -3825 59852
rect -3881 59798 -3825 59800
rect -3725 59013 -3669 59015
rect -3725 58961 -3723 59013
rect -3723 58961 -3671 59013
rect -3671 58961 -3669 59013
rect -3725 58959 -3669 58961
rect -3725 52879 -3669 52935
rect 50369 60164 50425 60220
rect 650 58510 44466 58806
rect 47930 58163 47986 58219
rect 47730 57803 47786 57859
rect 47530 57203 47586 57259
rect 47330 55723 47386 55779
rect 50375 51283 50431 51339
rect 49266 48323 49322 48379
rect 49718 49803 49774 49859
rect -3437 43507 -3381 43563
rect 46499 5371 46635 5507
rect -3437 -328 -3381 -272
rect 46499 -668 46509 -452
rect 46509 -668 46625 -452
rect 46625 -668 46635 -452
rect 59159 62523 59215 62579
rect 59159 61643 59215 61699
rect 58919 60163 58975 60219
rect 58919 58163 58975 58219
rect 59159 58683 59215 58739
rect 59159 57803 59215 57859
rect 58679 54243 58735 54299
rect 58439 52763 58495 52819
rect 64091 -1693 64093 -1477
rect 64093 -1693 64465 -1477
rect 64465 -1693 64467 -1477
<< metal3 >>
rect 61069 122081 61489 122102
rect 61069 121857 61087 122081
rect 61471 121857 61489 122081
rect 61069 121836 61489 121857
rect 67069 122081 67489 122102
rect 67069 121857 67087 122081
rect 67471 121857 67489 122081
rect 67069 121836 67489 121857
rect -3911 121565 -3793 121590
rect -3911 121509 -3880 121565
rect -3824 121509 -3793 121565
rect -3911 121485 -3793 121509
rect -3911 121429 -3880 121485
rect -3824 121429 -3793 121485
rect -3911 121405 -3793 121429
rect -3911 121349 -3880 121405
rect -3824 121349 -3793 121405
rect -3911 121324 -3793 121349
rect -3901 64788 -3803 121324
rect 46767 121052 46927 121077
rect 46767 120836 46779 121052
rect 46915 120836 46927 121052
rect 46767 120811 46927 120836
rect 46777 115226 46917 120811
rect 46767 115219 46927 115226
rect 46767 115083 46779 115219
rect 46915 115083 46927 115219
rect 46767 115076 46927 115083
rect 70049 73155 70849 73275
rect 49251 72091 49335 72096
rect 49251 72059 59263 72091
rect 49251 72003 49265 72059
rect 49321 72003 59263 72059
rect 49251 71971 59263 72003
rect 49251 71966 49335 71971
rect 58637 70611 58777 70616
rect 58637 70579 59127 70611
rect 58637 70523 58679 70579
rect 58735 70523 59127 70579
rect 58637 70491 59127 70523
rect 58637 70486 58777 70491
rect 49087 69131 49227 69136
rect 49087 69099 59247 69131
rect 49087 69043 49129 69099
rect 49185 69043 59247 69099
rect 49087 69011 59247 69043
rect 49087 69006 49227 69011
rect 70049 68419 70849 68539
rect 48887 67651 49027 67656
rect 48887 67619 59267 67651
rect 48887 67563 48929 67619
rect 48985 67563 59267 67619
rect 48887 67531 59267 67563
rect 48887 67526 49027 67531
rect -3739 67511 -3655 67520
rect -3739 67455 -3725 67511
rect -3669 67455 -3655 67511
rect -3739 67446 -3655 67455
rect -10586 61041 -10320 62853
rect -3729 61440 -3665 67446
rect 48687 66171 48827 66176
rect 48687 66139 59247 66171
rect 48687 66083 48729 66139
rect 48785 66083 59247 66139
rect 48687 66051 59247 66083
rect 70049 66051 70849 66171
rect 48687 66046 48827 66051
rect 48487 64691 48627 64696
rect 48487 64659 59247 64691
rect 48487 64603 48529 64659
rect 48585 64603 59247 64659
rect 48487 64571 59247 64603
rect 48487 64566 48627 64571
rect 70049 63683 70849 63803
rect 48287 63211 48427 63216
rect 48287 63179 59247 63211
rect 48287 63123 48329 63179
rect 48385 63123 59247 63179
rect 48287 63091 59247 63123
rect 48287 63086 48427 63091
rect 48087 62611 48227 62616
rect 59117 62611 59257 62616
rect 48087 62579 59257 62611
rect 48087 62523 48129 62579
rect 48185 62523 59159 62579
rect 59215 62523 59257 62579
rect 48087 62491 59257 62523
rect 48087 62486 48227 62491
rect 59117 62486 59257 62491
rect 614 61883 44502 61905
rect 614 61579 646 61883
rect 44470 61579 44502 61883
rect 59117 61699 59257 61736
rect 59117 61643 59159 61699
rect 59215 61643 59257 61699
rect 59117 61606 59257 61643
rect 614 61558 44502 61579
rect -3739 61431 -3655 61440
rect -3739 61375 -3725 61431
rect -3669 61375 -3655 61431
rect -3739 61366 -3655 61375
rect 70049 61315 70849 61435
rect -4576 60658 -4460 60683
rect -4576 60602 -4546 60658
rect -4490 60602 -4460 60658
rect -4576 60577 -4460 60602
rect 58877 60251 59017 60256
rect -3290 60224 -3206 60229
rect 50355 60224 50439 60229
rect -3290 60220 50439 60224
rect -3290 60164 -3276 60220
rect -3220 60164 50369 60220
rect 50425 60164 50439 60220
rect -3290 60160 50439 60164
rect -3290 60155 -3206 60160
rect 50355 60155 50439 60160
rect 58877 60219 59127 60251
rect 58877 60163 58919 60219
rect 58975 60163 59127 60219
rect 58877 60131 59127 60163
rect 58877 60126 59017 60131
rect -3911 59854 -3795 59879
rect -3911 59798 -3881 59854
rect -3825 59798 -3795 59854
rect -3911 59773 -3795 59798
rect -10581 57547 -10325 59339
rect -3739 59015 -3655 59024
rect -3739 58959 -3725 59015
rect -3669 58959 -3655 59015
rect -3739 58950 -3655 58959
rect -3729 52944 -3665 58950
rect 70049 58947 70849 59067
rect 614 58810 44502 58832
rect 614 58506 646 58810
rect 44470 58506 44502 58810
rect 59117 58739 59257 58776
rect 59117 58683 59159 58739
rect 59215 58683 59257 58739
rect 59117 58646 59257 58683
rect 614 58485 44502 58506
rect 47888 58251 48028 58256
rect 58877 58251 59017 58256
rect 47888 58219 59017 58251
rect 47888 58163 47930 58219
rect 47986 58163 58919 58219
rect 58975 58163 59017 58219
rect 47888 58131 59017 58163
rect 47888 58126 48028 58131
rect 58877 58126 59017 58131
rect 47688 57891 47828 57896
rect 59117 57891 59257 57896
rect 47688 57859 59257 57891
rect 47688 57803 47730 57859
rect 47786 57803 59159 57859
rect 59215 57803 59257 57859
rect 47688 57771 59257 57803
rect 47688 57766 47828 57771
rect 59117 57766 59257 57771
rect 47488 57291 47628 57296
rect 47488 57259 59247 57291
rect 47488 57203 47530 57259
rect 47586 57203 59247 57259
rect 47488 57171 59247 57203
rect 47488 57166 47628 57171
rect 70049 56579 70849 56699
rect 47288 55811 47428 55816
rect 47288 55779 59248 55811
rect 47288 55723 47330 55779
rect 47386 55723 59248 55779
rect 47288 55691 59248 55723
rect 47288 55686 47428 55691
rect 58637 54331 58777 54336
rect 58637 54299 59127 54331
rect 58637 54243 58679 54299
rect 58735 54243 59127 54299
rect 58637 54211 59127 54243
rect 70049 54211 70849 54331
rect 58637 54206 58777 54211
rect -3739 52935 -3655 52944
rect -3739 52879 -3725 52935
rect -3669 52879 -3655 52935
rect -3739 52870 -3655 52879
rect 58397 52851 58537 52856
rect 58397 52819 59127 52851
rect 58397 52763 58439 52819
rect 58495 52763 59127 52819
rect 58397 52731 59127 52763
rect 58397 52726 58537 52731
rect 70049 51843 70849 51963
rect 50365 51371 50441 51376
rect 50365 51339 59288 51371
rect 50365 51283 50375 51339
rect 50431 51283 59288 51339
rect 50365 51251 59288 51283
rect 50365 51246 50441 51251
rect 49676 49891 49816 49896
rect 49676 49859 59279 49891
rect 49676 49803 49718 49859
rect 49774 49803 59279 49859
rect 49676 49771 59279 49803
rect 49676 49766 49816 49771
rect 70049 49475 70849 49595
rect 49252 48411 49336 48416
rect 49252 48379 59391 48411
rect 49252 48323 49266 48379
rect 49322 48323 59391 48379
rect 49252 48291 59391 48323
rect 49252 48286 49336 48291
rect 70049 47107 70849 47227
rect -3479 43563 -3339 43600
rect -3479 43507 -3437 43563
rect -3381 43507 -3339 43563
rect -3479 43470 -3339 43507
rect -3469 -235 -3349 43470
rect 46487 5507 46648 5515
rect 46487 5371 46499 5507
rect 46635 5371 46648 5507
rect 46487 5364 46648 5371
rect -3479 -272 -3339 -235
rect -3479 -328 -3437 -272
rect -3381 -328 -3339 -272
rect -3479 -365 -3339 -328
rect 46497 -427 46638 5364
rect 46487 -452 46648 -427
rect 46487 -668 46499 -452
rect 46635 -668 46648 -452
rect 46487 -693 46648 -668
rect 64069 -1473 64489 -1452
rect 64069 -1697 64087 -1473
rect 64471 -1697 64489 -1473
rect 64069 -1718 64489 -1697
<< via3 >>
rect 61087 122077 61471 122081
rect 61087 121861 61091 122077
rect 61091 121861 61467 122077
rect 61467 121861 61471 122077
rect 61087 121857 61471 121861
rect 67087 122077 67471 122081
rect 67087 121861 67091 122077
rect 67091 121861 67467 122077
rect 67467 121861 67471 122077
rect 67087 121857 67471 121861
rect 646 61879 44470 61883
rect 646 61583 650 61879
rect 650 61583 44466 61879
rect 44466 61583 44470 61879
rect 646 61579 44470 61583
rect 646 58806 44470 58810
rect 646 58510 650 58806
rect 650 58510 44466 58806
rect 44466 58510 44470 58806
rect 646 58506 44470 58510
rect 64087 -1477 64471 -1473
rect 64087 -1693 64091 -1477
rect 64091 -1693 64467 -1477
rect 64467 -1693 64471 -1477
rect 64087 -1697 64471 -1693
<< metal4 >>
rect 61078 122081 61480 122098
rect 61078 121857 61087 122081
rect 61471 121857 61480 122081
rect 61078 121840 61480 121857
rect 67078 122081 67480 122098
rect 67078 121857 67087 122081
rect 67471 121857 67480 122081
rect 67078 121840 67480 121857
rect 61079 71451 61479 121840
rect 67079 71328 67479 121840
rect 623 61883 44493 61901
rect 623 61579 646 61883
rect 44470 61579 44493 61883
rect 623 61562 44493 61579
rect 623 58810 44493 58828
rect 623 58506 646 58810
rect 44470 58506 44493 58810
rect 623 58489 44493 58506
rect 64079 -1456 64479 49005
rect 64078 -1473 64480 -1456
rect 64078 -1697 64087 -1473
rect 64471 -1697 64480 -1473
rect 64078 -1714 64480 -1697
use cdac  cdac_0
timestamp 1750100919
transform 1 0 -1274 0 1 2329
box -1099 -705 50472 116437
use sar10b  sar10b_0
timestamp 1750100919
transform 1 0 59127 0 1 45909
box 0 0 11722 28874
use tdc  tdc_0
timestamp 1750100919
transform 1 0 50703 0 1 59011
box -224 -646 5424 3006
use th_dif_sw  th_dif_sw_0
timestamp 1750100919
transform 0 -1 -4206 1 0 44365
box -1 -413 31660 6385
<< labels >>
flabel metal1 s -10590 43715 -10470 43835 0 FreeSans 1000 0 0 0 VCM
port 1 nsew
flabel metal1 s -10590 43475 -10470 43595 0 FreeSans 1000 0 0 0 EN
port 2 nsew
flabel metal1 s -11103 121329 -10847 121585 0 FreeSans 1000 0 0 0 VDDA
port 3 nsew
flabel metal1 s -11103 120816 -10847 121072 0 FreeSans 1000 0 0 0 VDDR
port 4 nsew
flabel metal1 s -10590 43955 -10470 44075 0 FreeSans 1000 0 0 0 CLK
port 5 nsew
flabel metal3 s 70729 73155 70849 73275 0 FreeSans 1000 0 0 0 CKO
port 6 nsew
flabel metal3 s -10485 61786 -10455 61816 0 FreeSans 1000 0 0 0 VINP
port 7 nsew
flabel metal3 s 70729 66051 70849 66171 0 FreeSans 1000 0 0 0 DATA[8]
port 8 nsew
flabel metal3 s 70729 63683 70849 63803 0 FreeSans 1000 0 0 0 DATA[7]
port 9 nsew
flabel metal3 s 70729 61315 70849 61435 0 FreeSans 1000 0 0 0 DATA[6]
port 10 nsew
flabel metal3 s 70729 58947 70849 59067 0 FreeSans 1000 0 0 0 DATA[5]
port 11 nsew
flabel metal3 s 70729 56579 70849 56699 0 FreeSans 1000 0 0 0 DATA[4]
port 12 nsew
flabel metal3 s 70729 54211 70849 54331 0 FreeSans 1000 0 0 0 DATA[3]
port 13 nsew
flabel metal3 s 70729 51843 70849 51963 0 FreeSans 1000 0 0 0 DATA[2]
port 14 nsew
flabel metal3 s 70729 49475 70849 49595 0 FreeSans 1000 0 0 0 DATA[1]
port 15 nsew
flabel metal3 s 70729 47107 70849 47227 0 FreeSans 1000 0 0 0 DATA[0]
port 16 nsew
flabel metal1 s -11102 -688 -10846 -432 0 FreeSans 500 0 0 0 VSSR
port 17 nsew
flabel metal1 s -11102 -1200 -10846 -944 0 FreeSans 500 0 0 0 VSSA
port 18 nsew
flabel metal1 s -11102 -1713 -10846 -1457 0 FreeSans 500 0 0 0 VSSD
port 19 nsew
flabel metal1 s -11039 121933 -10943 122029 0 FreeSans 500 0 0 0 VDDD
port 20 nsew
flabel metal3 s 70777 68452 70822 68500 0 FreeSans 500 0 0 0 DATA[9]
port 21 nsew
flabel metal3 s -10479 58608 -10449 58638 0 FreeSans 1000 0 0 0 VINN
port 22 nsew
<< end >>
