magic
tech sky130A
magscale 1 2
timestamp 1749226129
<< pwell >>
rect 42 -49 1464 212
<< viali >>
rect 1393 325 1433 365
rect 77 208 117 248
rect 239 201 299 261
rect 353 201 413 261
rect 535 208 575 248
rect 805 214 865 274
rect 967 230 1027 290
rect 241 113 281 153
rect 529 34 569 74
<< metal1 >>
rect 38 568 1478 666
rect 0 451 353 511
rect 413 451 805 511
rect 865 451 875 511
rect 0 331 239 391
rect 299 331 967 391
rect 1027 331 1037 391
rect 1381 365 1445 371
rect 1381 325 1393 365
rect 1433 325 1516 365
rect 1381 319 1445 325
rect 955 290 1039 296
rect 793 274 877 280
rect 227 261 311 267
rect 65 248 129 254
rect 65 208 77 248
rect 117 208 129 248
rect 65 202 129 208
rect 77 74 117 202
rect 227 201 239 261
rect 299 201 311 261
rect 227 195 311 201
rect 341 261 425 267
rect 341 201 353 261
rect 413 201 425 261
rect 523 248 587 254
rect 523 208 535 248
rect 575 208 587 248
rect 793 214 805 274
rect 865 214 877 274
rect 955 230 967 290
rect 1027 230 1039 290
rect 955 224 1039 230
rect 793 208 877 214
rect 523 202 587 208
rect 341 195 425 201
rect 229 153 293 159
rect 535 153 575 202
rect 229 113 241 153
rect 281 113 1516 153
rect 229 107 293 113
rect 517 74 581 80
rect 77 34 529 74
rect 569 34 1516 74
rect 517 28 581 34
rect 38 -98 1478 0
<< via1 >>
rect 353 451 413 511
rect 805 451 865 511
rect 239 331 299 391
rect 967 331 1027 391
rect 239 201 299 261
rect 353 201 413 261
rect 805 214 865 274
rect 967 230 1027 290
<< metal2 >>
rect 353 511 413 521
rect 239 391 299 401
rect 239 261 299 331
rect 239 191 299 201
rect 353 261 413 451
rect 805 511 865 521
rect 805 274 865 451
rect 967 391 1027 401
rect 967 290 1027 331
rect 967 220 1027 230
rect 805 204 865 214
rect 353 191 413 201
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749010377
transform 1 0 614 0 1 -49
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749010377
transform 1 0 38 0 1 -49
box -38 -49 326 715
use sky130_fd_sc_hs__nand2_1  x2
timestamp 1749010377
transform 1 0 326 0 1 -49
box -38 -49 326 715
use sky130_fd_sc_hs__xor2_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 710 0 1 -49
box -38 -49 806 715
<< labels >>
flabel metal1 0 451 30 511 0 FreeSans 400 0 0 0 A
port 0 nsew
flabel metal1 0 331 30 391 0 FreeSans 400 0 0 0 B
port 1 nsew
flabel metal1 91 568 189 666 0 FreeSans 400 0 0 0 VDD
port 2 nsew
flabel metal1 95 -98 193 0 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 1496 325 1516 365 0 FreeSans 400 0 0 0 RDY
port 4 nsew
flabel metal1 1476 113 1516 153 0 FreeSans 400 0 0 0 OUTP
port 5 nsew
flabel metal1 1476 34 1516 74 0 FreeSans 400 0 0 0 OUTN
port 7 nsew
<< end >>
