* NGSPICE file created from sar10b.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

.subckt sar10b CF[0] CF[1] CF[2] CF[3] CF[4] CF[5] CF[6] CF[7] CF[8] CF[9] CKO CKS
+ CKSB CLK CMP_N CMP_P DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7]
+ DATA[8] DATA[9] EN RDY SWN[0] SWN[1] SWN[2] SWN[3] SWN[4] SWN[5] SWN[6] SWN[7] SWN[8]
+ SWN[9] SWP[0] SWP[1] SWP[2] SWP[3] SWP[4] SWP[5] SWP[6] SWP[7] SWP[8] SWP[9] VGND
+ VPWR
X_83_ cyclic_flag_0.FINAL net40 net3 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_66_ net14 net1 net16 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_49_ net4 net12 net16 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput7 net7 VGND VGND VPWR VPWR CF[2] sky130_fd_sc_hd__buf_1
Xoutput42 net42 VGND VGND VPWR VPWR SWP[4] sky130_fd_sc_hd__buf_1
Xoutput20 net20 VGND VGND VPWR VPWR DATA[2] sky130_fd_sc_hd__buf_1
Xoutput31 net31 VGND VGND VPWR VPWR SWN[3] sky130_fd_sc_hd__buf_1
XFILLER_0_1_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_82_ cyclic_flag_0.FINAL net41 net3 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfrtp_1
X_65_ net5 net2 net16 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_48_ net4 net11 net16 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput10 net10 VGND VGND VPWR VPWR CF[5] sky130_fd_sc_hd__buf_1
Xoutput8 net8 VGND VGND VPWR VPWR CF[3] sky130_fd_sc_hd__buf_1
Xoutput43 net43 VGND VGND VPWR VPWR SWP[5] sky130_fd_sc_hd__buf_1
Xoutput32 net32 VGND VGND VPWR VPWR SWN[4] sky130_fd_sc_hd__buf_1
Xoutput21 net21 VGND VGND VPWR VPWR DATA[3] sky130_fd_sc_hd__buf_1
X_81_ cyclic_flag_0.FINAL net42 net3 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_19_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_64_ net6 net2 net16 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_4_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_47_ net4 net10 net16 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput9 net9 VGND VGND VPWR VPWR CF[4] sky130_fd_sc_hd__buf_1
Xoutput11 net11 VGND VGND VPWR VPWR CF[6] sky130_fd_sc_hd__buf_1
Xoutput44 net44 VGND VGND VPWR VPWR SWP[6] sky130_fd_sc_hd__buf_1
Xoutput33 net33 VGND VGND VPWR VPWR SWN[5] sky130_fd_sc_hd__buf_1
Xoutput22 net22 VGND VGND VPWR VPWR DATA[4] sky130_fd_sc_hd__buf_1
XFILLER_0_11_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_80_ cyclic_flag_0.FINAL net43 net3 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_63_ net7 net2 net16 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_20_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_46_ net4 net9 net16 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_29_ clk_div_0.COUNT\[1\] clk_div_0.COUNT\[0\] _11_ VGND VGND VPWR VPWR _03_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput12 net12 VGND VGND VPWR VPWR CF[7] sky130_fd_sc_hd__buf_1
Xoutput45 net45 VGND VGND VPWR VPWR SWP[7] sky130_fd_sc_hd__buf_1
Xoutput34 net34 VGND VGND VPWR VPWR SWN[6] sky130_fd_sc_hd__buf_1
Xoutput23 net23 VGND VGND VPWR VPWR DATA[5] sky130_fd_sc_hd__buf_1
XFILLER_0_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_62_ net8 net2 net16 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_45_ net4 net8 net16 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfrtp_1
Xclkload0 clknet_1_0__leaf_CLK VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_28_ clk_div_0.COUNT\[1\] clk_div_0.COUNT\[0\] net3 VGND VGND VPWR VPWR _11_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput13 net13 VGND VGND VPWR VPWR CF[8] sky130_fd_sc_hd__buf_1
Xoutput46 net46 VGND VGND VPWR VPWR SWP[8] sky130_fd_sc_hd__buf_1
Xoutput35 net35 VGND VGND VPWR VPWR SWN[7] sky130_fd_sc_hd__buf_1
Xoutput24 net24 VGND VGND VPWR VPWR DATA[6] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_21_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_61_ net9 net2 net16 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_1__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_1_1__leaf_CLK sky130_fd_sc_hd__clkbuf_16
X_44_ net4 net7 net16 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_27_ clk_div_0.COUNT\[0\] _08_ VGND VGND VPWR VPWR _02_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput14 net14 VGND VGND VPWR VPWR CF[9] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_21_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput47 net47 VGND VGND VPWR VPWR SWP[9] sky130_fd_sc_hd__buf_1
Xoutput36 net36 VGND VGND VPWR VPWR SWN[8] sky130_fd_sc_hd__buf_1
Xoutput25 net25 VGND VGND VPWR VPWR DATA[7] sky130_fd_sc_hd__buf_1
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_60_ net10 net2 net16 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_43_ net4 net6 net16 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_26_ net16 _10_ _09_ VGND VGND VPWR VPWR _01_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_11_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net15 VGND VGND VPWR VPWR CKO sky130_fd_sc_hd__buf_1
Xoutput37 net37 VGND VGND VPWR VPWR SWN[9] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput26 net26 VGND VGND VPWR VPWR DATA[8] sky130_fd_sc_hd__buf_1
XFILLER_0_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_42_ net4 net5 net16 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25_ net3 _07_ VGND VGND VPWR VPWR _10_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput38 net38 VGND VGND VPWR VPWR SWP[0] sky130_fd_sc_hd__buf_1
Xoutput27 net27 VGND VGND VPWR VPWR DATA[9] sky130_fd_sc_hd__buf_1
Xoutput16 net16 VGND VGND VPWR VPWR CKS sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_41_ net4 net16 net16 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24_ net17 _08_ _09_ VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput39 net39 VGND VGND VPWR VPWR SWP[1] sky130_fd_sc_hd__buf_1
Xoutput28 net28 VGND VGND VPWR VPWR SWN[0] sky130_fd_sc_hd__buf_1
Xoutput17 net17 VGND VGND VPWR VPWR CKSB sky130_fd_sc_hd__buf_1
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_40_ clknet_1_1__leaf_CLK _01_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfxtp_4
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_23_ _07_ net16 net3 VGND VGND VPWR VPWR _09_ sky130_fd_sc_hd__or3b_1
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput18 net18 VGND VGND VPWR VPWR DATA[0] sky130_fd_sc_hd__buf_1
Xoutput29 net29 VGND VGND VPWR VPWR SWN[1] sky130_fd_sc_hd__buf_1
XFILLER_0_7_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_15_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22_ net3 _07_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_19_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput19 net19 VGND VGND VPWR VPWR DATA[1] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21_ clk_div_0.COUNT\[1\] clk_div_0.COUNT\[0\] clk_div_0.COUNT\[2\] clk_div_0.COUNT\[3\]
+ VGND VGND VPWR VPWR _07_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20_ _06_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 CMP_N VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 CMP_P VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
X_79_ cyclic_flag_0.FINAL net44 net3 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_21_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput3 EN VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_4
XFILLER_0_11_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_78_ cyclic_flag_0.FINAL net45 net3 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_77_ cyclic_flag_0.FINAL net46 net3 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfrtp_1
Xinput4 RDY VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_76_ cyclic_flag_0.FINAL net47 net3 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_59_ net11 net2 net16 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_75_ net5 net1 net16 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_58_ net12 net2 net16 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_74_ net6 net1 net16 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_2_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_57_ net13 net2 net16 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_73_ net7 net1 net16 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_56_ net14 net2 net16 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_39_ clknet_1_1__leaf_CLK _00_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_72_ net8 net1 net16 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_55_ clknet_1_0__leaf_CLK _05_ VGND VGND VPWR VPWR clk_div_0.COUNT\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_38_ _18_ VGND VGND VPWR VPWR _05_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_71_ net9 net1 net16 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_54_ clknet_1_0__leaf_CLK _04_ VGND VGND VPWR VPWR clk_div_0.COUNT\[2\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_6_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_37_ _10_ _16_ _17_ VGND VGND VPWR VPWR _18_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_70_ net10 net1 net16 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_53_ clknet_1_0__leaf_CLK _03_ VGND VGND VPWR VPWR clk_div_0.COUNT\[1\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0_CLK CLK VGND VGND VPWR VPWR clknet_0_CLK sky130_fd_sc_hd__clkbuf_16
X_36_ _15_ _12_ VGND VGND VPWR VPWR _17_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19_ net16 cyclic_flag_0.FINAL VGND VGND VPWR VPWR _06_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_4_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_52_ clknet_1_1__leaf_CLK _02_ VGND VGND VPWR VPWR clk_div_0.COUNT\[0\] sky130_fd_sc_hd__dfxtp_1
X_35_ _15_ _12_ VGND VGND VPWR VPWR _16_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_51_ net4 net14 net16 VGND VGND VPWR VPWR cyclic_flag_0.FINAL sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_34_ clk_div_0.COUNT\[3\] VGND VGND VPWR VPWR _15_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_50_ net4 net13 net16 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_33_ _14_ VGND VGND VPWR VPWR _04_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32_ _10_ _12_ _13_ VGND VGND VPWR VPWR _14_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_31_ clk_div_0.COUNT\[1\] clk_div_0.COUNT\[0\] clk_div_0.COUNT\[2\] VGND VGND VPWR
+ VPWR _13_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_30_ clk_div_0.COUNT\[1\] clk_div_0.COUNT\[0\] clk_div_0.COUNT\[2\] VGND VGND VPWR
+ VPWR _12_ sky130_fd_sc_hd__nand3_1
XFILLER_0_20_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_45 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_69_ net11 net1 net16 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_85_ cyclic_flag_0.FINAL net38 net3 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_68_ net12 net1 net16 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_12_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput5 net5 VGND VGND VPWR VPWR CF[0] sky130_fd_sc_hd__buf_1
Xoutput40 net40 VGND VGND VPWR VPWR SWP[2] sky130_fd_sc_hd__buf_1
XFILLER_0_5_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_1_0__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_84_ cyclic_flag_0.FINAL net39 net3 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_0_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_67_ net13 net1 net16 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput6 net6 VGND VGND VPWR VPWR CF[1] sky130_fd_sc_hd__buf_1
Xoutput41 net41 VGND VGND VPWR VPWR SWP[3] sky130_fd_sc_hd__buf_1
Xoutput30 net30 VGND VGND VPWR VPWR SWN[2] sky130_fd_sc_hd__buf_1
.ends

