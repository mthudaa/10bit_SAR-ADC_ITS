magic
tech sky130A
magscale 1 2
timestamp 1748792115
<< viali >>
rect 142 1527 6372 1561
rect 142 -123 3320 -89
<< metal1 >>
rect 106 1561 6408 1597
rect 106 1527 142 1561
rect 6372 1527 6408 1561
rect 106 1521 6408 1527
rect 325 1447 6189 1521
rect 106 1301 176 1401
rect 228 1301 284 1401
rect 325 1061 6189 1255
rect 106 915 284 1015
rect 106 569 6408 869
rect 106 423 284 523
rect 316 183 3146 377
rect 166 37 176 137
rect 228 37 284 137
rect 316 -83 3146 -9
rect 106 -89 6408 -83
rect 106 -123 142 -89
rect 3320 -123 6408 -89
rect 106 -159 6408 -123
<< via1 >>
rect 176 1301 228 1401
rect 176 37 228 137
<< metal2 >>
rect 176 1401 228 1411
rect 176 137 228 1301
rect 176 27 228 37
use sky130_fd_pr__nfet_01v8_H9ZN2D  sky130_fd_pr__nfet_01v8_H9ZN2D_0
timestamp 1746380519
transform 0 1 1731 -1 0 87
box -246 -1625 246 1625
use sky130_fd_pr__pfet_01v8_D9Q956  sky130_fd_pr__pfet_01v8_D9Q956_0
timestamp 1746380519
transform 0 1 3257 -1 0 965
box -246 -3151 246 3151
use sky130_fd_pr__pfet_01v8_D9Q956  XM1
timestamp 1746380519
transform 0 1 3257 -1 0 1351
box -246 -3151 246 3151
use sky130_fd_pr__nfet_01v8_H9ZN2D  XM3
timestamp 1746380519
transform 0 1 1731 -1 0 473
box -246 -1625 246 1625
<< labels >>
flabel metal1 113 1556 120 1563 0 FreeSans 400 0 0 0 VDD
port 0 nsew
flabel metal1 119 1345 126 1352 0 FreeSans 400 0 0 0 IN
port 1 nsew
flabel metal1 119 960 126 967 0 FreeSans 400 0 0 0 CKB
port 2 nsew
flabel metal1 119 469 126 476 0 FreeSans 400 0 0 0 CK
port 3 nsew
flabel metal1 122 -125 129 -118 0 FreeSans 400 0 0 0 VSS
port 4 nsew
flabel metal1 6347 690 6354 697 0 FreeSans 400 0 0 0 OUT
port 6 nsew
<< end >>
