* NGSPICE file created from sar10b.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hs__dfrtp_1 abstract view
.subckt sky130_fd_sc_hs__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hs__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__fill_1 abstract view
.subckt sky130_fd_sc_hs__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__fill_8 abstract view
.subckt sky130_fd_sc_hs__fill_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__decap_4 abstract view
.subckt sky130_fd_sc_hs__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__dfrtp_2 abstract view
.subckt sky130_fd_sc_hs__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__fill_2 abstract view
.subckt sky130_fd_sc_hs__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__and2_1 abstract view
.subckt sky130_fd_sc_hs__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__xor2_1 abstract view
.subckt sky130_fd_sc_hs__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__clkbuf_16 abstract view
.subckt sky130_fd_sc_hs__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nor2_1 abstract view
.subckt sky130_fd_sc_hs__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__clkbuf_1 abstract view
.subckt sky130_fd_sc_hs__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__a21bo_1 abstract view
.subckt sky130_fd_sc_hs__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__o21a_1 abstract view
.subckt sky130_fd_sc_hs__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__or3b_1 abstract view
.subckt sky130_fd_sc_hs__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nand2_1 abstract view
.subckt sky130_fd_sc_hs__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__or4bb_1 abstract view
.subckt sky130_fd_sc_hs__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__clkbuf_2 abstract view
.subckt sky130_fd_sc_hs__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__buf_8 abstract view
.subckt sky130_fd_sc_hs__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__clkbuf_4 abstract view
.subckt sky130_fd_sc_hs__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__dfxtp_4 abstract view
.subckt sky130_fd_sc_hs__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__dfxtp_1 abstract view
.subckt sky130_fd_sc_hs__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__nor3_1 abstract view
.subckt sky130_fd_sc_hs__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__a21oi_1 abstract view
.subckt sky130_fd_sc_hs__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hs__and3_1 abstract view
.subckt sky130_fd_sc_hs__and3_1 A B C VGND VNB VPB VPWR X
.ends

.subckt sar10b CF[0] CF[1] CF[2] CF[3] CF[4] CF[5] CF[6] CF[7] CF[8] CF[9] CKO CKS
+ CKSB CLK CMP_N CMP_P DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7]
+ DATA[8] DATA[9] EN RDY SWN[0] SWN[1] SWN[2] SWN[3] SWN[4] SWN[5] SWN[6] SWN[7] SWN[8]
+ SWN[9] SWP[0] SWP[1] SWP[2] SWP[3] SWP[4] SWP[5] SWP[6] SWP[7] SWP[8] SWP[9] VGND
+ VPWR
X_83_ cyclic_flag_0.FINAL SWP[0] net3 VGND VGND VPWR VPWR DATA[0] sky130_fd_sc_hs__dfrtp_1
XTAP_TAPCELL_ROW_12_76 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_18_18 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XTAP_TAPCELL_ROW_8_66 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_66_ CF[7] net1 CKS VGND VGND VPWR VPWR SWN[7] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_4_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_19_61 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_49_ net4 CF[9] CKS VGND VGND VPWR VPWR cyclic_flag_0.FINAL sky130_fd_sc_hs__dfrtp_2
XTAP_TAPCELL_ROW_20_98 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_6_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_4_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_82_ cyclic_flag_0.FINAL SWP[1] net3 VGND VGND VPWR VPWR DATA[1] sky130_fd_sc_hs__dfrtp_1
XTAP_TAPCELL_ROW_12_77 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_67 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_65_ CF[8] net1 CKS VGND VGND VPWR VPWR SWN[8] sky130_fd_sc_hs__dfrtp_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_48_ net4 CF[8] CKS VGND VGND VPWR VPWR CF[9] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_10_42 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_21_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_1_95 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_16_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_12_110 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_81_ cyclic_flag_0.FINAL SWP[2] net3 VGND VGND VPWR VPWR DATA[2] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_13_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_19_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_12_78 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_64_ CF[9] net1 CKS VGND VGND VPWR VPWR SWN[9] sky130_fd_sc_hs__dfrtp_1
XTAP_TAPCELL_ROW_8_68 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_47_ net4 CF[7] CKS VGND VGND VPWR VPWR CF[8] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_21_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_1_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_21_144 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_7_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_80_ cyclic_flag_0.FINAL SWP[3] net3 VGND VGND VPWR VPWR DATA[3] sky130_fd_sc_hs__dfrtp_1
XPHY_EDGE_ROW_20_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_4_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_63_ CF[0] net2 CKS VGND VGND VPWR VPWR SWP[0] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_46_ net4 CF[6] CKS VGND VGND VPWR VPWR CF[7] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_19_117 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_18_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XTAP_TAPCELL_ROW_5_59 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_29_ net3 _12_ VGND VGND VPWR VPWR _13_ sky130_fd_sc_hs__and2_1
XFILLER_0_16_98 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_9_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_11_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_62_ CF[1] net2 CKS VGND VGND VPWR VPWR SWP[1] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_45_ net4 CF[5] CKS VGND VGND VPWR VPWR CF[6] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_1_87 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_28_ clk_div_0.COUNT\[1\] clk_div_0.COUNT\[0\] VGND VGND VPWR VPWR _12_ sky130_fd_sc_hs__xor2_1
XFILLER_0_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_22 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_13_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_61_ CF[2] net2 CKS VGND VGND VPWR VPWR SWP[2] sky130_fd_sc_hs__dfrtp_1
Xclkbuf_1_1__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_1_1__leaf_CLK sky130_fd_sc_hs__clkbuf_16
XFILLER_0_19_22 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_13_80 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_44_ net4 CF[4] CKS VGND VGND VPWR VPWR CF[5] sky130_fd_sc_hs__dfrtp_1
XTAP_TAPCELL_ROW_9_70 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_21_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_27_ clk_div_0.COUNT\[0\] _08_ VGND VGND VPWR VPWR _02_ sky130_fd_sc_hs__nor2_1
XFILLER_0_21_136 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_16_45 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_16_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_7_10 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_60_ CF[3] net2 CKS VGND VGND VPWR VPWR SWP[3] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_10_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_43_ net4 CF[3] CKS VGND VGND VPWR VPWR CF[4] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_26_ _11_ VGND VGND VPWR VPWR _01_ sky130_fd_sc_hs__clkbuf_1
XFILLER_0_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_10_71 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_18_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_6_61 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_12_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_4_134 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_4_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_42_ net4 CF[2] CKS VGND VGND VPWR VPWR CF[3] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_25_ CKS _10_ _09_ VGND VGND VPWR VPWR _11_ sky130_fd_sc_hs__a21bo_1
XFILLER_0_1_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_10_72 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_16_69 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_6_62 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_41_ net4 CF[1] CKS VGND VGND VPWR VPWR CF[2] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_21_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_24_ net3 _07_ VGND VGND VPWR VPWR _10_ sky130_fd_sc_hs__and2_1
XFILLER_0_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_21_117 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_10_73 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XTAP_TAPCELL_ROW_6_63 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_12_106 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_1_139 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_40_ net4 CF[0] CKS VGND VGND VPWR VPWR CF[1] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_10_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_23_ CKSB _08_ _09_ VGND VGND VPWR VPWR _00_ sky130_fd_sc_hs__o21a_1
XTAP_TAPCELL_ROW_19_94 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_15_104 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_11_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_4_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_7_14 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_15_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_3_54 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_1_107 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_13_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_5_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_18_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_0_44 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_22_ _07_ CKS net3 VGND VGND VPWR VPWR _09_ sky130_fd_sc_hs__or3b_1
XTAP_TAPCELL_ROW_19_95 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_7_102 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_4_116 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_3_55 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_0_45 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_21_ net3 _07_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hs__nand2_1
XFILLER_0_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_21_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_14_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_7_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XTAP_TAPCELL_ROW_16_86 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_3_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_21_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_4_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_0_46 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_5_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_20_ clk_div_0.COUNT\[1\] clk_div_0.COUNT\[0\] clk_div_0.COUNT\[2\] clk_div_0.COUNT\[3\]
+ VGND VGND VPWR VPWR _07_ sky130_fd_sc_hs__or4bb_1
XFILLER_0_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_11_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
Xinput1 CMP_N VGND VGND VPWR VPWR net1 sky130_fd_sc_hs__clkbuf_2
XFILLER_0_20_143 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_17_95 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_16_87 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_14_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_0_47 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_15_119 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_7_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_79_ cyclic_flag_0.FINAL SWP[4] net3 VGND VGND VPWR VPWR DATA[4] sky130_fd_sc_hs__dfrtp_1
Xinput2 CMP_P VGND VGND VPWR VPWR net2 sky130_fd_sc_hs__clkbuf_2
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_21_99 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_17_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_16_88 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_8_94 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_0_48 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
Xinput3 EN VGND VGND VPWR VPWR net3 sky130_fd_sc_hs__buf_8
XFILLER_0_11_32 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_11_87 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_78_ cyclic_flag_0.FINAL SWP[5] net3 VGND VGND VPWR VPWR DATA[5] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_2_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_6_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_3_142 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_10_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_13_79 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_69 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
Xinput4 RDY VGND VGND VPWR VPWR net4 sky130_fd_sc_hs__clkbuf_4
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_77_ cyclic_flag_0.FINAL SWP[6] net3 VGND VGND VPWR VPWR DATA[6] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_2_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_8_96 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_12_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_1_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_76_ cyclic_flag_0.FINAL SWP[7] net3 VGND VGND VPWR VPWR DATA[7] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_59_ CF[4] net2 CKS VGND VGND VPWR VPWR SWP[4] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_3_100 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_14_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_17_90 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_1_50 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_75_ cyclic_flag_0.FINAL SWP[8] net3 VGND VGND VPWR VPWR DATA[8] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_9_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_58_ CF[5] net2 CKS VGND VGND VPWR VPWR SWP[5] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_17_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_14_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_14_81 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_74_ cyclic_flag_0.FINAL SWP[9] net3 VGND VGND VPWR VPWR DATA[9] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_20_127 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_2_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_2_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_12_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_57_ CF[6] net2 CKS VGND VGND VPWR VPWR SWP[6] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_17_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_14_82 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_73_ CF[0] net1 CKS VGND VGND VPWR VPWR SWN[0] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_14_125 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_56_ CF[7] net2 CKS VGND VGND VPWR VPWR SWP[7] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
X_39_ net4 CKS CKS VGND VGND VPWR VPWR CF[0] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_8_34 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_5_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_14_83 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_72_ CF[1] net1 CKS VGND VGND VPWR VPWR SWN[1] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_11_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_55_ CF[8] net2 CKS VGND VGND VPWR VPWR SWP[8] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_38_ clknet_1_1__leaf_CLK _01_ VGND VGND VPWR VPWR CKS sky130_fd_sc_hs__dfxtp_4
XFILLER_0_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_71_ CF[2] net1 CKS VGND VGND VPWR VPWR SWN[2] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_54_ CF[9] net2 CKS VGND VGND VPWR VPWR SWP[9] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_6_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_11_74 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XTAP_TAPCELL_ROW_7_64 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_37_ clknet_1_1__leaf_CLK _00_ VGND VGND VPWR VPWR CKSB sky130_fd_sc_hs__dfxtp_1
XPHY_EDGE_ROW_9_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_15_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_70_ CF[3] net1 CKS VGND VGND VPWR VPWR SWN[3] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_13_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
Xclkbuf_0_CLK CLK VGND VGND VPWR VPWR clknet_0_CLK sky130_fd_sc_hs__clkbuf_16
X_53_ clknet_1_1__leaf_CLK _05_ VGND VGND VPWR VPWR clk_div_0.COUNT\[3\] sky130_fd_sc_hs__dfxtp_1
XFILLER_0_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_11_75 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_12_72 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_7_65 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
X_36_ _17_ VGND VGND VPWR VPWR _05_ sky130_fd_sc_hs__clkbuf_1
XFILLER_0_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_19_ _06_ VGND VGND VPWR VPWR CKO sky130_fd_sc_hs__clkbuf_1
XFILLER_0_19_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_20_72 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_2_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_52_ clknet_1_0__leaf_CLK _04_ VGND VGND VPWR VPWR clk_div_0.COUNT\[2\] sky130_fd_sc_hs__dfxtp_1
XFILLER_0_6_115 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_6_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_35_ _10_ _16_ VGND VGND VPWR VPWR _17_ sky130_fd_sc_hs__and2_1
X_18_ CKS cyclic_flag_0.FINAL VGND VGND VPWR VPWR _06_ sky130_fd_sc_hs__and2_1
XFILLER_0_18_50 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_4_56 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_20_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_51_ clknet_1_0__leaf_CLK _03_ VGND VGND VPWR VPWR clk_div_0.COUNT\[1\] sky130_fd_sc_hs__dfxtp_1
X_34_ clk_div_0.COUNT\[3\] _14_ VGND VGND VPWR VPWR _16_ sky130_fd_sc_hs__xor2_1
XFILLER_0_8_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_4_57 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_117 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_15_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_12_20 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_50_ clknet_1_0__leaf_CLK _02_ VGND VGND VPWR VPWR clk_div_0.COUNT\[0\] sky130_fd_sc_hs__dfxtp_1
XFILLER_0_5_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_33_ _08_ _14_ _15_ VGND VGND VPWR VPWR _04_ sky130_fd_sc_hs__nor3_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_4_58 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_9_83 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_13_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_9_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_10_113 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_12_98 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XPHY_EDGE_ROW_1_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
X_32_ clk_div_0.COUNT\[1\] clk_div_0.COUNT\[0\] clk_div_0.COUNT\[2\] VGND VGND VPWR
+ VPWR _15_ sky130_fd_sc_hs__a21oi_1
XTAP_TAPCELL_ROW_21_100 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_18_86 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_17_89 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_130 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_1_49 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_144 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_31_ clk_div_0.COUNT\[1\] clk_div_0.COUNT\[0\] clk_div_0.COUNT\[2\] VGND VGND VPWR
+ VPWR _14_ sky130_fd_sc_hs__and3_1
XFILLER_0_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_21_101 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_8_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_12_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_30_ _13_ VGND VGND VPWR VPWR _03_ sky130_fd_sc_hs__clkbuf_1
XTAP_TAPCELL_ROW_21_102 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_3_43 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_18_66 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XPHY_EDGE_ROW_17_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_5_60 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_4_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_21_103 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_18_12 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_18_91 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_2_51 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_3_67 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XTAP_TAPCELL_ROW_18_92 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_2_52 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_2_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_18_58 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_20_48 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_0_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_18_93 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_2_53 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_2_4 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
X_69_ CF[4] net1 CKS VGND VGND VPWR VPWR SWN[4] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_4_90 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_9_35 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_15_8 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_117 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XTAP_TAPCELL_ROW_15_84 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XFILLER_0_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_12_150 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_2_128 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_18_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_68_ CF[5] net1 CKS VGND VGND VPWR VPWR SWN[5] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_0_16 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_16_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XPHY_EDGE_ROW_12_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_21_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XTAP_TAPCELL_ROW_20_96 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XFILLER_0_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XTAP_TAPCELL_ROW_15_85 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
Xclkbuf_1_0__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_1_0__leaf_CLK sky130_fd_sc_hs__clkbuf_16
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
XPHY_EDGE_ROW_0_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hs__decap_4
X_67_ CF[6] net1 CKS VGND VGND VPWR VPWR SWN[6] sky130_fd_sc_hs__dfrtp_1
XFILLER_0_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_1
XFILLER_0_0_28 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_2
XTAP_TAPCELL_ROW_20_97 VGND VPWR sky130_fd_sc_hs__tapvpwrvgnd_1
XFILLER_0_1_71 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
XFILLER_0_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hs__fill_8
.ends

