magic
tech sky130A
magscale 1 2
timestamp 1748962581
<< metal1 >>
rect -268 115138 -258 115238
rect -158 115138 -148 115238
rect -258 113198 -158 115138
rect -58 113198 42 115443
rect 4534 114938 4544 115038
rect 4644 114938 4654 115038
rect 4544 113198 4644 114938
rect 4744 113198 4844 115443
rect 9346 114827 9446 114838
rect 9336 114727 9346 114827
rect 9446 114727 9456 114827
rect 9346 113198 9446 114727
rect 9546 113198 9646 115443
rect 14148 114625 14248 114638
rect 14138 114525 14148 114625
rect 14248 114525 14258 114625
rect 14148 113198 14248 114525
rect 14348 113308 14448 115443
rect 18950 114433 19050 114438
rect 18940 114333 18950 114433
rect 19050 114333 19060 114433
rect 14347 113198 14448 113308
rect 18950 113198 19050 114333
rect 19150 113198 19250 115443
rect 23742 114138 23752 114238
rect 23852 114138 23862 114238
rect 23752 113198 23852 114138
rect 23952 113198 24052 115443
rect 28544 113938 28554 114038
rect 28654 113938 28664 114038
rect 28554 113198 28654 113938
rect 28754 113198 28854 115443
rect 33346 113738 33356 113838
rect 33456 113738 33466 113838
rect 33356 113198 33456 113738
rect 33556 113198 33656 115443
rect 38148 113538 38158 113638
rect 38258 113538 38268 113638
rect 38158 113198 38258 113538
rect 38358 113198 38458 115443
rect 42950 113338 42960 113438
rect 43060 113338 43070 113438
rect 42960 113198 43060 113338
rect 43160 113198 43260 115443
rect -258 -400 -158 1640
rect -268 -500 -258 -400
rect -158 -500 -148 -400
rect -58 -705 42 1440
rect 4544 -200 4644 1640
rect 4534 -300 4544 -200
rect 4644 -300 4654 -200
rect 4744 -705 4844 1440
rect 9346 11 9446 1640
rect 9336 -89 9346 11
rect 9446 -89 9456 11
rect 9346 -100 9446 -89
rect 9546 -705 9646 1440
rect 14148 213 14248 1640
rect 14138 113 14148 213
rect 14248 113 14258 213
rect 14148 100 14248 113
rect 14348 -705 14448 1440
rect 18950 405 19050 1640
rect 18940 305 18950 405
rect 19050 305 19060 405
rect 18950 300 19050 305
rect 19150 -705 19250 1440
rect 23752 600 23852 1640
rect 23742 500 23752 600
rect 23852 500 23862 600
rect 23952 -705 24052 1440
rect 28554 800 28654 1640
rect 28544 700 28554 800
rect 28654 700 28664 800
rect 28754 -705 28854 1440
rect 33356 1000 33456 1640
rect 33346 900 33356 1000
rect 33456 900 33466 1000
rect 33556 -705 33656 1436
rect 38158 1200 38258 1640
rect 38148 1100 38158 1200
rect 38258 1100 38268 1200
rect 38358 -705 38458 1440
rect 42960 1400 43060 1640
rect 42950 1300 42960 1400
rect 43060 1300 43070 1400
rect 43160 -705 43260 1440
<< via1 >>
rect -258 115138 -158 115238
rect 4544 114938 4644 115038
rect 9346 114727 9446 114827
rect 14148 114525 14248 114625
rect 18950 114333 19050 114433
rect 23752 114138 23852 114238
rect 28554 113938 28654 114038
rect 33356 113738 33456 113838
rect 38158 113538 38258 113638
rect 42960 113338 43060 113438
rect -258 -500 -158 -400
rect 4544 -300 4644 -200
rect 9346 -89 9446 11
rect 14148 113 14248 213
rect 18950 305 19050 405
rect 23752 500 23852 600
rect 28554 700 28654 800
rect 33356 900 33456 1000
rect 38158 1100 38258 1200
rect 42960 1300 43060 1400
<< metal2 >>
rect -258 115238 -158 115248
rect -158 115138 50472 115238
rect -258 115128 -158 115138
rect 4544 115038 4644 115048
rect 4644 114938 50272 115038
rect 4544 114928 4644 114938
rect 9346 114827 9446 114837
rect 9446 114727 50072 114827
rect 9346 114717 9446 114727
rect 14148 114625 14248 114635
rect 14248 114526 49872 114625
rect 14248 114525 14347 114526
rect 14148 114515 14248 114525
rect 18950 114433 19050 114443
rect 19050 114333 49672 114433
rect 18950 114323 19050 114333
rect 23752 114238 23852 114248
rect 23852 114138 49472 114238
rect 23752 114128 23852 114138
rect 28554 114038 28654 114048
rect 28654 113938 49272 114038
rect 28554 113928 28654 113938
rect 33356 113838 33456 113848
rect 33456 113738 49072 113838
rect 33356 113728 33456 113738
rect 38158 113638 38258 113648
rect 38258 113538 48872 113638
rect 38158 113528 38258 113538
rect 42960 113438 43060 113448
rect 43060 113338 48672 113438
rect 42960 113328 43060 113338
rect -1088 6313 -948 103865
rect -808 18026 -668 103809
rect -528 18124 -388 98943
rect 47772 3040 47912 111698
rect 48052 2840 48192 111898
rect 48332 1840 48472 112898
rect 42960 1400 43060 1410
rect 48572 1400 48672 113338
rect 43060 1300 48672 1400
rect 42960 1290 43060 1300
rect 38158 1200 38258 1210
rect 48772 1200 48872 113538
rect 38258 1100 48872 1200
rect 38158 1090 38258 1100
rect 33356 1000 33456 1010
rect 48972 1000 49072 113738
rect 33456 900 49072 1000
rect 33356 890 33456 900
rect 28554 800 28654 810
rect 49172 800 49272 113938
rect 28654 700 49272 800
rect 28554 690 28654 700
rect 23752 600 23852 610
rect 49372 600 49472 114138
rect 23852 500 49472 600
rect 23752 490 23852 500
rect 18950 405 19050 415
rect 49572 405 49672 114333
rect 19050 305 49672 405
rect 18950 295 19050 305
rect 14148 213 14248 223
rect 14248 212 14347 213
rect 49772 212 49872 114526
rect 14248 113 49872 212
rect 14148 103 14248 113
rect 9346 11 9446 21
rect 49972 11 50072 114727
rect 9446 -89 50072 11
rect 9346 -99 9446 -89
rect 4544 -200 4644 -190
rect 50172 -200 50272 114938
rect 4644 -300 50272 -200
rect 4544 -310 4644 -300
rect -258 -400 -158 -390
rect 50372 -400 50472 115138
rect -158 -500 50472 -400
rect -258 -510 -158 -500
<< metal4 >>
rect 1586 57728 46080 58450
rect 1586 56288 46080 57010
use single_10b_cdac  single_10b_cdac_0
timestamp 1748851250
transform -1 0 47388 0 1 41235
box -1094 -39935 48486 15775
use single_10b_cdac  single_10b_cdac_1
timestamp 1748851250
transform -1 0 47388 0 -1 73503
box -1094 -39935 48486 15775
<< labels >>
flabel metal1 43180 115367 43240 115427 0 FreeSans 400 0 0 0 SWP_IN[0]
port 0 nsew
flabel metal1 38378 115365 38438 115425 0 FreeSans 400 0 0 0 SWP_IN[1]
port 1 nsew
flabel metal1 33575 115357 33635 115417 0 FreeSans 400 0 0 0 SWP_IN[2]
port 2 nsew
flabel metal1 28774 115364 28834 115424 0 FreeSans 400 0 0 0 SWP_IN[3]
port 3 nsew
flabel metal1 23967 115349 24027 115409 0 FreeSans 400 0 0 0 SWP_IN[4]
port 4 nsew
flabel metal1 19170 115345 19230 115405 0 FreeSans 400 0 0 0 SWP_IN[5]
port 5 nsew
flabel metal1 14367 115362 14427 115422 0 FreeSans 400 0 0 0 SWP_IN[6]
port 6 nsew
flabel metal1 9568 115359 9628 115419 0 FreeSans 400 0 0 0 SWP_IN[7]
port 7 nsew
flabel metal1 4766 115364 4826 115424 0 FreeSans 400 0 0 0 SWP_IN[8]
port 8 nsew
flabel metal1 -37 115370 23 115430 0 FreeSans 400 0 0 0 SWP_IN[9]
port 9 nsew
flabel metal1 43181 -683 43241 -623 0 FreeSans 400 0 0 0 SWN_IN[0]
port 10 nsew
flabel metal1 38375 -683 38435 -623 0 FreeSans 400 0 0 0 SWN_IN[1]
port 11 nsew
flabel metal1 33571 -693 33631 -633 0 FreeSans 400 0 0 0 SWN_IN[2]
port 12 nsew
flabel metal1 28774 -691 28834 -631 0 FreeSans 400 0 0 0 SWN_IN[3]
port 13 nsew
flabel metal1 23968 -689 24028 -629 0 FreeSans 400 0 0 0 SWN_IN[4]
port 14 nsew
flabel metal1 19166 -687 19226 -627 0 FreeSans 400 0 0 0 SWN_IN[5]
port 15 nsew
flabel metal1 14366 -687 14426 -627 0 FreeSans 400 0 0 0 SWN_IN[6]
port 16 nsew
flabel metal1 9562 -683 9622 -623 0 FreeSans 400 0 0 0 SWN_IN[7]
port 17 nsew
flabel metal1 4760 -683 4820 -623 0 FreeSans 400 0 0 0 SWN_IN[8]
port 18 nsew
flabel metal1 -42 -683 18 -623 0 FreeSans 400 0 0 0 SWN_IN[9]
port 19 nsew
flabel metal2 48594 1567 48654 1627 0 FreeSans 400 0 0 0 CF[0]
port 20 nsew
flabel metal2 48796 1577 48856 1637 0 FreeSans 400 0 0 0 CF[1]
port 21 nsew
flabel metal2 48992 1577 49052 1637 0 FreeSans 400 0 0 0 CF[2]
port 22 nsew
flabel metal2 49192 1579 49252 1639 0 FreeSans 400 0 0 0 CF[3]
port 23 nsew
flabel metal2 49390 1577 49450 1637 0 FreeSans 400 0 0 0 CF[4]
port 24 nsew
flabel metal2 49590 1571 49650 1631 0 FreeSans 400 0 0 0 CF[5]
port 25 nsew
flabel metal2 49790 1573 49850 1633 0 FreeSans 400 0 0 0 CF[6]
port 26 nsew
flabel metal2 49996 1567 50056 1627 0 FreeSans 400 0 0 0 CF[7]
port 28 nsew
flabel metal2 50190 1561 50250 1621 0 FreeSans 400 0 0 0 CF[8]
port 29 nsew
flabel metal2 50390 1563 50450 1623 0 FreeSans 400 0 0 0 CF[9]
port 30 nsew
flabel metal2 48373 3281 48433 3341 0 FreeSans 400 0 0 0 VCM
port 31 nsew
flabel metal2 48092 3275 48152 3335 0 FreeSans 400 0 0 0 VDD
port 32 nsew
flabel metal2 47805 3284 47865 3344 0 FreeSans 400 0 0 0 VSS
port 33 nsew
flabel metal4 24857 58063 24917 58123 0 FreeSans 400 0 0 0 VCP
port 34 nsew
flabel metal4 24853 56584 24913 56644 0 FreeSans 400 0 0 0 VCN
port 35 nsew
<< end >>
