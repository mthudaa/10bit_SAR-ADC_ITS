magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect -17 369 13 403
rect 47 369 85 403
rect 119 369 157 403
rect 191 369 229 403
rect 263 369 301 403
rect 335 369 373 403
rect 407 369 445 403
rect 479 369 517 403
rect 551 369 589 403
rect 623 369 661 403
rect 695 369 733 403
rect 767 369 805 403
rect 839 369 877 403
rect 911 369 949 403
rect 983 369 1021 403
rect 1055 369 1093 403
rect 1127 369 1165 403
rect 1199 369 1237 403
rect 1271 369 1309 403
rect 1343 369 1381 403
rect 1415 369 1453 403
rect 1487 369 1525 403
rect 1559 369 1597 403
rect 1631 369 1669 403
rect 1703 369 1741 403
rect 1775 369 1813 403
rect 1847 369 1885 403
rect 1919 369 1957 403
rect 1991 369 2029 403
rect 2063 369 2101 403
rect 2135 369 2173 403
rect 2207 369 2245 403
rect 2279 369 2317 403
rect 2351 369 2389 403
rect 2423 369 2461 403
rect 2495 369 2533 403
rect 2567 369 2605 403
rect 2639 369 2677 403
rect 2711 369 2749 403
rect 2783 369 2821 403
rect 2855 369 2893 403
rect 2927 369 2965 403
rect 2999 369 3037 403
rect 3071 369 3109 403
rect 3143 369 3181 403
rect 3215 369 3253 403
rect 3287 369 3325 403
rect 3359 369 3397 403
rect 3431 369 3469 403
rect 3503 369 3541 403
rect 3575 369 3613 403
rect 3647 369 3685 403
rect 3719 369 3757 403
rect 3791 369 3829 403
rect 3863 369 3901 403
rect 3935 369 3973 403
rect 4007 369 4045 403
rect 4079 369 4117 403
rect 4151 369 4189 403
rect 4223 369 4261 403
rect 4295 369 4333 403
rect 4367 369 4405 403
rect 4439 369 4477 403
rect 4511 369 4549 403
rect 4583 369 4621 403
rect 4655 369 4693 403
rect 4727 369 4765 403
rect 4799 369 4837 403
rect 4871 369 4909 403
rect 4943 369 4981 403
rect 5015 369 5053 403
rect 5087 369 5125 403
rect 5159 369 5197 403
rect 5231 369 5269 403
rect 5303 369 5341 403
rect 5375 369 5413 403
rect 5447 369 5485 403
rect 5519 369 5557 403
rect 5591 369 5629 403
rect 5663 369 5701 403
rect 5735 369 5773 403
rect 5807 369 5845 403
rect 5879 369 5917 403
rect 5951 369 5989 403
rect 6023 369 6061 403
rect 6095 369 6133 403
rect 6167 369 6205 403
rect 6239 369 6277 403
rect 6311 369 6349 403
rect 6383 369 6421 403
rect 6455 369 6493 403
rect 6527 369 6565 403
rect 6599 369 6637 403
rect 6671 369 6709 403
rect 6743 369 6781 403
rect 6815 369 6853 403
rect 6887 369 6925 403
rect 6959 369 6997 403
rect 7031 369 7069 403
rect 7103 369 7141 403
rect 7175 369 7213 403
rect 7247 369 7285 403
rect 7319 369 7357 403
rect 7391 369 7429 403
rect 7463 369 7501 403
rect 7535 369 7573 403
rect 7607 369 7645 403
rect 7679 369 7717 403
rect 7751 369 7789 403
rect 7823 369 7861 403
rect 7895 369 7925 403
rect 7997 -17 8009 17
rect 8043 -17 8081 17
rect 8115 -17 8153 17
rect 8187 -17 8225 17
rect 8259 -17 8297 17
rect 8331 -17 8369 17
rect 8403 -17 8441 17
rect 8475 -17 8513 17
rect 8547 -17 8585 17
rect 8619 -17 8657 17
rect 8691 -17 8729 17
rect 8763 -17 8801 17
rect 8835 -17 8873 17
rect 8907 -17 8945 17
rect 8979 -17 9017 17
rect 9051 -17 9089 17
rect 9123 -17 9161 17
rect 9195 -17 9233 17
rect 9267 -17 9305 17
rect 9339 -17 9377 17
rect 9411 -17 9449 17
rect 9483 -17 9521 17
rect 9555 -17 9593 17
rect 9627 -17 9665 17
rect 9699 -17 9737 17
rect 9771 -17 9809 17
rect 9843 -17 9881 17
rect 9915 -17 9953 17
rect 9987 -17 10025 17
rect 10059 -17 10097 17
rect 10131 -17 10169 17
rect 10203 -17 10241 17
rect 10275 -17 10313 17
rect 10347 -17 10385 17
rect 10419 -17 10457 17
rect 10491 -17 10529 17
rect 10563 -17 10601 17
rect 10635 -17 10673 17
rect 10707 -17 10745 17
rect 10779 -17 10817 17
rect 10851 -17 10889 17
rect 10923 -17 10961 17
rect 10995 -17 11033 17
rect 11067 -17 11105 17
rect 11139 -17 11177 17
rect 11211 -17 11249 17
rect 11283 -17 11321 17
rect 11355 -17 11393 17
rect 11427 -17 11465 17
rect 11499 -17 11537 17
rect 11571 -17 11609 17
rect 11643 -17 11681 17
rect 11715 -17 11753 17
rect 11787 -17 11825 17
rect 11859 -17 11897 17
rect 11931 -17 11969 17
rect 12003 -17 12015 17
<< viali >>
rect 13 369 47 403
rect 85 369 119 403
rect 157 369 191 403
rect 229 369 263 403
rect 301 369 335 403
rect 373 369 407 403
rect 445 369 479 403
rect 517 369 551 403
rect 589 369 623 403
rect 661 369 695 403
rect 733 369 767 403
rect 805 369 839 403
rect 877 369 911 403
rect 949 369 983 403
rect 1021 369 1055 403
rect 1093 369 1127 403
rect 1165 369 1199 403
rect 1237 369 1271 403
rect 1309 369 1343 403
rect 1381 369 1415 403
rect 1453 369 1487 403
rect 1525 369 1559 403
rect 1597 369 1631 403
rect 1669 369 1703 403
rect 1741 369 1775 403
rect 1813 369 1847 403
rect 1885 369 1919 403
rect 1957 369 1991 403
rect 2029 369 2063 403
rect 2101 369 2135 403
rect 2173 369 2207 403
rect 2245 369 2279 403
rect 2317 369 2351 403
rect 2389 369 2423 403
rect 2461 369 2495 403
rect 2533 369 2567 403
rect 2605 369 2639 403
rect 2677 369 2711 403
rect 2749 369 2783 403
rect 2821 369 2855 403
rect 2893 369 2927 403
rect 2965 369 2999 403
rect 3037 369 3071 403
rect 3109 369 3143 403
rect 3181 369 3215 403
rect 3253 369 3287 403
rect 3325 369 3359 403
rect 3397 369 3431 403
rect 3469 369 3503 403
rect 3541 369 3575 403
rect 3613 369 3647 403
rect 3685 369 3719 403
rect 3757 369 3791 403
rect 3829 369 3863 403
rect 3901 369 3935 403
rect 3973 369 4007 403
rect 4045 369 4079 403
rect 4117 369 4151 403
rect 4189 369 4223 403
rect 4261 369 4295 403
rect 4333 369 4367 403
rect 4405 369 4439 403
rect 4477 369 4511 403
rect 4549 369 4583 403
rect 4621 369 4655 403
rect 4693 369 4727 403
rect 4765 369 4799 403
rect 4837 369 4871 403
rect 4909 369 4943 403
rect 4981 369 5015 403
rect 5053 369 5087 403
rect 5125 369 5159 403
rect 5197 369 5231 403
rect 5269 369 5303 403
rect 5341 369 5375 403
rect 5413 369 5447 403
rect 5485 369 5519 403
rect 5557 369 5591 403
rect 5629 369 5663 403
rect 5701 369 5735 403
rect 5773 369 5807 403
rect 5845 369 5879 403
rect 5917 369 5951 403
rect 5989 369 6023 403
rect 6061 369 6095 403
rect 6133 369 6167 403
rect 6205 369 6239 403
rect 6277 369 6311 403
rect 6349 369 6383 403
rect 6421 369 6455 403
rect 6493 369 6527 403
rect 6565 369 6599 403
rect 6637 369 6671 403
rect 6709 369 6743 403
rect 6781 369 6815 403
rect 6853 369 6887 403
rect 6925 369 6959 403
rect 6997 369 7031 403
rect 7069 369 7103 403
rect 7141 369 7175 403
rect 7213 369 7247 403
rect 7285 369 7319 403
rect 7357 369 7391 403
rect 7429 369 7463 403
rect 7501 369 7535 403
rect 7573 369 7607 403
rect 7645 369 7679 403
rect 7717 369 7751 403
rect 7789 369 7823 403
rect 7861 369 7895 403
rect 8009 -17 8043 17
rect 8081 -17 8115 17
rect 8153 -17 8187 17
rect 8225 -17 8259 17
rect 8297 -17 8331 17
rect 8369 -17 8403 17
rect 8441 -17 8475 17
rect 8513 -17 8547 17
rect 8585 -17 8619 17
rect 8657 -17 8691 17
rect 8729 -17 8763 17
rect 8801 -17 8835 17
rect 8873 -17 8907 17
rect 8945 -17 8979 17
rect 9017 -17 9051 17
rect 9089 -17 9123 17
rect 9161 -17 9195 17
rect 9233 -17 9267 17
rect 9305 -17 9339 17
rect 9377 -17 9411 17
rect 9449 -17 9483 17
rect 9521 -17 9555 17
rect 9593 -17 9627 17
rect 9665 -17 9699 17
rect 9737 -17 9771 17
rect 9809 -17 9843 17
rect 9881 -17 9915 17
rect 9953 -17 9987 17
rect 10025 -17 10059 17
rect 10097 -17 10131 17
rect 10169 -17 10203 17
rect 10241 -17 10275 17
rect 10313 -17 10347 17
rect 10385 -17 10419 17
rect 10457 -17 10491 17
rect 10529 -17 10563 17
rect 10601 -17 10635 17
rect 10673 -17 10707 17
rect 10745 -17 10779 17
rect 10817 -17 10851 17
rect 10889 -17 10923 17
rect 10961 -17 10995 17
rect 11033 -17 11067 17
rect 11105 -17 11139 17
rect 11177 -17 11211 17
rect 11249 -17 11283 17
rect 11321 -17 11355 17
rect 11393 -17 11427 17
rect 11465 -17 11499 17
rect 11537 -17 11571 17
rect 11609 -17 11643 17
rect 11681 -17 11715 17
rect 11753 -17 11787 17
rect 11825 -17 11859 17
rect 11897 -17 11931 17
rect 11969 -17 12003 17
<< metal1 >>
rect -53 403 12051 439
rect -53 369 13 403
rect 47 369 85 403
rect 119 369 157 403
rect 191 369 229 403
rect 263 369 301 403
rect 335 369 373 403
rect 407 369 445 403
rect 479 369 517 403
rect 551 369 589 403
rect 623 369 661 403
rect 695 369 733 403
rect 767 369 805 403
rect 839 369 877 403
rect 911 369 949 403
rect 983 369 1021 403
rect 1055 369 1093 403
rect 1127 369 1165 403
rect 1199 369 1237 403
rect 1271 369 1309 403
rect 1343 369 1381 403
rect 1415 369 1453 403
rect 1487 369 1525 403
rect 1559 369 1597 403
rect 1631 369 1669 403
rect 1703 369 1741 403
rect 1775 369 1813 403
rect 1847 369 1885 403
rect 1919 369 1957 403
rect 1991 369 2029 403
rect 2063 369 2101 403
rect 2135 369 2173 403
rect 2207 369 2245 403
rect 2279 369 2317 403
rect 2351 369 2389 403
rect 2423 369 2461 403
rect 2495 369 2533 403
rect 2567 369 2605 403
rect 2639 369 2677 403
rect 2711 369 2749 403
rect 2783 369 2821 403
rect 2855 369 2893 403
rect 2927 369 2965 403
rect 2999 369 3037 403
rect 3071 369 3109 403
rect 3143 369 3181 403
rect 3215 369 3253 403
rect 3287 369 3325 403
rect 3359 369 3397 403
rect 3431 369 3469 403
rect 3503 369 3541 403
rect 3575 369 3613 403
rect 3647 369 3685 403
rect 3719 369 3757 403
rect 3791 369 3829 403
rect 3863 369 3901 403
rect 3935 369 3973 403
rect 4007 369 4045 403
rect 4079 369 4117 403
rect 4151 369 4189 403
rect 4223 369 4261 403
rect 4295 369 4333 403
rect 4367 369 4405 403
rect 4439 369 4477 403
rect 4511 369 4549 403
rect 4583 369 4621 403
rect 4655 369 4693 403
rect 4727 369 4765 403
rect 4799 369 4837 403
rect 4871 369 4909 403
rect 4943 369 4981 403
rect 5015 369 5053 403
rect 5087 369 5125 403
rect 5159 369 5197 403
rect 5231 369 5269 403
rect 5303 369 5341 403
rect 5375 369 5413 403
rect 5447 369 5485 403
rect 5519 369 5557 403
rect 5591 369 5629 403
rect 5663 369 5701 403
rect 5735 369 5773 403
rect 5807 369 5845 403
rect 5879 369 5917 403
rect 5951 369 5989 403
rect 6023 369 6061 403
rect 6095 369 6133 403
rect 6167 369 6205 403
rect 6239 369 6277 403
rect 6311 369 6349 403
rect 6383 369 6421 403
rect 6455 369 6493 403
rect 6527 369 6565 403
rect 6599 369 6637 403
rect 6671 369 6709 403
rect 6743 369 6781 403
rect 6815 369 6853 403
rect 6887 369 6925 403
rect 6959 369 6997 403
rect 7031 369 7069 403
rect 7103 369 7141 403
rect 7175 369 7213 403
rect 7247 369 7285 403
rect 7319 369 7357 403
rect 7391 369 7429 403
rect 7463 369 7501 403
rect 7535 369 7573 403
rect 7607 369 7645 403
rect 7679 369 7717 403
rect 7751 369 7789 403
rect 7823 369 7861 403
rect 7895 369 12051 403
rect -53 363 12051 369
rect -53 289 11841 323
rect -53 147 125 239
rect 11873 147 12051 239
rect 166 63 12051 97
rect -53 17 12051 23
rect -53 -17 8009 17
rect 8043 -17 8081 17
rect 8115 -17 8153 17
rect 8187 -17 8225 17
rect 8259 -17 8297 17
rect 8331 -17 8369 17
rect 8403 -17 8441 17
rect 8475 -17 8513 17
rect 8547 -17 8585 17
rect 8619 -17 8657 17
rect 8691 -17 8729 17
rect 8763 -17 8801 17
rect 8835 -17 8873 17
rect 8907 -17 8945 17
rect 8979 -17 9017 17
rect 9051 -17 9089 17
rect 9123 -17 9161 17
rect 9195 -17 9233 17
rect 9267 -17 9305 17
rect 9339 -17 9377 17
rect 9411 -17 9449 17
rect 9483 -17 9521 17
rect 9555 -17 9593 17
rect 9627 -17 9665 17
rect 9699 -17 9737 17
rect 9771 -17 9809 17
rect 9843 -17 9881 17
rect 9915 -17 9953 17
rect 9987 -17 10025 17
rect 10059 -17 10097 17
rect 10131 -17 10169 17
rect 10203 -17 10241 17
rect 10275 -17 10313 17
rect 10347 -17 10385 17
rect 10419 -17 10457 17
rect 10491 -17 10529 17
rect 10563 -17 10601 17
rect 10635 -17 10673 17
rect 10707 -17 10745 17
rect 10779 -17 10817 17
rect 10851 -17 10889 17
rect 10923 -17 10961 17
rect 10995 -17 11033 17
rect 11067 -17 11105 17
rect 11139 -17 11177 17
rect 11211 -17 11249 17
rect 11283 -17 11321 17
rect 11355 -17 11393 17
rect 11427 -17 11465 17
rect 11499 -17 11537 17
rect 11571 -17 11609 17
rect 11643 -17 11681 17
rect 11715 -17 11753 17
rect 11787 -17 11825 17
rect 11859 -17 11897 17
rect 11931 -17 11969 17
rect 12003 -17 12051 17
rect -53 -53 12051 -17
use sky130_fd_pr__pfet_01v8_D9QHA6  XM1
timestamp 1750100919
transform 0 1 3954 -1 0 193
box -246 -4007 246 4007
use sky130_fd_pr__nfet_01v8_DPTN2D  XM2
timestamp 1750100919
transform 0 1 10006 -1 0 193
box -236 -2035 236 2035
<< labels >>
flabel metal1 s -38 401 -28 412 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s -39 -34 -29 -23 0 FreeSans 500 0 0 0 VSS
port 2 nsew
flabel metal1 s -39 189 -29 200 0 FreeSans 500 0 0 0 SWP
port 3 nsew
flabel metal1 s -44 299 -34 310 0 FreeSans 500 0 0 0 IN
port 4 nsew
flabel metal1 s 12024 181 12035 195 0 FreeSans 500 0 0 0 SWN
port 5 nsew
flabel metal1 s 12032 73 12043 87 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
