magic
tech sky130A
magscale 1 2
timestamp 1748803925
<< metal1 >>
rect 1421 2274 14902 2574
rect -519 260 -379 360
rect -279 260 -269 360
rect -519 60 -179 160
rect -79 60 -69 160
rect 8488 -2528 13626 -2228
rect -519 -4542 -379 -4442
rect -279 -4542 -269 -4442
rect -519 -4742 -179 -4642
rect -79 -4742 -69 -4642
rect 1421 -7330 12350 -7030
rect -519 -9344 -383 -9244
rect -283 -9344 -273 -9244
rect -519 -9544 -179 -9444
rect -79 -9544 -69 -9444
rect 1421 -12132 11074 -11832
rect -519 -14146 -379 -14046
rect -279 -14146 -269 -14046
rect -189 -14246 -179 -14245
rect -519 -14345 -179 -14246
rect -79 -14345 -69 -14245
rect -519 -14346 -79 -14345
rect 1421 -16934 9798 -16634
rect -519 -18948 -379 -18848
rect -279 -18948 -269 -18848
rect -519 -19148 -179 -19048
rect -79 -19148 -69 -19048
rect 1631 -21736 8522 -21436
rect -519 -23750 -379 -23650
rect -279 -23750 -269 -23650
rect -519 -23950 -179 -23850
rect -79 -23950 -69 -23850
rect 4208 -26538 7246 -26238
rect -519 -28453 -279 -28452
rect -519 -28552 -379 -28453
rect -389 -28553 -379 -28552
rect -279 -28553 -269 -28453
rect -519 -28752 -179 -28652
rect -79 -28752 -69 -28652
rect 1421 -31340 5970 -31040
rect -519 -33354 -379 -33254
rect -279 -33354 -269 -33254
rect -519 -33554 -179 -33454
rect -79 -33554 -69 -33454
rect 2978 -36142 4694 -35842
rect -519 -38156 -379 -38056
rect -279 -38156 -269 -38056
rect -519 -38356 -179 -38256
rect -79 -38356 -69 -38256
rect 2277 -40944 3418 -40644
rect -519 -42958 -379 -42858
rect -279 -42958 -269 -42858
rect -519 -43158 -179 -43058
rect -79 -43158 -69 -43058
<< via1 >>
rect -379 260 -279 360
rect -179 60 -79 160
rect -379 -4542 -279 -4442
rect -179 -4742 -79 -4642
rect -383 -9344 -283 -9244
rect -179 -9544 -79 -9444
rect -379 -14146 -279 -14046
rect -179 -14345 -79 -14245
rect -379 -18948 -279 -18848
rect -179 -19148 -79 -19048
rect -379 -23750 -279 -23650
rect -179 -23950 -79 -23850
rect -379 -28553 -279 -28453
rect -179 -28752 -79 -28652
rect -379 -33354 -279 -33254
rect -179 -33554 -79 -33454
rect -379 -38156 -279 -38056
rect -179 -38356 -79 -38256
rect -379 -42958 -279 -42858
rect -179 -43158 -79 -43058
<< metal2 >>
rect -379 360 -279 370
rect -379 250 -279 260
rect -179 160 -79 170
rect -179 50 -79 60
rect -379 -4442 -279 -4432
rect -379 -4552 -279 -4542
rect -179 -4642 -79 -4632
rect -179 -4752 -79 -4742
rect -383 -9244 -283 -9234
rect -383 -9354 -283 -9344
rect -179 -9444 -79 -9434
rect -179 -9554 -79 -9544
rect -379 -14046 -279 -14036
rect -379 -14156 -279 -14146
rect -179 -14245 -79 -14235
rect -179 -14355 -79 -14345
rect -379 -18848 -279 -18835
rect -379 -18958 -279 -18948
rect -179 -19048 -79 -19038
rect -179 -19158 -79 -19148
rect -379 -23650 -279 -23640
rect -379 -23760 -279 -23750
rect -179 -23850 -79 -23840
rect -179 -23960 -79 -23950
rect -379 -28453 -279 -28443
rect -379 -28563 -279 -28553
rect -179 -28652 -79 -28642
rect -179 -28762 -79 -28752
rect -379 -33254 -279 -33244
rect -379 -33364 -279 -33354
rect -179 -33454 -79 -33444
rect -179 -33564 -79 -33554
rect -379 -38056 -279 -38046
rect -379 -38166 -279 -38156
rect -179 -38256 -79 -38246
rect -179 -38366 -79 -38356
rect -379 -42858 -279 -42848
rect 21 -42880 121 4462
rect 1021 -42907 1121 4728
rect 1221 -42872 1321 4634
rect -379 -42968 -279 -42958
rect -179 -43058 -79 -43048
rect -179 -43168 -79 -43158
use cdac_sw_1  cdac_sw_1_0
timestamp 1748800002
transform 1 0 1439 0 1 3332
box -1828 -3272 13573 1410
use cdac_sw_2  cdac_sw_2_0
timestamp 1748789316
transform 1 0 1439 0 1 -1470
box -1828 -3272 12297 1410
use cdac_sw_3  cdac_sw_3_0
timestamp 1748790148
transform 1 0 1439 0 1 -6272
box -1828 -3272 11021 1410
use cdac_sw_4  cdac_sw_4_0
timestamp 1748792579
transform 1 0 1439 0 1 -11074
box -1828 -3272 9745 1410
use cdac_sw_5  cdac_sw_5_0
timestamp 1748794220
transform 1 0 1439 0 1 -15876
box -1828 -3272 8469 1410
use cdac_sw_6  cdac_sw_6_0
timestamp 1748794577
transform 1 0 1439 0 1 -20678
box -1828 -3272 7193 1410
use cdac_sw_7  cdac_sw_7_0
timestamp 1748795123
transform 1 0 1439 0 1 -25480
box -1828 -3272 5917 1410
use cdac_sw_8  cdac_sw_8_0
timestamp 1748795623
transform 1 0 1439 0 1 -30282
box -1828 -3272 4641 1410
use cdac_sw_9  cdac_sw_9_0
timestamp 1748796169
transform 1 0 1439 0 1 -35084
box -1828 -3272 3610 1410
use cdac_sw_10  cdac_sw_10_0
timestamp 1748803164
transform 1 0 1439 0 1 -39886
box -1828 -3272 3610 1410
<< labels >>
flabel metal2 1052 4651 1092 4691 0 FreeSans 800 0 0 0 VDD
port 0 nsew
flabel metal2 1249 4437 1289 4477 0 FreeSans 800 0 0 0 VSS
port 1 nsew
flabel metal2 55 4351 95 4391 0 FreeSans 800 0 0 0 VCM
port 2 nsew
flabel metal1 -501 281 -461 321 0 FreeSans 800 0 0 0 SW_IN[0]
port 3 nsew
flabel metal1 -492 -4511 -452 -4471 0 FreeSans 800 0 0 0 SW_IN[1]
port 4 nsew
flabel metal1 -503 -9309 -463 -9269 0 FreeSans 800 0 0 0 SW_IN[2]
port 5 nsew
flabel metal1 -499 -14115 -459 -14075 0 FreeSans 800 0 0 0 SW_IN[3]
port 6 nsew
flabel metal1 -503 -18914 -463 -18874 0 FreeSans 800 0 0 0 SW_IN[4]
port 7 nsew
flabel metal1 -498 -23716 -458 -23676 0 FreeSans 800 0 0 0 SW_IN[5]
port 8 nsew
flabel metal1 -500 -28521 -460 -28481 0 FreeSans 800 0 0 0 SW_IN[6]
port 9 nsew
flabel metal1 -497 -33321 -457 -33281 0 FreeSans 800 0 0 0 SW_IN[7]
port 10 nsew
flabel metal1 -496 -38127 -456 -38087 0 FreeSans 800 0 0 0 SW_IN[8]
port 11 nsew
flabel metal1 -492 -42927 -452 -42887 0 FreeSans 800 0 0 0 SW_IN[9]
port 12 nsew
flabel metal1 -496 88 -456 128 0 FreeSans 800 0 0 0 CF[0]
port 13 nsew
flabel metal1 -497 -4710 -457 -4670 0 FreeSans 800 0 0 0 CF[1]
port 14 nsew
flabel metal1 -500 -9513 -460 -9473 0 FreeSans 800 0 0 0 CF[2]
port 15 nsew
flabel metal1 -490 -14319 -450 -14279 0 FreeSans 800 0 0 0 CF[3]
port 16 nsew
flabel metal1 -497 -19117 -457 -19077 0 FreeSans 800 0 0 0 CF[4]
port 17 nsew
flabel metal1 -495 -23917 -455 -23877 0 FreeSans 800 0 0 0 CF[5]
port 18 nsew
flabel metal1 -500 -28722 -460 -28682 0 FreeSans 800 0 0 0 CF[6]
port 19 nsew
flabel metal1 -497 -33525 -457 -33485 0 FreeSans 800 0 0 0 CF[7]
port 20 nsew
flabel metal1 -495 -38323 -455 -38283 0 FreeSans 800 0 0 0 CF[8]
port 21 nsew
flabel metal1 -500 -43131 -460 -43091 0 FreeSans 800 0 0 0 CF[9]
port 22 nsew
flabel metal1 14719 2393 14759 2433 0 FreeSans 800 0 0 0 SWN[0]
port 23 nsew
flabel metal1 13429 -2410 13469 -2370 0 FreeSans 800 0 0 0 SWN[1]
port 24 nsew
flabel metal1 12158 -7204 12198 -7164 0 FreeSans 800 0 0 0 SWN[2]
port 25 nsew
flabel metal1 10887 -11997 10927 -11957 0 FreeSans 800 0 0 0 SWN[3]
port 26 nsew
flabel metal1 9616 -16801 9656 -16761 0 FreeSans 800 0 0 0 SWN[4]
port 27 nsew
flabel metal1 8331 -21599 8371 -21559 0 FreeSans 800 0 0 0 SWN[5]
port 28 nsew
flabel metal1 7065 -26418 7105 -26378 0 FreeSans 800 0 0 0 SWN[6]
port 29 nsew
flabel metal1 5784 -31216 5824 -31176 0 FreeSans 800 0 0 0 SWN[7]
port 30 nsew
flabel metal1 4504 -36010 4544 -35970 0 FreeSans 800 0 0 0 SWN[8]
port 31 nsew
flabel metal1 3223 -40818 3263 -40778 0 FreeSans 800 0 0 0 SWN[9]
port 32 nsew
<< end >>
