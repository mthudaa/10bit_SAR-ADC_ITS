magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< metal1 >>
rect -20212 -12192 -19884 -12166
rect -20212 -12244 -20176 -12192
rect -20124 -12244 -19972 -12192
rect -19920 -12244 -19884 -12192
rect -20212 -12270 -19884 -12244
rect -22696 -14432 -21500 -14406
rect -22696 -14484 -22660 -14432
rect -22608 -14484 -21588 -14432
rect -21536 -14484 -21500 -14432
rect -22696 -14510 -21500 -14484
rect -21628 -15552 -21504 -15526
rect -21628 -15604 -21592 -15552
rect -21540 -15604 -21504 -15552
rect -21628 -15630 -21504 -15604
rect -21618 -18886 -21514 -15630
rect -20216 -16672 -20092 -16646
rect -20216 -16724 -20180 -16672
rect -20128 -16724 -20092 -16672
rect -20216 -16750 -20092 -16724
rect -20206 -17910 -20102 -16750
rect -20216 -17936 -20092 -17910
rect -20216 -17988 -20180 -17936
rect -20128 -17988 -20092 -17936
rect -20216 -18014 -20092 -17988
rect -21628 -18912 -21504 -18886
rect -21628 -18964 -21592 -18912
rect -21540 -18964 -21504 -18912
rect -21628 -18990 -21504 -18964
rect -22488 -20312 -22364 -20286
rect -22488 -20364 -22452 -20312
rect -22400 -20364 -22364 -20312
rect -22488 -20390 -22364 -20364
rect -21628 -20312 -21504 -20286
rect -21628 -20364 -21592 -20312
rect -21540 -20364 -21504 -20312
rect -21628 -20390 -21504 -20364
rect -22478 -21406 -22374 -20390
rect -21618 -21406 -21514 -20390
rect -22488 -21432 -22364 -21406
rect -22488 -21484 -22452 -21432
rect -22400 -21484 -22364 -21432
rect -22488 -21510 -22364 -21484
rect -21628 -21432 -21504 -21406
rect -21628 -21484 -21592 -21432
rect -21540 -21484 -21504 -21432
rect -21628 -21510 -21504 -21484
rect -20216 -24792 -20092 -24766
rect -20216 -24844 -20180 -24792
rect -20128 -24844 -20092 -24792
rect -20216 -24870 -20092 -24844
rect -20206 -25886 -20102 -24870
rect -20216 -25912 -20092 -25886
rect -20216 -25964 -20180 -25912
rect -20128 -25964 -20092 -25912
rect -20216 -25990 -20092 -25964
rect -21628 -32632 -21504 -32606
rect -21628 -32684 -21592 -32632
rect -21540 -32684 -21504 -32632
rect -21628 -32710 -21504 -32684
rect -21618 -33726 -21514 -32710
rect -21628 -33752 -21504 -33726
rect -21628 -33804 -21592 -33752
rect -21540 -33804 -21504 -33752
rect -21628 -33830 -21504 -33804
rect -18800 -34592 -18676 -34566
rect -18800 -34606 -18764 -34592
rect -23036 -34632 -18764 -34606
rect -23036 -34684 -23016 -34632
rect -22964 -34684 -22952 -34632
rect -22900 -34684 -22888 -34632
rect -22836 -34644 -18764 -34632
rect -18712 -34606 -18676 -34592
rect -18712 -34632 -18336 -34606
rect -18712 -34644 -18424 -34632
rect -22836 -34684 -18424 -34644
rect -18372 -34684 -18336 -34632
rect -23036 -34710 -18336 -34684
rect -24448 -34845 -17060 -34819
rect -24448 -34897 -24412 -34845
rect -24360 -34897 -17352 -34845
rect -17300 -34897 -17148 -34845
rect -17096 -34897 -17060 -34845
rect -24448 -34923 -17060 -34897
rect -27272 -35053 -14440 -35027
rect -27272 -35105 -27236 -35053
rect -27184 -35105 -27032 -35053
rect -26980 -35105 -14524 -35053
rect -14472 -35105 -14440 -35053
rect -27272 -35131 -14440 -35105
rect -32920 -35260 -8588 -35234
rect -32920 -35312 -32884 -35260
rect -32832 -35312 -8876 -35260
rect -8824 -35312 -8676 -35260
rect -8624 -35312 -8588 -35260
rect -32920 -35338 -8588 -35312
rect -45174 -35960 2594 -35934
rect -45174 -36012 -20180 -35960
rect -20128 -36012 2594 -35960
rect -45174 -36038 2594 -36012
rect -45174 -36168 2594 -36142
rect -45174 -36220 -21144 -36168
rect -21092 -36220 2594 -36168
rect -45174 -36246 2594 -36220
rect -45174 -36376 2594 -36350
rect -45174 -36428 -22452 -36376
rect -22400 -36428 2594 -36376
rect -45174 -36454 2594 -36428
rect -45174 -36584 2594 -36558
rect -45174 -36636 -21592 -36584
rect -21540 -36636 2594 -36584
rect -45174 -36662 2594 -36636
rect -45174 -36792 2594 -36766
rect -45174 -36844 -22660 -36792
rect -22608 -36844 2594 -36792
rect -45174 -36870 2594 -36844
rect -45174 -37000 2594 -36974
rect -45174 -37052 -19972 -37000
rect -19920 -37052 2594 -37000
rect -45174 -37078 2594 -37052
rect -45174 -37208 2594 -37182
rect -45174 -37260 -21384 -37208
rect -21332 -37260 2594 -37208
rect -45174 -37286 2594 -37260
rect -45174 -37416 2594 -37390
rect -45174 -37468 -18424 -37416
rect -18372 -37468 2594 -37416
rect -45174 -37494 2594 -37468
rect -45174 -37624 2594 -37598
rect -45174 -37676 -17148 -37624
rect -17096 -37676 2594 -37624
rect -45174 -37702 2594 -37676
rect -45174 -37832 2594 -37806
rect -45174 -37884 -27032 -37832
rect -26980 -37884 2594 -37832
rect -45174 -37910 2594 -37884
rect -45174 -38040 2594 -38014
rect -45174 -38092 -8676 -38040
rect -8624 -38092 2594 -38040
rect -45174 -38118 2594 -38092
<< via1 >>
rect -20176 -12244 -20124 -12192
rect -19972 -12244 -19920 -12192
rect -22660 -14484 -22608 -14432
rect -21588 -14484 -21536 -14432
rect -21592 -15604 -21540 -15552
rect -20180 -16724 -20128 -16672
rect -20180 -17988 -20128 -17936
rect -21592 -18964 -21540 -18912
rect -22452 -20364 -22400 -20312
rect -21592 -20364 -21540 -20312
rect -22452 -21484 -22400 -21432
rect -21592 -21484 -21540 -21432
rect -20180 -24844 -20128 -24792
rect -20180 -25964 -20128 -25912
rect -21592 -32684 -21540 -32632
rect -21592 -33804 -21540 -33752
rect -23016 -34684 -22964 -34632
rect -22952 -34684 -22900 -34632
rect -22888 -34684 -22836 -34632
rect -18764 -34644 -18712 -34592
rect -18424 -34684 -18372 -34632
rect -24412 -34897 -24360 -34845
rect -17352 -34897 -17300 -34845
rect -17148 -34897 -17096 -34845
rect -27236 -35105 -27184 -35053
rect -27032 -35105 -26980 -35053
rect -14524 -35105 -14472 -35053
rect -32884 -35312 -32832 -35260
rect -8876 -35312 -8824 -35260
rect -8676 -35312 -8624 -35260
rect -20180 -36012 -20128 -35960
rect -21144 -36220 -21092 -36168
rect -22452 -36428 -22400 -36376
rect -21592 -36636 -21540 -36584
rect -22660 -36844 -22608 -36792
rect -19972 -37052 -19920 -37000
rect -21384 -37260 -21332 -37208
rect -18424 -37468 -18372 -37416
rect -17148 -37676 -17096 -37624
rect -27032 -37884 -26980 -37832
rect -8676 -38092 -8624 -38040
<< metal2 >>
rect -21614 -7686 -21510 -7676
rect -21614 -7710 -21306 -7686
rect -21614 -7766 -21590 -7710
rect -21534 -7766 -21306 -7710
rect -21614 -7790 -21306 -7766
rect -21614 -7800 -21510 -7790
rect -22686 -14432 -22582 -14396
rect -22686 -14484 -22660 -14432
rect -22608 -14484 -22582 -14432
rect -22686 -21126 -22582 -14484
rect -21614 -14430 -21510 -14396
rect -21614 -14486 -21590 -14430
rect -21534 -14486 -21510 -14430
rect -21614 -14520 -21510 -14486
rect -21618 -15550 -21514 -15516
rect -21618 -15606 -21594 -15550
rect -21538 -15606 -21514 -15550
rect -21618 -15640 -21514 -15606
rect -21614 -17766 -21510 -17756
rect -22478 -17790 -21510 -17766
rect -22478 -17846 -21590 -17790
rect -21534 -17846 -21510 -17790
rect -22478 -17870 -21510 -17846
rect -22478 -20312 -22374 -17870
rect -21614 -17880 -21510 -17870
rect -22478 -20364 -22452 -20312
rect -22400 -20364 -22374 -20312
rect -22478 -20400 -22374 -20364
rect -21618 -18910 -21514 -18876
rect -21618 -18966 -21594 -18910
rect -21538 -18966 -21514 -18910
rect -21618 -20312 -21514 -18966
rect -21618 -20364 -21592 -20312
rect -21540 -20364 -21514 -20312
rect -21618 -20400 -21514 -20364
rect -21614 -21126 -21510 -21116
rect -22686 -21150 -21510 -21126
rect -22686 -21206 -21590 -21150
rect -21534 -21206 -21510 -21150
rect -22686 -21230 -21510 -21206
rect -32910 -34590 -32806 -34556
rect -32910 -34646 -32886 -34590
rect -32830 -34646 -32806 -34590
rect -32910 -35260 -32806 -34646
rect -27262 -34576 -27158 -34556
rect -27262 -34590 -27062 -34576
rect -27262 -34646 -27238 -34590
rect -27182 -34646 -27062 -34590
rect -27262 -34682 -27062 -34646
rect -24438 -34590 -24334 -34556
rect -24438 -34646 -24414 -34590
rect -24358 -34646 -24334 -34590
rect -27262 -35053 -27158 -34682
rect -24438 -34845 -24334 -34646
rect -23026 -34576 -22922 -34556
rect -23026 -34590 -22826 -34576
rect -23026 -34632 -23002 -34590
rect -22946 -34632 -22826 -34590
rect -23026 -34684 -23016 -34632
rect -22964 -34684 -22952 -34646
rect -22900 -34684 -22888 -34632
rect -22836 -34684 -22826 -34632
rect -23026 -34720 -22826 -34684
rect -24438 -34897 -24412 -34845
rect -24360 -34897 -24334 -34845
rect -24438 -34933 -24334 -34897
rect -27262 -35105 -27236 -35053
rect -27184 -35105 -27158 -35053
rect -27262 -35141 -27158 -35105
rect -27058 -35053 -26954 -35017
rect -27058 -35105 -27032 -35053
rect -26980 -35105 -26954 -35053
rect -32910 -35312 -32884 -35260
rect -32832 -35312 -32806 -35260
rect -32910 -35348 -32806 -35312
rect -27058 -37832 -26954 -35105
rect -22686 -36792 -22582 -21230
rect -21614 -21240 -21510 -21230
rect -22478 -21432 -22374 -21396
rect -22478 -21484 -22452 -21432
rect -22400 -21484 -22374 -21432
rect -22478 -36376 -22374 -21484
rect -21618 -21432 -21514 -21396
rect -21618 -21484 -21592 -21432
rect -21540 -21484 -21514 -21432
rect -21618 -32632 -21514 -21484
rect -21618 -32684 -21592 -32632
rect -21540 -32684 -21514 -32632
rect -21618 -32720 -21514 -32684
rect -21614 -33446 -21510 -33436
rect -21410 -33446 -21306 -7790
rect -20202 -12190 -20098 -12156
rect -20202 -12246 -20178 -12190
rect -20122 -12246 -20098 -12190
rect -20202 -12280 -20098 -12246
rect -19998 -12192 -19894 -12156
rect -19998 -12244 -19972 -12192
rect -19920 -12244 -19894 -12192
rect -20206 -16670 -20102 -16636
rect -20206 -16726 -20182 -16670
rect -20126 -16726 -20102 -16670
rect -20206 -16760 -20102 -16726
rect -20206 -17070 -20102 -17060
rect -21614 -33470 -21306 -33446
rect -21614 -33526 -21590 -33470
rect -21534 -33526 -21306 -33470
rect -21614 -33550 -21306 -33526
rect -21614 -33560 -21510 -33550
rect -22478 -36428 -22452 -36376
rect -22400 -36428 -22374 -36376
rect -22478 -36464 -22374 -36428
rect -21618 -33752 -21514 -33716
rect -21618 -33804 -21592 -33752
rect -21540 -33804 -21514 -33752
rect -21618 -36584 -21514 -33804
rect -21618 -36636 -21592 -36584
rect -21540 -36636 -21514 -36584
rect -21618 -36672 -21514 -36636
rect -22686 -36844 -22660 -36792
rect -22608 -36844 -22582 -36792
rect -22686 -36880 -22582 -36844
rect -21410 -37208 -21306 -33550
rect -21170 -17094 -20102 -17070
rect -21170 -17150 -20182 -17094
rect -20126 -17150 -20102 -17094
rect -21170 -17174 -20102 -17150
rect -21170 -36168 -21066 -17174
rect -20206 -17184 -20102 -17174
rect -20206 -17936 -20102 -17900
rect -20206 -17988 -20180 -17936
rect -20128 -17988 -20102 -17936
rect -20206 -24792 -20102 -17988
rect -20206 -24844 -20180 -24792
rect -20128 -24844 -20102 -24792
rect -20206 -24880 -20102 -24844
rect -20202 -25606 -20098 -25596
rect -19998 -25606 -19894 -12244
rect -20202 -25630 -19894 -25606
rect -20202 -25686 -20178 -25630
rect -20122 -25686 -19894 -25630
rect -20202 -25710 -19894 -25686
rect -20202 -25720 -20098 -25710
rect -20206 -25912 -20102 -25876
rect -20206 -25964 -20180 -25912
rect -20128 -25964 -20102 -25912
rect -20206 -35960 -20102 -25964
rect -20206 -36012 -20180 -35960
rect -20128 -36012 -20102 -35960
rect -20206 -36048 -20102 -36012
rect -21170 -36220 -21144 -36168
rect -21092 -36220 -21066 -36168
rect -21170 -36256 -21066 -36220
rect -19998 -37000 -19894 -25710
rect -18790 -34590 -18686 -34556
rect -18790 -34646 -18766 -34590
rect -18710 -34646 -18686 -34590
rect -17378 -34576 -17274 -34555
rect -17378 -34589 -17178 -34576
rect -18790 -34680 -18686 -34646
rect -18450 -34632 -18346 -34596
rect -19998 -37052 -19972 -37000
rect -19920 -37052 -19894 -37000
rect -19998 -37088 -19894 -37052
rect -18450 -34684 -18424 -34632
rect -18372 -34684 -18346 -34632
rect -21410 -37260 -21384 -37208
rect -21332 -37260 -21306 -37208
rect -21410 -37296 -21306 -37260
rect -18450 -37416 -18346 -34684
rect -17378 -34645 -17354 -34589
rect -17298 -34645 -17178 -34589
rect -17378 -34682 -17178 -34645
rect -14546 -34594 -14450 -34564
rect -14546 -34650 -14526 -34594
rect -14470 -34650 -14450 -34594
rect -17378 -34845 -17274 -34682
rect -17378 -34897 -17352 -34845
rect -17300 -34897 -17274 -34845
rect -17378 -34933 -17274 -34897
rect -17174 -34845 -17070 -34809
rect -17174 -34897 -17148 -34845
rect -17096 -34897 -17070 -34845
rect -18450 -37468 -18424 -37416
rect -18372 -37468 -18346 -37416
rect -18450 -37504 -18346 -37468
rect -17174 -37624 -17070 -34897
rect -14546 -35053 -14450 -34650
rect -14546 -35105 -14524 -35053
rect -14472 -35105 -14450 -35053
rect -14546 -35141 -14450 -35105
rect -8898 -34594 -8802 -34564
rect -8898 -34650 -8878 -34594
rect -8822 -34650 -8802 -34594
rect -8898 -35260 -8802 -34650
rect -8898 -35312 -8876 -35260
rect -8824 -35312 -8802 -35260
rect -8898 -35348 -8802 -35312
rect -8702 -35260 -8598 -35224
rect -8702 -35312 -8676 -35260
rect -8624 -35312 -8598 -35260
rect -17174 -37676 -17148 -37624
rect -17096 -37676 -17070 -37624
rect -17174 -37712 -17070 -37676
rect -27058 -37884 -27032 -37832
rect -26980 -37884 -26954 -37832
rect -27058 -37920 -26954 -37884
rect -8702 -38040 -8598 -35312
rect -8702 -38092 -8676 -38040
rect -8624 -38092 -8598 -38040
rect -8702 -38128 -8598 -38092
<< via2 >>
rect -21590 -7766 -21534 -7710
rect -21590 -14432 -21534 -14430
rect -21590 -14484 -21588 -14432
rect -21588 -14484 -21536 -14432
rect -21536 -14484 -21534 -14432
rect -21590 -14486 -21534 -14484
rect -21594 -15552 -21538 -15550
rect -21594 -15604 -21592 -15552
rect -21592 -15604 -21540 -15552
rect -21540 -15604 -21538 -15552
rect -21594 -15606 -21538 -15604
rect -21590 -17846 -21534 -17790
rect -21594 -18912 -21538 -18910
rect -21594 -18964 -21592 -18912
rect -21592 -18964 -21540 -18912
rect -21540 -18964 -21538 -18912
rect -21594 -18966 -21538 -18964
rect -21590 -21206 -21534 -21150
rect -32886 -34646 -32830 -34590
rect -27238 -34646 -27182 -34590
rect -24414 -34646 -24358 -34590
rect -23002 -34632 -22946 -34590
rect -23002 -34646 -22964 -34632
rect -22964 -34646 -22952 -34632
rect -22952 -34646 -22946 -34632
rect -20178 -12192 -20122 -12190
rect -20178 -12244 -20176 -12192
rect -20176 -12244 -20124 -12192
rect -20124 -12244 -20122 -12192
rect -20178 -12246 -20122 -12244
rect -20182 -16672 -20126 -16670
rect -20182 -16724 -20180 -16672
rect -20180 -16724 -20128 -16672
rect -20128 -16724 -20126 -16672
rect -20182 -16726 -20126 -16724
rect -21590 -33526 -21534 -33470
rect -20182 -17150 -20126 -17094
rect -20178 -25686 -20122 -25630
rect -18766 -34592 -18710 -34590
rect -18766 -34644 -18764 -34592
rect -18764 -34644 -18712 -34592
rect -18712 -34644 -18710 -34592
rect -18766 -34646 -18710 -34644
rect -17354 -34645 -17298 -34589
rect -14526 -34650 -14470 -34594
rect -8878 -34650 -8822 -34594
<< metal3 >>
rect -21624 -7710 -21500 -7681
rect -21624 -7766 -21590 -7710
rect -21534 -7766 -21500 -7710
rect -21624 -7795 -21500 -7766
rect -21520 -7918 -19992 -7910
rect -21520 -7982 -21494 -7918
rect -21430 -7982 -20082 -7918
rect -20018 -7982 -19992 -7918
rect -21520 -7990 -19992 -7982
rect -20212 -12190 -20088 -12161
rect -20212 -12246 -20178 -12190
rect -20122 -12246 -20088 -12190
rect -20212 -12275 -20088 -12246
rect -21520 -12398 -19992 -12390
rect -21520 -12462 -21494 -12398
rect -21430 -12462 -20082 -12398
rect -20018 -12462 -19992 -12398
rect -21520 -12470 -19992 -12462
rect -21624 -14430 -21500 -14401
rect -21624 -14486 -21590 -14430
rect -21534 -14486 -21500 -14430
rect -21624 -14515 -21500 -14486
rect -21520 -14638 -19992 -14630
rect -21520 -14702 -21494 -14638
rect -21430 -14702 -20082 -14638
rect -20018 -14702 -19992 -14638
rect -21520 -14710 -19992 -14702
rect -21628 -15550 -21504 -15521
rect -21628 -15606 -21594 -15550
rect -21538 -15606 -21504 -15550
rect -21628 -15635 -21504 -15606
rect -21520 -15758 -19992 -15750
rect -21520 -15822 -21494 -15758
rect -21430 -15822 -20082 -15758
rect -20018 -15822 -19992 -15758
rect -21520 -15830 -19992 -15822
rect -20216 -16670 -20092 -16641
rect -20216 -16726 -20182 -16670
rect -20126 -16726 -20092 -16670
rect -20216 -16755 -20092 -16726
rect -20216 -17094 -20092 -17065
rect -20216 -17150 -20182 -17094
rect -20126 -17150 -20092 -17094
rect -20216 -17179 -20092 -17150
rect -21624 -17790 -21500 -17761
rect -21624 -17846 -21590 -17790
rect -21534 -17846 -21500 -17790
rect -21624 -17875 -21500 -17846
rect -21628 -18910 -21504 -18881
rect -21628 -18966 -21594 -18910
rect -21538 -18966 -21504 -18910
rect -21628 -18995 -21504 -18966
rect -21488 -19030 -21410 -19014
rect -21520 -19118 -19992 -19110
rect -21520 -19182 -21494 -19118
rect -21430 -19182 -20082 -19118
rect -20018 -19182 -19992 -19118
rect -21520 -19190 -19992 -19182
rect -21624 -21150 -21500 -21121
rect -21624 -21206 -21590 -21150
rect -21534 -21206 -21500 -21150
rect -21624 -21235 -21500 -21206
rect -21520 -21358 -19992 -21350
rect -21520 -21422 -21494 -21358
rect -21430 -21422 -20082 -21358
rect -20018 -21422 -19992 -21358
rect -21520 -21430 -19992 -21422
rect -20212 -25630 -20088 -25601
rect -20212 -25686 -20178 -25630
rect -20122 -25686 -20088 -25630
rect -20212 -25715 -20088 -25686
rect -21520 -25838 -19992 -25830
rect -21520 -25902 -21494 -25838
rect -21430 -25902 -20082 -25838
rect -20018 -25902 -19992 -25838
rect -21520 -25910 -19992 -25902
rect -21624 -33470 -21500 -33441
rect -21624 -33526 -21590 -33470
rect -21534 -33526 -21500 -33470
rect -21624 -33555 -21500 -33526
rect -32920 -34590 -32796 -34561
rect -32920 -34646 -32886 -34590
rect -32830 -34646 -32796 -34590
rect -32920 -34675 -32796 -34646
rect -27272 -34590 -27148 -34561
rect -27272 -34646 -27238 -34590
rect -27182 -34646 -27148 -34590
rect -27272 -34675 -27148 -34646
rect -24448 -34590 -24324 -34561
rect -24448 -34646 -24414 -34590
rect -24358 -34646 -24324 -34590
rect -24448 -34675 -24324 -34646
rect -23036 -34590 -22912 -34561
rect -23036 -34646 -23002 -34590
rect -22946 -34646 -22912 -34590
rect -23036 -34675 -22912 -34646
rect -18800 -34590 -18676 -34561
rect -18800 -34646 -18766 -34590
rect -18710 -34646 -18676 -34590
rect -18800 -34675 -18676 -34646
rect -17388 -34589 -17264 -34560
rect -17388 -34645 -17354 -34589
rect -17298 -34645 -17264 -34589
rect -17388 -34674 -17264 -34645
rect -14556 -34594 -14440 -34569
rect -14556 -34650 -14526 -34594
rect -14470 -34650 -14440 -34594
rect -14556 -34675 -14440 -34650
rect -8908 -34594 -8792 -34569
rect -8908 -34650 -8878 -34594
rect -8822 -34650 -8792 -34594
rect -8908 -34675 -8792 -34650
<< via3 >>
rect -21494 -7982 -21430 -7918
rect -20082 -7982 -20018 -7918
rect -21494 -12462 -21430 -12398
rect -20082 -12462 -20018 -12398
rect -21494 -14702 -21430 -14638
rect -20082 -14702 -20018 -14638
rect -21494 -15822 -21430 -15758
rect -20082 -15822 -20018 -15758
rect -21494 -19182 -21430 -19118
rect -20082 -19182 -20018 -19118
rect -21494 -21422 -21430 -21358
rect -20082 -21422 -20018 -21358
rect -21494 -25902 -21430 -25838
rect -20082 -25902 -20018 -25838
<< metal4 >>
rect -43370 986 498 1082
rect -43370 -34318 -43274 986
rect -42690 -34794 -42594 878
rect -41958 -34318 -41862 986
rect -41278 -34794 -41182 878
rect -40546 -34318 -40450 986
rect -39866 -34794 -39770 878
rect -39134 -34318 -39038 986
rect -38454 -34794 -38358 878
rect -37722 -34318 -37626 986
rect -37042 -34794 -36946 878
rect -36310 -34318 -36214 986
rect -35630 -34794 -35534 878
rect -34898 -34318 -34802 986
rect -34218 -34794 -34122 878
rect -33486 -34318 -33390 986
rect -32806 -34794 -32710 878
rect -32074 -34318 -31978 986
rect -42690 -34890 -32710 -34794
rect -31394 -34794 -31298 878
rect -30662 -34318 -30566 986
rect -29982 -34794 -29886 878
rect -29250 -34318 -29154 986
rect -28570 -34794 -28474 878
rect -27838 -34318 -27742 986
rect -27158 -34794 -27062 878
rect -26426 -34318 -26330 986
rect -31394 -34890 -27062 -34794
rect -25746 -34794 -25650 878
rect -25014 -34318 -24918 986
rect -24334 -34794 -24238 878
rect -23602 -34318 -23506 986
rect -25746 -34890 -24238 -34794
rect -22922 -34890 -22826 878
rect -22190 -34318 -22094 986
rect -21510 -6962 -21414 439
rect -21510 -7909 -21414 -7818
rect -21511 -7918 -21413 -7909
rect -21511 -7982 -21494 -7918
rect -21430 -7982 -21413 -7918
rect -21511 -7991 -21413 -7982
rect -21510 -11442 -21414 -8420
rect -21510 -12389 -21414 -12298
rect -21511 -12398 -21413 -12389
rect -21511 -12462 -21494 -12398
rect -21430 -12462 -21413 -12398
rect -21511 -12471 -21413 -12462
rect -21510 -13689 -21414 -13332
rect -21510 -14629 -21414 -14538
rect -21511 -14638 -21413 -14629
rect -21511 -14702 -21494 -14638
rect -21430 -14702 -21413 -14638
rect -21511 -14711 -21413 -14702
rect -21510 -15749 -21414 -15658
rect -21511 -15758 -21413 -15749
rect -21511 -15822 -21494 -15758
rect -21430 -15822 -21413 -15758
rect -21511 -15831 -21413 -15822
rect -21510 -17046 -21414 -16702
rect -21510 -19109 -21414 -19018
rect -21511 -19118 -21413 -19109
rect -21511 -19182 -21494 -19118
rect -21430 -19182 -21413 -19118
rect -21511 -19191 -21413 -19182
rect -21510 -20418 -21414 -19979
rect -21510 -21349 -21414 -21258
rect -21511 -21358 -21413 -21349
rect -21511 -21422 -21494 -21358
rect -21430 -21422 -21413 -21358
rect -21511 -21431 -21413 -21422
rect -21510 -24891 -21414 -21864
rect -21510 -25829 -21414 -25738
rect -21511 -25838 -21413 -25829
rect -21511 -25902 -21494 -25838
rect -21430 -25902 -21413 -25838
rect -21511 -25911 -21413 -25902
rect -21510 -33842 -21414 -26331
rect -20778 -34318 -20682 986
rect -20098 -6962 -20002 148
rect -20098 -7909 -20002 -7818
rect -20099 -7918 -20001 -7909
rect -20099 -7982 -20082 -7918
rect -20018 -7982 -20001 -7918
rect -20099 -7991 -20001 -7982
rect -20098 -11442 -20002 -8451
rect -20098 -12389 -20002 -12298
rect -20099 -12398 -20001 -12389
rect -20099 -12462 -20082 -12398
rect -20018 -12462 -20001 -12398
rect -20099 -12471 -20001 -12462
rect -20098 -13682 -20002 -13323
rect -20098 -14629 -20002 -14538
rect -20099 -14638 -20001 -14629
rect -20099 -14702 -20082 -14638
rect -20018 -14702 -20001 -14638
rect -20099 -14711 -20001 -14702
rect -20098 -15749 -20002 -15658
rect -20099 -15758 -20001 -15749
rect -20099 -15822 -20082 -15758
rect -20018 -15822 -20001 -15758
rect -20099 -15831 -20001 -15822
rect -20098 -19109 -20002 -19018
rect -20099 -19118 -20001 -19109
rect -20099 -19182 -20082 -19118
rect -20018 -19182 -20001 -19118
rect -20099 -19191 -20001 -19182
rect -20098 -20402 -20002 -20096
rect -20098 -21349 -20002 -21258
rect -20099 -21358 -20001 -21349
rect -20099 -21422 -20082 -21358
rect -20018 -21422 -20001 -21358
rect -20099 -21431 -20001 -21422
rect -20098 -24898 -20002 -21857
rect -20098 -25829 -20002 -25738
rect -20099 -25838 -20001 -25829
rect -20099 -25902 -20082 -25838
rect -20018 -25902 -20001 -25838
rect -20099 -25911 -20001 -25902
rect -20098 -34553 -20002 -26858
rect -19366 -34316 -19270 986
rect -21510 -34794 -21414 -34698
rect -20098 -34794 -20002 -34698
rect -21510 -34890 -20002 -34794
rect -18686 -34888 -18590 880
rect -17954 -34318 -17858 986
rect -17274 -34794 -17178 878
rect -16542 -34318 -16446 986
rect -15862 -34794 -15766 878
rect -15130 -34318 -15034 986
rect -17274 -34890 -15766 -34794
rect -14450 -34794 -14354 878
rect -13718 -34318 -13622 986
rect -13038 -34794 -12942 878
rect -12306 -34318 -12210 986
rect -11626 -34794 -11530 878
rect -10894 -34318 -10798 986
rect -10214 -34794 -10118 878
rect -9482 -34318 -9386 986
rect -14450 -34890 -10118 -34794
rect -8802 -34794 -8706 878
rect -8070 -34318 -7974 986
rect -7390 -34794 -7294 878
rect -6658 -34318 -6562 986
rect -5978 -34794 -5882 878
rect -5246 -34318 -5150 986
rect -4566 -34794 -4470 878
rect -3834 -34318 -3738 986
rect -3154 -34794 -3058 878
rect -2422 -34318 -2326 986
rect -1742 -34794 -1646 878
rect -1010 -34318 -914 986
rect -330 -34794 -234 878
rect 402 -34318 498 986
rect 1082 -34794 1178 878
rect -8802 -34890 1178 -34794
use sky130_fd_pr__cap_mim_m3_1_8CZEMF  sky130_fd_pr__cap_mim_m3_1_8CZEMF_0
timestamp 1750100919
transform 1 0 -21290 0 1 -17470
box -23884 -18360 23884 18360
<< labels >>
flabel metal1 s -45174 -36038 -20206 -35934 0 FreeSans 1000 0 0 0 VCM
port 1 nsew
flabel metal1 s -45174 -36246 -21170 -36142 0 FreeSans 1000 0 0 0 SW[9]
port 2 nsew
flabel metal1 s -45174 -36454 -22478 -36350 0 FreeSans 1000 0 0 0 SW[8]
port 3 nsew
flabel metal1 s -45174 -36662 -21618 -36558 0 FreeSans 1000 0 0 0 SW[7]
port 4 nsew
flabel metal1 s -45174 -36870 -22686 -36766 0 FreeSans 1000 0 0 0 SW[6]
port 5 nsew
flabel metal1 s -45174 -37078 -19998 -36974 0 FreeSans 1000 0 0 0 SW[5]
port 6 nsew
flabel metal1 s -45174 -37286 -21410 -37182 0 FreeSans 1000 0 0 0 SW[4]
port 7 nsew
flabel metal1 s -45174 -37494 -18586 -37390 0 FreeSans 1000 0 0 0 SW[3]
port 8 nsew
flabel metal1 s -45174 -37702 -17174 -37598 0 FreeSans 1000 0 0 0 SW[2]
port 9 nsew
flabel metal1 s -45174 -37910 -28470 -37806 0 FreeSans 1000 0 0 0 SW[1]
port 10 nsew
flabel metal1 s -45174 -38118 -8702 -38014 0 FreeSans 1000 0 0 0 SW[0]
port 11 nsew
flabel metal4 s -21498 1009 -21442 1065 0 FreeSans 1000 0 0 0 VC
port 12 nsew
<< end >>
