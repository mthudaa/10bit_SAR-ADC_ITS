magic
tech sky130A
magscale 1 2
timestamp 1749497323
<< metal1 >>
rect -18696 -34606 -18686 -34586
rect -22932 -34710 -22922 -34606
rect -22826 -34631 -19679 -34606
rect -18957 -34631 -18686 -34606
rect -22826 -34682 -18686 -34631
rect -18590 -34606 -18580 -34586
rect -18590 -34682 -18450 -34606
rect -22826 -34710 -18450 -34682
rect -18346 -34710 -18336 -34606
rect -24344 -34923 -24334 -34819
rect -24238 -34923 -17274 -34819
rect -17070 -34923 -17060 -34819
rect -27168 -35131 -27158 -35027
rect -26954 -35131 -14450 -35027
rect -14354 -35131 -14344 -35027
rect -32816 -35338 -32806 -35234
rect -32710 -35338 -8802 -35234
rect -8598 -35338 -8588 -35234
rect -45174 -36038 -20206 -35934
rect -20102 -36038 2594 -35934
rect -45174 -36246 -21170 -36142
rect -21066 -36246 2594 -36142
rect -45174 -36454 -22478 -36350
rect -22374 -36454 2594 -36350
rect -45174 -36662 -21618 -36558
rect -21514 -36662 2594 -36558
rect -45174 -36870 -22686 -36766
rect -22582 -36870 2594 -36766
rect -45174 -37078 -19998 -36974
rect -19894 -37078 2594 -36974
rect -45174 -37286 -21410 -37182
rect -21306 -37286 2594 -37182
rect -45174 -37494 -18450 -37390
rect -18346 -37494 2594 -37390
rect -45174 -37702 -17174 -37598
rect -17070 -37702 2594 -37598
rect -45174 -37910 -27058 -37806
rect -26954 -37910 2594 -37806
rect -45174 -38118 -8702 -38014
rect -8598 -38118 2594 -38014
<< via1 >>
rect -22922 -34710 -22826 -34606
rect -18686 -34682 -18590 -34586
rect -18450 -34710 -18346 -34606
rect -24334 -34923 -24238 -34819
rect -17274 -34923 -17070 -34819
rect -27158 -35131 -26954 -35027
rect -14450 -35131 -14354 -35027
rect -32806 -35338 -32710 -35234
rect -8802 -35338 -8598 -35234
rect -20206 -36038 -20102 -35934
rect -21170 -36246 -21066 -36142
rect -22478 -36454 -22374 -36350
rect -21618 -36662 -21514 -36558
rect -22686 -36870 -22582 -36766
rect -19998 -37078 -19894 -36974
rect -21410 -37286 -21306 -37182
rect -18450 -37494 -18346 -37390
rect -17174 -37702 -17070 -37598
rect -27058 -37910 -26954 -37806
rect -8702 -38118 -8598 -38014
<< metal2 >>
rect -21410 -7716 -21306 -7706
rect -22686 -14436 -22582 -14426
rect -22686 -21156 -22582 -14550
rect -21618 -15566 -21514 -15556
rect -32806 -34586 -32710 -34576
rect -32806 -35234 -32710 -34682
rect -27158 -34586 -27062 -34576
rect -27158 -35017 -27062 -34682
rect -24334 -34586 -24238 -34576
rect -24334 -34819 -24238 -34682
rect -22922 -34586 -22826 -34576
rect -22922 -34720 -22826 -34710
rect -24334 -34933 -24238 -34923
rect -27158 -35027 -26954 -35017
rect -27158 -35141 -26954 -35131
rect -32806 -35348 -32710 -35338
rect -27058 -37806 -26954 -35141
rect -22686 -36766 -22582 -21270
rect -22478 -16926 -22374 -16916
rect -22478 -36350 -22374 -17030
rect -22478 -36464 -22374 -36454
rect -21618 -18926 -21514 -15670
rect -21618 -36558 -21514 -19030
rect -21618 -36672 -21514 -36662
rect -21410 -34606 -21306 -7830
rect -19998 -12196 -19894 -12186
rect -20206 -16686 -20102 -16676
rect -22686 -36880 -22582 -36870
rect -21410 -37182 -21306 -34710
rect -21170 -16926 -21066 -16916
rect -21170 -36142 -21066 -17030
rect -20206 -35934 -20102 -16790
rect -20206 -36048 -20102 -36038
rect -19998 -25646 -19894 -12310
rect -21170 -36256 -21066 -36246
rect -19998 -36974 -19894 -25750
rect -18686 -34586 -18590 -34576
rect -17274 -34586 -17178 -34576
rect -18686 -34692 -18590 -34682
rect -18450 -34606 -18346 -34596
rect -19998 -37088 -19894 -37078
rect -21410 -37296 -21306 -37286
rect -18450 -37390 -18346 -34710
rect -17274 -34809 -17178 -34682
rect -14450 -34586 -14354 -34576
rect -17274 -34819 -17070 -34809
rect -17274 -34933 -17070 -34923
rect -18450 -37504 -18346 -37494
rect -17174 -37598 -17070 -34933
rect -14450 -35027 -14354 -34682
rect -14450 -35141 -14354 -35131
rect -8802 -34586 -8706 -34576
rect -8802 -35224 -8706 -34682
rect -8802 -35234 -8598 -35224
rect -8802 -35348 -8598 -35338
rect -17174 -37712 -17070 -37702
rect -27058 -37920 -26954 -37910
rect -8702 -38014 -8598 -35348
rect -8702 -38128 -8598 -38118
<< via2 >>
rect -21410 -7830 -21306 -7716
rect -22686 -14550 -22582 -14436
rect -21618 -15670 -21514 -15566
rect -22686 -21270 -22582 -21156
rect -32806 -34682 -32710 -34586
rect -27158 -34682 -27062 -34586
rect -24334 -34682 -24238 -34586
rect -22922 -34606 -22826 -34586
rect -22922 -34682 -22826 -34606
rect -22478 -17030 -22374 -16926
rect -21618 -19030 -21514 -18926
rect -19998 -12310 -19894 -12196
rect -20206 -16790 -20102 -16686
rect -21410 -34710 -21306 -34606
rect -21170 -17030 -21066 -16926
rect -19998 -25750 -19894 -25646
rect -18686 -34682 -18590 -34586
rect -17274 -34682 -17178 -34586
rect -14450 -34682 -14354 -34586
rect -8802 -34682 -8706 -34586
<< metal3 >>
rect -21420 -7716 -21296 -7711
rect -21420 -7830 -21410 -7716
rect -21306 -7830 -21296 -7716
rect -21420 -7835 -21296 -7830
rect -21520 -7990 -21510 -7910
rect -21414 -7990 -20098 -7910
rect -20002 -7990 -19992 -7910
rect -20008 -12196 -19884 -12191
rect -20008 -12310 -19998 -12196
rect -19894 -12310 -19884 -12196
rect -20008 -12315 -19884 -12310
rect -21520 -12470 -21510 -12390
rect -21414 -12470 -20098 -12390
rect -20002 -12470 -19992 -12390
rect -22696 -14436 -22572 -14431
rect -22696 -14550 -22686 -14436
rect -22582 -14550 -22572 -14436
rect -22696 -14555 -22572 -14550
rect -21520 -14710 -21510 -14630
rect -21414 -14710 -20098 -14630
rect -20002 -14710 -19992 -14630
rect -21628 -15566 -21504 -15561
rect -21628 -15670 -21618 -15566
rect -21514 -15670 -21504 -15566
rect -21628 -15675 -21504 -15670
rect -21520 -15830 -21510 -15750
rect -21414 -15830 -20098 -15750
rect -20002 -15830 -19992 -15750
rect -20216 -16686 -20092 -16681
rect -20216 -16790 -20206 -16686
rect -20102 -16790 -20092 -16686
rect -20216 -16795 -20092 -16790
rect -22488 -16926 -22364 -16921
rect -22488 -17030 -22478 -16926
rect -22374 -17030 -22364 -16926
rect -22488 -17035 -22364 -17030
rect -21180 -16926 -21056 -16921
rect -21180 -17030 -21170 -16926
rect -21066 -17030 -21056 -16926
rect -21180 -17035 -21056 -17030
rect -21628 -18926 -21504 -18921
rect -21628 -19030 -21618 -18926
rect -21514 -19014 -21504 -18926
rect -21514 -19030 -21410 -19014
rect -21628 -19035 -21504 -19030
rect -21520 -19190 -21510 -19110
rect -21414 -19190 -20098 -19110
rect -20002 -19190 -19992 -19110
rect -22696 -21156 -22572 -21151
rect -22696 -21270 -22686 -21156
rect -22582 -21270 -22572 -21156
rect -22696 -21275 -22572 -21270
rect -21520 -21430 -21510 -21350
rect -21414 -21430 -20098 -21350
rect -20002 -21430 -19992 -21350
rect -20008 -25646 -19884 -25641
rect -20008 -25750 -19998 -25646
rect -19894 -25750 -19884 -25646
rect -20008 -25755 -19884 -25750
rect -21520 -25910 -21510 -25830
rect -21414 -25910 -20098 -25830
rect -20002 -25910 -19992 -25830
rect -32816 -34586 -32700 -34581
rect -32816 -34682 -32806 -34586
rect -32710 -34682 -32700 -34586
rect -32816 -34687 -32700 -34682
rect -27168 -34586 -27052 -34581
rect -27168 -34682 -27158 -34586
rect -27062 -34682 -27052 -34586
rect -27168 -34687 -27052 -34682
rect -24344 -34586 -24228 -34581
rect -24344 -34682 -24334 -34586
rect -24238 -34682 -24228 -34586
rect -24344 -34687 -24228 -34682
rect -22932 -34586 -22816 -34581
rect -22932 -34682 -22922 -34586
rect -22826 -34682 -22816 -34586
rect -18696 -34586 -18580 -34581
rect -22932 -34687 -22816 -34682
rect -21420 -34606 -21296 -34601
rect -21420 -34710 -21410 -34606
rect -21306 -34710 -21296 -34606
rect -18696 -34682 -18686 -34586
rect -18590 -34682 -18580 -34586
rect -18696 -34687 -18580 -34682
rect -17284 -34586 -17168 -34581
rect -17284 -34682 -17274 -34586
rect -17178 -34682 -17168 -34586
rect -17284 -34687 -17168 -34682
rect -14460 -34586 -14344 -34581
rect -14460 -34682 -14450 -34586
rect -14354 -34682 -14344 -34586
rect -14460 -34687 -14344 -34682
rect -8812 -34586 -8696 -34581
rect -8812 -34682 -8802 -34586
rect -8706 -34682 -8696 -34586
rect -8812 -34687 -8696 -34682
rect -21420 -34715 -21296 -34710
<< via3 >>
rect -21510 -7990 -21414 -7910
rect -20098 -7990 -20002 -7910
rect -21510 -12470 -21414 -12390
rect -20098 -12470 -20002 -12390
rect -21510 -14710 -21414 -14630
rect -20098 -14710 -20002 -14630
rect -21510 -15830 -21414 -15750
rect -20098 -15830 -20002 -15750
rect -21510 -19190 -21414 -19110
rect -20098 -19190 -20002 -19110
rect -21510 -21430 -21414 -21350
rect -20098 -21430 -20002 -21350
rect -21510 -25910 -21414 -25830
rect -20098 -25910 -20002 -25830
<< metal4 >>
rect -43370 986 498 1082
rect -43370 -34318 -43274 986
rect -42690 -34794 -42594 878
rect -41958 -34318 -41862 986
rect -41278 -34794 -41182 878
rect -40546 -34318 -40450 986
rect -39866 -34794 -39770 878
rect -39134 -34318 -39038 986
rect -38454 -34794 -38358 878
rect -37722 -34318 -37626 986
rect -37042 -34794 -36946 878
rect -36310 -34318 -36214 986
rect -35630 -34794 -35534 878
rect -34898 -34318 -34802 986
rect -34218 -34794 -34122 878
rect -33486 -34318 -33390 986
rect -32806 -34794 -32710 878
rect -32074 -34318 -31978 986
rect -42690 -34890 -32710 -34794
rect -31394 -34794 -31298 878
rect -30662 -34318 -30566 986
rect -29982 -34794 -29886 878
rect -29250 -34318 -29154 986
rect -28570 -34794 -28474 878
rect -27838 -34318 -27742 986
rect -27158 -34794 -27062 878
rect -26426 -34318 -26330 986
rect -31394 -34890 -27062 -34794
rect -25746 -34794 -25650 878
rect -25014 -34318 -24918 986
rect -24334 -34794 -24238 878
rect -23602 -34318 -23506 986
rect -25746 -34890 -24238 -34794
rect -22922 -34890 -22826 878
rect -22190 -34318 -22094 986
rect -21510 -6962 -21414 439
rect -21510 -7909 -21414 -7818
rect -21511 -7910 -21413 -7909
rect -21511 -7990 -21510 -7910
rect -21414 -7990 -21413 -7910
rect -21511 -7991 -21413 -7990
rect -21510 -11442 -21414 -8420
rect -21510 -12389 -21414 -12298
rect -21511 -12390 -21413 -12389
rect -21511 -12470 -21510 -12390
rect -21414 -12470 -21413 -12390
rect -21511 -12471 -21413 -12470
rect -21510 -13689 -21414 -13332
rect -21510 -14629 -21414 -14538
rect -21511 -14630 -21413 -14629
rect -21511 -14710 -21510 -14630
rect -21414 -14710 -21413 -14630
rect -21511 -14711 -21413 -14710
rect -21510 -15749 -21414 -15658
rect -21511 -15750 -21413 -15749
rect -21511 -15830 -21510 -15750
rect -21414 -15830 -21413 -15750
rect -21511 -15831 -21413 -15830
rect -21510 -17046 -21414 -16702
rect -21510 -19109 -21414 -19018
rect -21511 -19110 -21413 -19109
rect -21511 -19190 -21510 -19110
rect -21414 -19190 -21413 -19110
rect -21511 -19191 -21413 -19190
rect -21510 -20418 -21414 -19979
rect -21510 -21349 -21414 -21258
rect -21511 -21350 -21413 -21349
rect -21511 -21430 -21510 -21350
rect -21414 -21430 -21413 -21350
rect -21511 -21431 -21413 -21430
rect -21510 -24891 -21414 -21864
rect -21510 -25829 -21414 -25738
rect -21511 -25830 -21413 -25829
rect -21511 -25910 -21510 -25830
rect -21414 -25910 -21413 -25830
rect -21511 -25911 -21413 -25910
rect -21510 -33842 -21414 -26331
rect -20778 -34318 -20682 986
rect -20098 -6962 -20002 148
rect -20098 -7909 -20002 -7818
rect -20099 -7910 -20001 -7909
rect -20099 -7990 -20098 -7910
rect -20002 -7990 -20001 -7910
rect -20099 -7991 -20001 -7990
rect -20098 -11442 -20002 -8451
rect -20098 -12389 -20002 -12298
rect -20099 -12390 -20001 -12389
rect -20099 -12470 -20098 -12390
rect -20002 -12470 -20001 -12390
rect -20099 -12471 -20001 -12470
rect -20098 -13682 -20002 -13323
rect -20098 -14629 -20002 -14538
rect -20099 -14630 -20001 -14629
rect -20099 -14710 -20098 -14630
rect -20002 -14710 -20001 -14630
rect -20099 -14711 -20001 -14710
rect -20098 -15749 -20002 -15658
rect -20099 -15750 -20001 -15749
rect -20099 -15830 -20098 -15750
rect -20002 -15830 -20001 -15750
rect -20099 -15831 -20001 -15830
rect -20098 -19109 -20002 -19018
rect -20099 -19110 -20001 -19109
rect -20099 -19190 -20098 -19110
rect -20002 -19190 -20001 -19110
rect -20099 -19191 -20001 -19190
rect -20098 -20402 -20002 -20096
rect -20098 -21349 -20002 -21258
rect -20099 -21350 -20001 -21349
rect -20099 -21430 -20098 -21350
rect -20002 -21430 -20001 -21350
rect -20099 -21431 -20001 -21430
rect -20098 -24898 -20002 -21857
rect -20098 -25829 -20002 -25738
rect -20099 -25830 -20001 -25829
rect -20099 -25910 -20098 -25830
rect -20002 -25910 -20001 -25830
rect -20099 -25911 -20001 -25910
rect -20098 -34553 -20002 -26858
rect -19366 -34316 -19270 986
rect -21510 -34794 -21414 -34698
rect -20098 -34794 -20002 -34698
rect -21510 -34890 -20002 -34794
rect -18686 -34888 -18590 880
rect -17954 -34318 -17858 986
rect -17274 -34794 -17178 878
rect -16542 -34318 -16446 986
rect -15862 -34794 -15766 878
rect -15130 -34318 -15034 986
rect -17274 -34890 -15766 -34794
rect -14450 -34794 -14354 878
rect -13718 -34318 -13622 986
rect -13038 -34794 -12942 878
rect -12306 -34318 -12210 986
rect -11626 -34794 -11530 878
rect -10894 -34318 -10798 986
rect -10214 -34794 -10118 878
rect -9482 -34318 -9386 986
rect -14450 -34890 -10118 -34794
rect -8802 -34794 -8706 878
rect -8070 -34318 -7974 986
rect -7390 -34794 -7294 878
rect -6658 -34318 -6562 986
rect -5978 -34794 -5882 878
rect -5246 -34318 -5150 986
rect -4566 -34794 -4470 878
rect -3834 -34318 -3738 986
rect -3154 -34794 -3058 878
rect -2422 -34318 -2326 986
rect -1742 -34794 -1646 878
rect -1010 -34318 -914 986
rect -330 -34794 -234 878
rect 402 -34318 498 986
rect 1082 -34794 1178 878
rect -8802 -34890 1178 -34794
use sky130_fd_pr__cap_mim_m3_1_8CZEMF  sky130_fd_pr__cap_mim_m3_1_8CZEMF_0
timestamp 1748849030
transform 1 0 -21290 0 1 -17470
box -23884 -18360 23884 18360
<< labels >>
flabel metal1 -45174 -36038 -20206 -35934 0 FreeSans 800 0 0 0 VCM
port 0 nsew
flabel metal1 -45174 -36246 -21170 -36142 0 FreeSans 800 0 0 0 SW[9]
port 1 nsew
flabel metal1 -45174 -36454 -22478 -36350 0 FreeSans 800 0 0 0 SW[8]
port 2 nsew
flabel metal1 -45174 -36662 -21618 -36558 0 FreeSans 800 0 0 0 SW[7]
port 3 nsew
flabel metal1 -45174 -36870 -22686 -36766 0 FreeSans 800 0 0 0 SW[6]
port 4 nsew
flabel metal1 -45174 -37078 -19998 -36974 0 FreeSans 800 0 0 0 SW[5]
port 5 nsew
flabel metal1 -45174 -37286 -21410 -37182 0 FreeSans 800 0 0 0 SW[4]
port 6 nsew
flabel metal1 -45174 -37494 -18586 -37390 0 FreeSans 800 0 0 0 SW[3]
port 7 nsew
flabel metal1 -45174 -37702 -17174 -37598 0 FreeSans 800 0 0 0 SW[2]
port 8 nsew
flabel metal1 -45174 -37910 -28470 -37806 0 FreeSans 800 0 0 0 SW[1]
port 9 nsew
flabel metal1 -45174 -38118 -8702 -38014 0 FreeSans 800 0 0 0 SW[0]
port 10 nsew
flabel metal4 -21498 1009 -21442 1065 0 FreeSans 800 0 0 0 VC
port 11 nsew
<< end >>
