magic
tech sky130A
magscale 1 2
timestamp 1748851250
<< metal1 >>
rect -1094 -22194 -1084 -22090
rect -944 -22194 -38 -22090
rect 47481 -22194 48336 -22090
rect 48476 -22194 48486 -22090
rect 45426 -22402 45436 -22298
rect 45536 -22402 45546 -22298
rect 40620 -22610 40630 -22506
rect 40730 -22610 40740 -22506
rect 35818 -22818 35828 -22714
rect 35928 -22818 35938 -22714
rect 31016 -23026 31026 -22922
rect 31126 -23026 31136 -22922
rect 26219 -23234 26229 -23130
rect 26329 -23234 26339 -23130
rect 21412 -23442 21422 -23338
rect 21522 -23442 21532 -23338
rect 16612 -23650 16622 -23546
rect 16722 -23650 16732 -23546
rect 11808 -23858 11818 -23754
rect 11918 -23858 11928 -23754
rect 7006 -24066 7016 -23962
rect 7116 -24066 7126 -23962
rect 2204 -24274 2214 -24170
rect 2314 -24274 2324 -24170
rect 4128 -39935 4228 -39795
rect 4328 -39935 4428 -39595
rect 8930 -39935 9030 -39795
rect 9130 -39935 9230 -39595
rect 13732 -39935 13832 -39799
rect 13932 -39935 14032 -39595
rect 18534 -39935 18634 -39795
rect 18734 -39935 18834 -39595
rect 23336 -39935 23436 -39795
rect 23536 -39935 23636 -39595
rect 28138 -39935 28238 -39795
rect 28338 -39935 28438 -39595
rect 32940 -39935 33040 -39795
rect 33140 -39935 33240 -39595
rect 37742 -39935 37842 -39795
rect 37942 -39935 38042 -39595
rect 42544 -39935 42644 -39795
rect 42744 -39935 42844 -39595
rect 47346 -39935 47446 -39795
rect 47546 -39935 47646 -39595
<< via1 >>
rect -1084 -22194 -944 -22090
rect 48336 -22194 48476 -22090
rect 45436 -22402 45536 -22298
rect 40630 -22610 40730 -22506
rect 35828 -22818 35928 -22714
rect 31026 -23026 31126 -22922
rect 26229 -23234 26329 -23130
rect 21422 -23442 21522 -23338
rect 16622 -23650 16722 -23546
rect 11818 -23858 11918 -23754
rect 7016 -24066 7116 -23962
rect 2214 -24274 2314 -24170
<< metal2 >>
rect -1084 -22090 -944 -22080
rect 48336 -22090 48476 -22080
rect -1084 -39295 -944 -22194
rect -804 -38295 -664 -22090
rect -524 -38095 -384 -22090
rect 45436 -22298 45536 -22288
rect 40630 -22506 40730 -22496
rect 35828 -22714 35928 -22704
rect 31026 -22922 31126 -22912
rect 26229 -23130 26329 -23120
rect 21422 -23338 21522 -23328
rect 16622 -23546 16722 -23536
rect 11818 -23754 11918 -23744
rect 7016 -23962 7116 -23952
rect 2214 -24170 2314 -24160
rect 2214 -24514 2314 -24274
rect 7016 -25790 7116 -24066
rect 11818 -27066 11918 -23858
rect 16622 -28342 16722 -23650
rect 21422 -29618 21522 -23442
rect 26229 -30894 26329 -23234
rect 31026 -32170 31126 -23026
rect 35828 -33446 35928 -22818
rect 40630 -34722 40730 -22610
rect 45436 -35998 45536 -22402
rect 47776 -38095 47916 -22090
rect -524 -38195 -46 -38095
rect 47392 -38195 47916 -38095
rect 48056 -38295 48196 -22090
rect -804 -38395 -63 -38295
rect 47337 -38395 48196 -38295
rect 48336 -39295 48476 -22194
rect -1084 -39395 -129 -39295
rect 47347 -39395 48476 -39295
<< metal4 >>
rect 1308 15053 45802 15775
use cdac_sw_10b  cdac_sw_10b_0
timestamp 1748803925
transform 0 -1 4488 1 0 -39416
box -519 -43168 15012 4742
use x10b_cap_array  x10b_cap_array_0
timestamp 1748849030
transform 1 0 44991 0 1 13844
box -45174 -38128 2594 1931
<< labels >>
flabel metal2 -471 -38074 -431 -38034 0 FreeSans 800 0 0 0 VSS
port 0 nsew
flabel metal2 -756 -38069 -716 -38029 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel metal2 -1044 -38074 -1004 -38034 0 FreeSans 800 0 0 0 VCM
port 2 nsew
flabel metal4 21449 15318 21489 15358 0 FreeSans 800 0 0 0 VC
port 3 nsew
flabel metal1 4160 -39905 4200 -39865 0 FreeSans 800 0 0 0 SW_IN[0]
port 4 nsew
flabel metal1 8957 -39902 8997 -39862 0 FreeSans 800 0 0 0 SW_IN[1]
port 5 nsew
flabel metal1 13755 -39914 13795 -39874 0 FreeSans 800 0 0 0 SW_IN[2]
port 6 nsew
flabel metal1 18561 -39918 18601 -39878 0 FreeSans 800 0 0 0 SW_IN[3]
port 7 nsew
flabel metal1 23354 -39923 23394 -39883 0 FreeSans 800 0 0 0 SW_IN[4]
port 8 nsew
flabel metal1 28164 -39914 28204 -39874 0 FreeSans 800 0 0 0 SW_IN[5]
port 9 nsew
flabel metal1 32969 -39916 33009 -39876 0 FreeSans 800 0 0 0 SW_IN[6]
port 10 nsew
flabel metal1 37770 -39911 37810 -39871 0 FreeSans 800 0 0 0 SW_IN[7]
port 11 nsew
flabel metal1 42576 -39911 42616 -39871 0 FreeSans 800 0 0 0 SW_IN[8]
port 12 nsew
flabel metal1 47374 -39910 47414 -39870 0 FreeSans 800 0 0 0 SW_IN[9]
port 13 nsew
flabel metal1 4355 -39667 4395 -39627 0 FreeSans 800 0 0 0 CF[0]
port 14 nsew
flabel metal1 9157 -39658 9197 -39618 0 FreeSans 800 0 0 0 CF[1]
port 15 nsew
flabel metal1 13962 -39657 14002 -39617 0 FreeSans 800 0 0 0 CF[2]
port 16 nsew
flabel metal1 18760 -39671 18800 -39631 0 FreeSans 800 0 0 0 CF[3]
port 17 nsew
flabel metal1 23565 -39662 23605 -39622 0 FreeSans 800 0 0 0 CF[4]
port 18 nsew
flabel metal1 28367 -39661 28407 -39621 0 FreeSans 800 0 0 0 CF[5]
port 19 nsew
flabel metal1 33165 -39670 33205 -39630 0 FreeSans 800 0 0 0 CF[6]
port 20 nsew
flabel metal1 37970 -39663 38010 -39623 0 FreeSans 800 0 0 0 CF[7]
port 21 nsew
flabel metal1 42769 -39670 42809 -39630 0 FreeSans 800 0 0 0 CF[8]
port 22 nsew
flabel metal1 47575 -39663 47615 -39623 0 FreeSans 800 0 0 0 CF[9]
port 24 nsew
<< end >>
