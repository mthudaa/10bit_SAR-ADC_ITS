magic
tech sky130A
magscale 1 2
timestamp 1749574357
<< viali >>
rect 1855 25846 1889 25880
rect 3007 25846 3041 25880
rect 4159 25846 4193 25880
rect 5311 25846 5345 25880
rect 6463 25846 6497 25880
rect 7615 25846 7649 25880
rect 9055 25846 9089 25880
rect 9727 25846 9761 25880
rect 9823 25846 9857 25880
rect 2239 25772 2273 25806
rect 2143 25624 2177 25658
rect 2431 25624 2465 25658
rect 3199 25624 3233 25658
rect 4447 25624 4481 25658
rect 5503 25624 5537 25658
rect 6655 25624 6689 25658
rect 7807 25624 7841 25658
rect 9247 25624 9281 25658
rect 9439 25624 9473 25658
rect 10015 25624 10049 25658
rect 1951 25180 1985 25214
rect 10111 25180 10145 25214
rect 2239 24958 2273 24992
rect 9823 24958 9857 24992
rect 1663 24884 1697 24918
rect 1759 24884 1793 24918
rect 8479 23848 8513 23882
rect 9055 23848 9089 23882
rect 1855 23626 1889 23660
rect 6847 23626 6881 23660
rect 8767 23626 8801 23660
rect 6463 23552 6497 23586
rect 1567 23404 1601 23438
rect 5599 22960 5633 22994
rect 5983 22960 6017 22994
rect 7615 22960 7649 22994
rect 9823 22960 9857 22994
rect 8095 22886 8129 22920
rect 8287 22812 8321 22846
rect 7903 22738 7937 22772
rect 10111 22738 10145 22772
rect 9823 22516 9857 22550
rect 7807 22368 7841 22402
rect 1855 22294 1889 22328
rect 8191 22294 8225 22328
rect 1567 22072 1601 22106
rect 3583 21702 3617 21736
rect 3871 21702 3905 21736
rect 1951 21628 1985 21662
rect 4255 21628 4289 21662
rect 5983 21628 6017 21662
rect 1567 21554 1601 21588
rect 7807 21036 7841 21070
rect 8191 20962 8225 20996
rect 9823 20740 9857 20774
rect 1759 20518 1793 20552
rect 7423 20518 7457 20552
rect 5407 20370 5441 20404
rect 3295 20296 3329 20330
rect 3679 20296 3713 20330
rect 5791 20296 5825 20330
rect 9823 20296 9857 20330
rect 10111 20148 10145 20182
rect 1567 19852 1601 19886
rect 7807 19704 7841 19738
rect 1855 19630 1889 19664
rect 8191 19630 8225 19664
rect 9823 19408 9857 19442
rect 1759 19186 1793 19220
rect 5023 19038 5057 19072
rect 3295 18964 3329 18998
rect 3679 18964 3713 18998
rect 5407 18964 5441 18998
rect 7039 18742 7073 18776
rect 1567 18520 1601 18554
rect 7807 18372 7841 18406
rect 1855 18298 1889 18332
rect 8191 18298 8225 18332
rect 9727 18076 9761 18110
rect 1759 17854 1793 17888
rect 6463 17854 6497 17888
rect 10111 17780 10145 17814
rect 4447 17706 4481 17740
rect 3295 17632 3329 17666
rect 3679 17632 3713 17666
rect 4831 17632 4865 17666
rect 9823 17632 9857 17666
rect 1567 17188 1601 17222
rect 7807 17040 7841 17074
rect 1855 16966 1889 17000
rect 3967 16966 4001 17000
rect 8191 16966 8225 17000
rect 3583 16892 3617 16926
rect 5599 16744 5633 16778
rect 9823 16744 9857 16778
rect 1759 16522 1793 16556
rect 3295 16300 3329 16334
rect 3679 16226 3713 16260
rect 1567 15708 1601 15742
rect 2911 15708 2945 15742
rect 7519 15708 7553 15742
rect 1855 15634 1889 15668
rect 3295 15634 3329 15668
rect 7903 15634 7937 15668
rect 9823 15634 9857 15668
rect 4927 15412 4961 15446
rect 9535 15412 9569 15446
rect 10111 15412 10145 15446
rect 3295 14968 3329 15002
rect 3679 14894 3713 14928
rect 1663 14746 1697 14780
rect 7519 14376 7553 14410
rect 1855 14302 1889 14336
rect 4543 14302 4577 14336
rect 7903 14302 7937 14336
rect 1567 14228 1601 14262
rect 4159 14228 4193 14262
rect 6175 14080 6209 14114
rect 9535 14080 9569 14114
rect 5503 13636 5537 13670
rect 9823 13636 9857 13670
rect 5119 13562 5153 13596
rect 7135 13414 7169 13448
rect 10111 13414 10145 13448
rect 7807 13044 7841 13078
rect 1567 12970 1601 13004
rect 1759 12970 1793 13004
rect 3007 12970 3041 13004
rect 3391 12970 3425 13004
rect 5023 12970 5057 13004
rect 8191 12970 8225 13004
rect 9727 12748 9761 12782
rect 6175 12378 6209 12412
rect 1951 12304 1985 12338
rect 6559 12304 6593 12338
rect 1567 12230 1601 12264
rect 3583 12082 3617 12116
rect 8191 12082 8225 12116
rect 4447 11860 4481 11894
rect 1855 11638 1889 11672
rect 2815 11638 2849 11672
rect 6847 11638 6881 11672
rect 2431 11564 2465 11598
rect 6463 11564 6497 11598
rect 8479 11564 8513 11598
rect 1567 11416 1601 11450
rect 3487 11194 3521 11228
rect 1567 11046 1601 11080
rect 6271 11046 6305 11080
rect 1951 10972 1985 11006
rect 4255 10972 4289 11006
rect 6655 10972 6689 11006
rect 9823 10972 9857 11006
rect 3871 10898 3905 10932
rect 5887 10750 5921 10784
rect 8287 10750 8321 10784
rect 10111 10750 10145 10784
rect 4351 10528 4385 10562
rect 2335 10380 2369 10414
rect 7711 10380 7745 10414
rect 1855 10306 1889 10340
rect 2719 10306 2753 10340
rect 8095 10306 8129 10340
rect 1567 10084 1601 10118
rect 9727 10084 9761 10118
rect 7807 9048 7841 9082
rect 8191 8974 8225 9008
rect 1663 8900 1697 8934
rect 1759 8900 1793 8934
rect 9823 8752 9857 8786
rect 1759 8530 1793 8564
rect 7711 8308 7745 8342
rect 9823 8308 9857 8342
rect 10111 8308 10145 8342
rect 1663 8234 1697 8268
rect 3679 7864 3713 7898
rect 8191 7864 8225 7898
rect 1663 7716 1697 7750
rect 8095 7716 8129 7750
rect 2047 7642 2081 7676
rect 7135 7642 7169 7676
rect 7903 7568 7937 7602
rect 6847 7420 6881 7454
rect 1663 7198 1697 7232
rect 8191 7198 8225 7232
rect 6655 7050 6689 7084
rect 3295 6976 3329 7010
rect 6271 6976 6305 7010
rect 8575 6976 8609 7010
rect 3679 6902 3713 6936
rect 8773 6902 8807 6936
rect 7807 6828 7841 6862
rect 1759 6532 1793 6566
rect 6271 6532 6305 6566
rect 8191 6458 8225 6492
rect 5791 6384 5825 6418
rect 8863 6384 8897 6418
rect 3391 6310 3425 6344
rect 5311 6310 5345 6344
rect 6079 6310 6113 6344
rect 6559 6310 6593 6344
rect 8383 6310 8417 6344
rect 9055 6310 9089 6344
rect 9343 6310 9377 6344
rect 9823 6310 9857 6344
rect 3775 6236 3809 6270
rect 5599 6236 5633 6270
rect 6943 6236 6977 6270
rect 8095 6162 8129 6196
rect 8479 6162 8513 6196
rect 5503 6088 5537 6122
rect 9151 6088 9185 6122
rect 10111 6088 10145 6122
rect 9631 5792 9665 5826
rect 9535 5718 9569 5752
rect 1951 5644 1985 5678
rect 5599 5644 5633 5678
rect 6367 5644 6401 5678
rect 9343 5644 9377 5678
rect 9631 5644 9665 5678
rect 9727 5644 9761 5678
rect 1567 5570 1601 5604
rect 4831 5570 4865 5604
rect 5023 5570 5057 5604
rect 5119 5570 5153 5604
rect 5503 5570 5537 5604
rect 9247 5570 9281 5604
rect 9919 5570 9953 5604
rect 4927 5496 4961 5530
rect 3583 5422 3617 5456
rect 5791 5422 5825 5456
rect 9151 5422 9185 5456
rect 7999 5200 8033 5234
rect 9343 5200 9377 5234
rect 1663 5052 1697 5086
rect 6847 5052 6881 5086
rect 9055 5052 9089 5086
rect 9151 5052 9185 5086
rect 9439 5052 9473 5086
rect 2047 4978 2081 5012
rect 6175 4978 6209 5012
rect 6463 4978 6497 5012
rect 8575 4978 8609 5012
rect 9247 4978 9281 5012
rect 5791 4904 5825 4938
rect 3583 4756 3617 4790
rect 4639 4756 4673 4790
rect 8383 4756 8417 4790
rect 6175 4534 6209 4568
rect 8191 4534 8225 4568
rect 7039 4386 7073 4420
rect 3295 4312 3329 4346
rect 5695 4312 5729 4346
rect 5791 4312 5825 4346
rect 5983 4312 6017 4346
rect 6271 4312 6305 4346
rect 6463 4312 6497 4346
rect 6655 4312 6689 4346
rect 3679 4238 3713 4272
rect 8479 4238 8513 4272
rect 8671 4164 8705 4198
rect 1663 4090 1697 4124
rect 6367 4090 6401 4124
rect 8383 4090 8417 4124
rect 5887 3868 5921 3902
rect 6175 3868 6209 3902
rect 8095 3868 8129 3902
rect 2527 3794 2561 3828
rect 6079 3720 6113 3754
rect 6943 3720 6977 3754
rect 1567 3646 1601 3680
rect 6559 3646 6593 3680
rect 8383 3646 8417 3680
rect 9439 3646 9473 3680
rect 9823 3646 9857 3680
rect 10111 3572 10145 3606
rect 8191 3498 8225 3532
rect 9727 3424 9761 3458
rect 2623 3054 2657 3088
rect 2047 2980 2081 3014
rect 2527 2980 2561 3014
rect 2911 2980 2945 3014
rect 3295 2980 3329 3014
rect 4447 2980 4481 3014
rect 5503 2980 5537 3014
rect 6751 2980 6785 3014
rect 7135 2980 7169 3014
rect 9247 2980 9281 3014
rect 9535 2980 9569 3014
rect 10111 2980 10145 3014
rect 1855 2906 1889 2940
rect 3007 2906 3041 2940
rect 4159 2906 4193 2940
rect 5311 2906 5345 2940
rect 6463 2906 6497 2940
rect 9055 2906 9089 2940
rect 9727 2906 9761 2940
rect 9823 2906 9857 2940
rect 2239 2758 2273 2792
<< metal1 >>
rect 1152 26000 10560 26022
rect 1152 25948 1966 26000
rect 2018 25948 2030 26000
rect 2082 25948 2094 26000
rect 2146 25948 2158 26000
rect 2210 25948 2222 26000
rect 2274 25948 2286 26000
rect 2338 25948 7966 26000
rect 8018 25948 8030 26000
rect 8082 25948 8094 26000
rect 8146 25948 8158 26000
rect 8210 25948 8222 26000
rect 8274 25948 8286 26000
rect 8338 25948 10560 26000
rect 1152 25926 10560 25948
rect 1744 25837 1750 25889
rect 1802 25877 1808 25889
rect 1843 25880 1901 25886
rect 1843 25877 1855 25880
rect 1802 25849 1855 25877
rect 1802 25837 1808 25849
rect 1843 25846 1855 25849
rect 1889 25846 1901 25880
rect 1843 25840 1901 25846
rect 2992 25837 2998 25889
rect 3050 25837 3056 25889
rect 4144 25837 4150 25889
rect 4202 25837 4208 25889
rect 5296 25837 5302 25889
rect 5354 25837 5360 25889
rect 6448 25837 6454 25889
rect 6506 25837 6512 25889
rect 7600 25837 7606 25889
rect 7658 25837 7664 25889
rect 8656 25837 8662 25889
rect 8714 25877 8720 25889
rect 9043 25880 9101 25886
rect 9043 25877 9055 25880
rect 8714 25849 9055 25877
rect 8714 25837 8720 25849
rect 9043 25846 9055 25849
rect 9089 25846 9101 25880
rect 9043 25840 9101 25846
rect 9712 25837 9718 25889
rect 9770 25837 9776 25889
rect 9808 25837 9814 25889
rect 9866 25837 9872 25889
rect 1648 25763 1654 25815
rect 1706 25803 1712 25815
rect 2227 25806 2285 25812
rect 2227 25803 2239 25806
rect 1706 25775 2239 25803
rect 1706 25763 1712 25775
rect 2227 25772 2239 25775
rect 2273 25772 2285 25806
rect 2227 25766 2285 25772
rect 2131 25658 2189 25664
rect 2131 25624 2143 25658
rect 2177 25624 2189 25658
rect 2131 25618 2189 25624
rect 2146 25581 2174 25618
rect 2416 25615 2422 25667
rect 2474 25615 2480 25667
rect 3184 25615 3190 25667
rect 3242 25615 3248 25667
rect 4435 25658 4493 25664
rect 4435 25624 4447 25658
rect 4481 25624 4493 25658
rect 4435 25618 4493 25624
rect 2704 25581 2710 25593
rect 2146 25553 2710 25581
rect 2704 25541 2710 25553
rect 2762 25541 2768 25593
rect 4450 25581 4478 25618
rect 5488 25615 5494 25667
rect 5546 25615 5552 25667
rect 6448 25615 6454 25667
rect 6506 25655 6512 25667
rect 6643 25658 6701 25664
rect 6643 25655 6655 25658
rect 6506 25627 6655 25655
rect 6506 25615 6512 25627
rect 6643 25624 6655 25627
rect 6689 25624 6701 25658
rect 6643 25618 6701 25624
rect 7792 25615 7798 25667
rect 7850 25615 7856 25667
rect 7888 25615 7894 25667
rect 7946 25655 7952 25667
rect 9235 25658 9293 25664
rect 9235 25655 9247 25658
rect 7946 25627 9247 25655
rect 7946 25615 7952 25627
rect 9235 25624 9247 25627
rect 9281 25624 9293 25658
rect 9235 25618 9293 25624
rect 9424 25615 9430 25667
rect 9482 25615 9488 25667
rect 10003 25658 10061 25664
rect 10003 25624 10015 25658
rect 10049 25624 10061 25658
rect 10003 25618 10061 25624
rect 5680 25581 5686 25593
rect 4450 25553 5686 25581
rect 5680 25541 5686 25553
rect 5738 25541 5744 25593
rect 7600 25541 7606 25593
rect 7658 25581 7664 25593
rect 10018 25581 10046 25618
rect 7658 25553 10046 25581
rect 7658 25541 7664 25553
rect 1152 25334 10560 25356
rect 1152 25282 4966 25334
rect 5018 25282 5030 25334
rect 5082 25282 5094 25334
rect 5146 25282 5158 25334
rect 5210 25282 5222 25334
rect 5274 25282 5286 25334
rect 5338 25282 10560 25334
rect 1152 25260 10560 25282
rect 592 25171 598 25223
rect 650 25211 656 25223
rect 1939 25214 1997 25220
rect 1939 25211 1951 25214
rect 650 25183 1951 25211
rect 650 25171 656 25183
rect 1939 25180 1951 25183
rect 1985 25180 1997 25214
rect 1939 25174 1997 25180
rect 10099 25214 10157 25220
rect 10099 25180 10111 25214
rect 10145 25211 10157 25214
rect 10960 25211 10966 25223
rect 10145 25183 10966 25211
rect 10145 25180 10157 25183
rect 10099 25174 10157 25180
rect 10960 25171 10966 25183
rect 11018 25171 11024 25223
rect 2227 24992 2285 24998
rect 2227 24958 2239 24992
rect 2273 24989 2285 24992
rect 2512 24989 2518 25001
rect 2273 24961 2518 24989
rect 2273 24958 2285 24961
rect 2227 24952 2285 24958
rect 2512 24949 2518 24961
rect 2570 24949 2576 25001
rect 8464 24949 8470 25001
rect 8522 24989 8528 25001
rect 9811 24992 9869 24998
rect 9811 24989 9823 24992
rect 8522 24961 9823 24989
rect 8522 24949 8528 24961
rect 9811 24958 9823 24961
rect 9857 24958 9869 24992
rect 9811 24952 9869 24958
rect 880 24875 886 24927
rect 938 24915 944 24927
rect 1651 24918 1709 24924
rect 1651 24915 1663 24918
rect 938 24887 1663 24915
rect 938 24875 944 24887
rect 1651 24884 1663 24887
rect 1697 24884 1709 24918
rect 1651 24878 1709 24884
rect 1747 24918 1805 24924
rect 1747 24884 1759 24918
rect 1793 24915 1805 24918
rect 5584 24915 5590 24927
rect 1793 24887 5590 24915
rect 1793 24884 1805 24887
rect 1747 24878 1805 24884
rect 5584 24875 5590 24887
rect 5642 24875 5648 24927
rect 1152 24668 10560 24690
rect 1152 24616 1966 24668
rect 2018 24616 2030 24668
rect 2082 24616 2094 24668
rect 2146 24616 2158 24668
rect 2210 24616 2222 24668
rect 2274 24616 2286 24668
rect 2338 24616 7966 24668
rect 8018 24616 8030 24668
rect 8082 24616 8094 24668
rect 8146 24616 8158 24668
rect 8210 24616 8222 24668
rect 8274 24616 8286 24668
rect 8338 24616 10560 24668
rect 1152 24594 10560 24616
rect 1152 24002 10560 24024
rect 1152 23950 4966 24002
rect 5018 23950 5030 24002
rect 5082 23950 5094 24002
rect 5146 23950 5158 24002
rect 5210 23950 5222 24002
rect 5274 23950 5286 24002
rect 5338 23950 10560 24002
rect 1152 23928 10560 23950
rect 8464 23839 8470 23891
rect 8522 23839 8528 23891
rect 9043 23882 9101 23888
rect 9043 23848 9055 23882
rect 9089 23879 9101 23882
rect 9424 23879 9430 23891
rect 9089 23851 9430 23879
rect 9089 23848 9101 23851
rect 9043 23842 9101 23848
rect 9424 23839 9430 23851
rect 9482 23839 9488 23891
rect 1843 23660 1901 23666
rect 1843 23626 1855 23660
rect 1889 23657 1901 23660
rect 3856 23657 3862 23669
rect 1889 23629 3862 23657
rect 1889 23626 1901 23629
rect 1843 23620 1901 23626
rect 3856 23617 3862 23629
rect 3914 23617 3920 23669
rect 6736 23617 6742 23669
rect 6794 23657 6800 23669
rect 6835 23660 6893 23666
rect 6835 23657 6847 23660
rect 6794 23629 6847 23657
rect 6794 23617 6800 23629
rect 6835 23626 6847 23629
rect 6881 23626 6893 23660
rect 6835 23620 6893 23626
rect 8752 23617 8758 23669
rect 8810 23617 8816 23669
rect 5584 23543 5590 23595
rect 5642 23583 5648 23595
rect 6451 23586 6509 23592
rect 6451 23583 6463 23586
rect 5642 23555 6463 23583
rect 5642 23543 5648 23555
rect 6451 23552 6463 23555
rect 6497 23552 6509 23586
rect 6451 23546 6509 23552
rect 6064 23469 6070 23521
rect 6122 23509 6128 23521
rect 6658 23509 6686 23569
rect 6122 23481 6686 23509
rect 6122 23469 6128 23481
rect 784 23395 790 23447
rect 842 23435 848 23447
rect 1555 23438 1613 23444
rect 1555 23435 1567 23438
rect 842 23407 1567 23435
rect 842 23395 848 23407
rect 1555 23404 1567 23407
rect 1601 23404 1613 23438
rect 1555 23398 1613 23404
rect 1152 23336 10560 23358
rect 1152 23284 1966 23336
rect 2018 23284 2030 23336
rect 2082 23284 2094 23336
rect 2146 23284 2158 23336
rect 2210 23284 2222 23336
rect 2274 23284 2286 23336
rect 2338 23284 7966 23336
rect 8018 23284 8030 23336
rect 8082 23284 8094 23336
rect 8146 23284 8158 23336
rect 8210 23284 8222 23336
rect 8274 23284 8286 23336
rect 8338 23284 10560 23336
rect 1152 23262 10560 23284
rect 3856 23099 3862 23151
rect 3914 23139 3920 23151
rect 6736 23139 6742 23151
rect 3914 23111 6742 23139
rect 3914 23099 3920 23111
rect 6736 23099 6742 23111
rect 6794 23099 6800 23151
rect 6064 23025 6070 23077
rect 6122 23025 6128 23077
rect 5584 22951 5590 23003
rect 5642 22951 5648 23003
rect 5971 22994 6029 23000
rect 5971 22960 5983 22994
rect 6017 22960 6029 22994
rect 5971 22954 6029 22960
rect 5986 22917 6014 22954
rect 7600 22951 7606 23003
rect 7658 22951 7664 23003
rect 9808 22951 9814 23003
rect 9866 22951 9872 23003
rect 6544 22917 6550 22929
rect 5986 22889 6550 22917
rect 6544 22877 6550 22889
rect 6602 22877 6608 22929
rect 8083 22920 8141 22926
rect 8083 22886 8095 22920
rect 8129 22917 8141 22920
rect 8368 22917 8374 22929
rect 8129 22889 8374 22917
rect 8129 22886 8141 22889
rect 8083 22880 8141 22886
rect 8368 22877 8374 22889
rect 8426 22877 8432 22929
rect 8275 22846 8333 22852
rect 7186 22815 7934 22843
rect 6064 22729 6070 22781
rect 6122 22769 6128 22781
rect 7186 22769 7214 22815
rect 7906 22778 7934 22815
rect 8275 22812 8287 22846
rect 8321 22843 8333 22846
rect 8752 22843 8758 22855
rect 8321 22815 8758 22843
rect 8321 22812 8333 22815
rect 8275 22806 8333 22812
rect 8752 22803 8758 22815
rect 8810 22803 8816 22855
rect 6122 22741 7214 22769
rect 7891 22772 7949 22778
rect 6122 22729 6128 22741
rect 7891 22738 7903 22772
rect 7937 22738 7949 22772
rect 7891 22732 7949 22738
rect 10096 22729 10102 22781
rect 10154 22729 10160 22781
rect 1152 22670 10560 22692
rect 1152 22618 4966 22670
rect 5018 22618 5030 22670
rect 5082 22618 5094 22670
rect 5146 22618 5158 22670
rect 5210 22618 5222 22670
rect 5274 22618 5286 22670
rect 5338 22618 10560 22670
rect 1152 22596 10560 22618
rect 9808 22507 9814 22559
rect 9866 22507 9872 22559
rect 7795 22402 7853 22408
rect 7795 22368 7807 22402
rect 7841 22399 7853 22402
rect 8464 22399 8470 22411
rect 7841 22371 8470 22399
rect 7841 22368 7853 22371
rect 7795 22362 7853 22368
rect 8464 22359 8470 22371
rect 8522 22359 8528 22411
rect 1840 22285 1846 22337
rect 1898 22325 1904 22337
rect 6544 22325 6550 22337
rect 1898 22297 6550 22325
rect 1898 22285 1904 22297
rect 6544 22285 6550 22297
rect 6602 22285 6608 22337
rect 8179 22328 8237 22334
rect 8179 22294 8191 22328
rect 8225 22325 8237 22328
rect 8368 22325 8374 22337
rect 8225 22297 8374 22325
rect 8225 22294 8237 22297
rect 8179 22288 8237 22294
rect 8368 22285 8374 22297
rect 8426 22285 8432 22337
rect 8656 22211 8662 22263
rect 8714 22211 8720 22263
rect 880 22063 886 22115
rect 938 22103 944 22115
rect 1555 22106 1613 22112
rect 1555 22103 1567 22106
rect 938 22075 1567 22103
rect 938 22063 944 22075
rect 1555 22072 1567 22075
rect 1601 22072 1613 22106
rect 1555 22066 1613 22072
rect 1152 22004 10560 22026
rect 1152 21952 1966 22004
rect 2018 21952 2030 22004
rect 2082 21952 2094 22004
rect 2146 21952 2158 22004
rect 2210 21952 2222 22004
rect 2274 21952 2286 22004
rect 2338 21952 7966 22004
rect 8018 21952 8030 22004
rect 8082 21952 8094 22004
rect 8146 21952 8158 22004
rect 8210 21952 8222 22004
rect 8274 21952 8286 22004
rect 8338 21952 10560 22004
rect 1152 21930 10560 21952
rect 2434 21779 4094 21807
rect 2434 21745 2462 21779
rect 2416 21693 2422 21745
rect 2474 21693 2480 21745
rect 3571 21736 3629 21742
rect 3571 21702 3583 21736
rect 3617 21733 3629 21736
rect 3856 21733 3862 21745
rect 3617 21705 3862 21733
rect 3617 21702 3629 21705
rect 3571 21696 3629 21702
rect 3856 21693 3862 21705
rect 3914 21693 3920 21745
rect 4066 21719 4094 21779
rect 1939 21662 1997 21668
rect 1939 21628 1951 21662
rect 1985 21659 1997 21662
rect 3280 21659 3286 21671
rect 1985 21631 3286 21659
rect 1985 21628 1997 21631
rect 1939 21622 1997 21628
rect 3280 21619 3286 21631
rect 3338 21659 3344 21671
rect 4243 21662 4301 21668
rect 4243 21659 4255 21662
rect 3338 21631 4255 21659
rect 3338 21619 3344 21631
rect 4243 21628 4255 21631
rect 4289 21628 4301 21662
rect 4243 21622 4301 21628
rect 5971 21662 6029 21668
rect 5971 21628 5983 21662
rect 6017 21659 6029 21662
rect 8368 21659 8374 21671
rect 6017 21631 8374 21659
rect 6017 21628 6029 21631
rect 5971 21622 6029 21628
rect 8368 21619 8374 21631
rect 8426 21619 8432 21671
rect 1555 21588 1613 21594
rect 1555 21554 1567 21588
rect 1601 21585 1613 21588
rect 1840 21585 1846 21597
rect 1601 21557 1846 21585
rect 1601 21554 1613 21557
rect 1555 21548 1613 21554
rect 1840 21545 1846 21557
rect 1898 21545 1904 21597
rect 1152 21338 10560 21360
rect 1152 21286 4966 21338
rect 5018 21286 5030 21338
rect 5082 21286 5094 21338
rect 5146 21286 5158 21338
rect 5210 21286 5222 21338
rect 5274 21286 5286 21338
rect 5338 21286 10560 21338
rect 1152 21264 10560 21286
rect 7600 21027 7606 21079
rect 7658 21067 7664 21079
rect 7795 21070 7853 21076
rect 7795 21067 7807 21070
rect 7658 21039 7807 21067
rect 7658 21027 7664 21039
rect 7795 21036 7807 21039
rect 7841 21036 7853 21070
rect 7795 21030 7853 21036
rect 8179 20996 8237 21002
rect 8179 20962 8191 20996
rect 8225 20993 8237 20996
rect 8368 20993 8374 21005
rect 8225 20965 8374 20993
rect 8225 20962 8237 20965
rect 8179 20956 8237 20962
rect 8368 20953 8374 20965
rect 8426 20953 8432 21005
rect 8656 20879 8662 20931
rect 8714 20879 8720 20931
rect 9808 20731 9814 20783
rect 9866 20731 9872 20783
rect 1152 20672 10560 20694
rect 1152 20620 1966 20672
rect 2018 20620 2030 20672
rect 2082 20620 2094 20672
rect 2146 20620 2158 20672
rect 2210 20620 2222 20672
rect 2274 20620 2286 20672
rect 2338 20620 7966 20672
rect 8018 20620 8030 20672
rect 8082 20620 8094 20672
rect 8146 20620 8158 20672
rect 8210 20620 8222 20672
rect 8274 20620 8286 20672
rect 8338 20620 10560 20672
rect 1152 20598 10560 20620
rect 1747 20552 1805 20558
rect 1747 20518 1759 20552
rect 1793 20549 1805 20552
rect 1840 20549 1846 20561
rect 1793 20521 1846 20549
rect 1793 20518 1805 20521
rect 1747 20512 1805 20518
rect 1840 20509 1846 20521
rect 1898 20509 1904 20561
rect 5584 20509 5590 20561
rect 5642 20509 5648 20561
rect 7411 20552 7469 20558
rect 7411 20518 7423 20552
rect 7457 20549 7469 20552
rect 7888 20549 7894 20561
rect 7457 20521 7894 20549
rect 7457 20518 7469 20521
rect 7411 20512 7469 20518
rect 7888 20509 7894 20521
rect 7946 20509 7952 20561
rect 5602 20475 5630 20509
rect 5410 20447 5630 20475
rect 5410 20413 5438 20447
rect 2416 20361 2422 20413
rect 2474 20361 2480 20413
rect 5392 20361 5398 20413
rect 5450 20361 5456 20413
rect 6064 20361 6070 20413
rect 6122 20361 6128 20413
rect 3280 20287 3286 20339
rect 3338 20287 3344 20339
rect 3664 20287 3670 20339
rect 3722 20327 3728 20339
rect 5779 20330 5837 20336
rect 5779 20327 5791 20330
rect 3722 20299 5791 20327
rect 3722 20287 3728 20299
rect 5779 20296 5791 20299
rect 5825 20327 5837 20330
rect 5872 20327 5878 20339
rect 5825 20299 5878 20327
rect 5825 20296 5837 20299
rect 5779 20290 5837 20296
rect 5872 20287 5878 20299
rect 5930 20287 5936 20339
rect 9808 20287 9814 20339
rect 9866 20287 9872 20339
rect 10096 20139 10102 20191
rect 10154 20139 10160 20191
rect 1152 20006 10560 20028
rect 1152 19954 4966 20006
rect 5018 19954 5030 20006
rect 5082 19954 5094 20006
rect 5146 19954 5158 20006
rect 5210 19954 5222 20006
rect 5274 19954 5286 20006
rect 5338 19954 10560 20006
rect 1152 19932 10560 19954
rect 1552 19843 1558 19895
rect 1610 19843 1616 19895
rect 7795 19738 7853 19744
rect 7795 19704 7807 19738
rect 7841 19735 7853 19738
rect 7888 19735 7894 19747
rect 7841 19707 7894 19735
rect 7841 19704 7853 19707
rect 7795 19698 7853 19704
rect 7888 19695 7894 19707
rect 7946 19695 7952 19747
rect 1744 19621 1750 19673
rect 1802 19661 1808 19673
rect 1843 19664 1901 19670
rect 1843 19661 1855 19664
rect 1802 19633 1855 19661
rect 1802 19621 1808 19633
rect 1843 19630 1855 19633
rect 1889 19661 1901 19664
rect 3664 19661 3670 19673
rect 1889 19633 3670 19661
rect 1889 19630 1901 19633
rect 1843 19624 1901 19630
rect 3664 19621 3670 19633
rect 3722 19621 3728 19673
rect 8179 19664 8237 19670
rect 8179 19661 8191 19664
rect 7906 19633 8191 19661
rect 7906 19599 7934 19633
rect 8179 19630 8191 19633
rect 8225 19661 8237 19664
rect 8368 19661 8374 19673
rect 8225 19633 8374 19661
rect 8225 19630 8237 19633
rect 8179 19624 8237 19630
rect 8368 19621 8374 19633
rect 8426 19621 8432 19673
rect 7888 19547 7894 19599
rect 7946 19547 7952 19599
rect 8656 19547 8662 19599
rect 8714 19547 8720 19599
rect 9808 19399 9814 19451
rect 9866 19399 9872 19451
rect 1152 19340 10560 19362
rect 1152 19288 1966 19340
rect 2018 19288 2030 19340
rect 2082 19288 2094 19340
rect 2146 19288 2158 19340
rect 2210 19288 2222 19340
rect 2274 19288 2286 19340
rect 2338 19288 7966 19340
rect 8018 19288 8030 19340
rect 8082 19288 8094 19340
rect 8146 19288 8158 19340
rect 8210 19288 8222 19340
rect 8274 19288 8286 19340
rect 8338 19288 10560 19340
rect 1152 19266 10560 19288
rect 1744 19177 1750 19229
rect 1802 19177 1808 19229
rect 5392 19143 5398 19155
rect 5026 19115 5398 19143
rect 2416 19029 2422 19081
rect 2474 19029 2480 19081
rect 4432 19029 4438 19081
rect 4490 19069 4496 19081
rect 5026 19078 5054 19115
rect 5392 19103 5398 19115
rect 5450 19103 5456 19155
rect 6064 19143 6070 19155
rect 5602 19115 6070 19143
rect 5602 19081 5630 19115
rect 6064 19103 6070 19115
rect 6122 19103 6128 19155
rect 5011 19072 5069 19078
rect 5011 19069 5023 19072
rect 4490 19041 5023 19069
rect 4490 19029 4496 19041
rect 5011 19038 5023 19041
rect 5057 19038 5069 19072
rect 5011 19032 5069 19038
rect 5584 19029 5590 19081
rect 5642 19029 5648 19081
rect 3280 18955 3286 19007
rect 3338 18955 3344 19007
rect 3667 18998 3725 19004
rect 3667 18964 3679 18998
rect 3713 18995 3725 18998
rect 4144 18995 4150 19007
rect 3713 18967 4150 18995
rect 3713 18964 3725 18967
rect 3667 18958 3725 18964
rect 4144 18955 4150 18967
rect 4202 18995 4208 19007
rect 5395 18998 5453 19004
rect 5395 18995 5407 18998
rect 4202 18967 5407 18995
rect 4202 18955 4208 18967
rect 5395 18964 5407 18967
rect 5441 18964 5453 18998
rect 5395 18958 5453 18964
rect 7027 18776 7085 18782
rect 7027 18742 7039 18776
rect 7073 18773 7085 18776
rect 7792 18773 7798 18785
rect 7073 18745 7798 18773
rect 7073 18742 7085 18745
rect 7027 18736 7085 18742
rect 7792 18733 7798 18745
rect 7850 18733 7856 18785
rect 1152 18674 10560 18696
rect 1152 18622 4966 18674
rect 5018 18622 5030 18674
rect 5082 18622 5094 18674
rect 5146 18622 5158 18674
rect 5210 18622 5222 18674
rect 5274 18622 5286 18674
rect 5338 18622 10560 18674
rect 1152 18600 10560 18622
rect 1552 18511 1558 18563
rect 1610 18511 1616 18563
rect 6448 18363 6454 18415
rect 6506 18403 6512 18415
rect 7795 18406 7853 18412
rect 7795 18403 7807 18406
rect 6506 18375 7807 18403
rect 6506 18363 6512 18375
rect 7795 18372 7807 18375
rect 7841 18372 7853 18406
rect 7795 18366 7853 18372
rect 1744 18289 1750 18341
rect 1802 18329 1808 18341
rect 1843 18332 1901 18338
rect 1843 18329 1855 18332
rect 1802 18301 1855 18329
rect 1802 18289 1808 18301
rect 1843 18298 1855 18301
rect 1889 18329 1901 18332
rect 4144 18329 4150 18341
rect 1889 18301 4150 18329
rect 1889 18298 1901 18301
rect 1843 18292 1901 18298
rect 4144 18289 4150 18301
rect 4202 18289 4208 18341
rect 7888 18289 7894 18341
rect 7946 18329 7952 18341
rect 8179 18332 8237 18338
rect 8179 18329 8191 18332
rect 7946 18301 8191 18329
rect 7946 18289 7952 18301
rect 8179 18298 8191 18301
rect 8225 18298 8237 18332
rect 8179 18292 8237 18298
rect 8656 18215 8662 18267
rect 8714 18215 8720 18267
rect 9712 18067 9718 18119
rect 9770 18067 9776 18119
rect 1152 18008 10560 18030
rect 1152 17956 1966 18008
rect 2018 17956 2030 18008
rect 2082 17956 2094 18008
rect 2146 17956 2158 18008
rect 2210 17956 2222 18008
rect 2274 17956 2286 18008
rect 2338 17956 7966 18008
rect 8018 17956 8030 18008
rect 8082 17956 8094 18008
rect 8146 17956 8158 18008
rect 8210 17956 8222 18008
rect 8274 17956 8286 18008
rect 8338 17956 10560 18008
rect 1152 17934 10560 17956
rect 1744 17845 1750 17897
rect 1802 17845 1808 17897
rect 6448 17845 6454 17897
rect 6506 17845 6512 17897
rect 5584 17811 5590 17823
rect 2818 17783 5590 17811
rect 2416 17697 2422 17749
rect 2474 17697 2480 17749
rect 2434 17663 2462 17697
rect 2818 17675 2846 17783
rect 4432 17697 4438 17749
rect 4490 17697 4496 17749
rect 4642 17723 4670 17783
rect 5584 17771 5590 17783
rect 5642 17771 5648 17823
rect 10096 17771 10102 17823
rect 10154 17771 10160 17823
rect 2800 17663 2806 17675
rect 2434 17635 2806 17663
rect 2800 17623 2806 17635
rect 2858 17623 2864 17675
rect 3280 17623 3286 17675
rect 3338 17623 3344 17675
rect 3667 17666 3725 17672
rect 3667 17632 3679 17666
rect 3713 17663 3725 17666
rect 4240 17663 4246 17675
rect 3713 17635 4246 17663
rect 3713 17632 3725 17635
rect 3667 17626 3725 17632
rect 4240 17623 4246 17635
rect 4298 17663 4304 17675
rect 4819 17666 4877 17672
rect 4819 17663 4831 17666
rect 4298 17635 4831 17663
rect 4298 17623 4304 17635
rect 4819 17632 4831 17635
rect 4865 17632 4877 17666
rect 4819 17626 4877 17632
rect 9808 17623 9814 17675
rect 9866 17623 9872 17675
rect 1152 17342 10560 17364
rect 1152 17290 4966 17342
rect 5018 17290 5030 17342
rect 5082 17290 5094 17342
rect 5146 17290 5158 17342
rect 5210 17290 5222 17342
rect 5274 17290 5286 17342
rect 5338 17290 10560 17342
rect 1152 17268 10560 17290
rect 1264 17179 1270 17231
rect 1322 17219 1328 17231
rect 1555 17222 1613 17228
rect 1555 17219 1567 17222
rect 1322 17191 1567 17219
rect 1322 17179 1328 17191
rect 1555 17188 1567 17191
rect 1601 17188 1613 17222
rect 1555 17182 1613 17188
rect 4240 17071 4246 17083
rect 1858 17043 4246 17071
rect 1744 16957 1750 17009
rect 1802 16997 1808 17009
rect 1858 17006 1886 17043
rect 4240 17031 4246 17043
rect 4298 17031 4304 17083
rect 7792 17031 7798 17083
rect 7850 17031 7856 17083
rect 1843 17000 1901 17006
rect 1843 16997 1855 17000
rect 1802 16969 1855 16997
rect 1802 16957 1808 16969
rect 1843 16966 1855 16969
rect 1889 16966 1901 17000
rect 1843 16960 1901 16966
rect 3952 16957 3958 17009
rect 4010 16957 4016 17009
rect 7888 16957 7894 17009
rect 7946 16997 7952 17009
rect 8179 17000 8237 17006
rect 8179 16997 8191 17000
rect 7946 16969 8191 16997
rect 7946 16957 7952 16969
rect 8179 16966 8191 16969
rect 8225 16966 8237 17000
rect 8179 16960 8237 16966
rect 8758 16935 8810 16941
rect 3571 16926 3629 16932
rect 3571 16892 3583 16926
rect 3617 16892 3629 16926
rect 5584 16923 5590 16935
rect 5136 16895 5590 16923
rect 3571 16886 3629 16892
rect 2896 16809 2902 16861
rect 2954 16849 2960 16861
rect 3586 16849 3614 16886
rect 5584 16883 5590 16895
rect 5642 16883 5648 16935
rect 8758 16877 8810 16883
rect 4432 16849 4438 16861
rect 2954 16821 4438 16849
rect 2954 16809 2960 16821
rect 4432 16809 4438 16821
rect 4490 16809 4496 16861
rect 5584 16735 5590 16787
rect 5642 16735 5648 16787
rect 9808 16735 9814 16787
rect 9866 16735 9872 16787
rect 1152 16676 10560 16698
rect 1152 16624 1966 16676
rect 2018 16624 2030 16676
rect 2082 16624 2094 16676
rect 2146 16624 2158 16676
rect 2210 16624 2222 16676
rect 2274 16624 2286 16676
rect 2338 16624 7966 16676
rect 8018 16624 8030 16676
rect 8082 16624 8094 16676
rect 8146 16624 8158 16676
rect 8210 16624 8222 16676
rect 8274 16624 8286 16676
rect 8338 16624 10560 16676
rect 1152 16602 10560 16624
rect 1744 16513 1750 16565
rect 1802 16513 1808 16565
rect 2800 16365 2806 16417
rect 2858 16365 2864 16417
rect 3280 16291 3286 16343
rect 3338 16291 3344 16343
rect 2992 16217 2998 16269
rect 3050 16257 3056 16269
rect 3667 16260 3725 16266
rect 3667 16257 3679 16260
rect 3050 16229 3679 16257
rect 3050 16217 3056 16229
rect 3667 16226 3679 16229
rect 3713 16257 3725 16260
rect 3952 16257 3958 16269
rect 3713 16229 3958 16257
rect 3713 16226 3725 16229
rect 3667 16220 3725 16226
rect 3952 16217 3958 16229
rect 4010 16217 4016 16269
rect 1152 16010 10560 16032
rect 1152 15958 4966 16010
rect 5018 15958 5030 16010
rect 5082 15958 5094 16010
rect 5146 15958 5158 16010
rect 5210 15958 5222 16010
rect 5274 15958 5286 16010
rect 5338 15958 10560 16010
rect 1152 15936 10560 15958
rect 784 15699 790 15751
rect 842 15739 848 15751
rect 1555 15742 1613 15748
rect 1555 15739 1567 15742
rect 842 15711 1567 15739
rect 842 15699 848 15711
rect 1555 15708 1567 15711
rect 1601 15708 1613 15742
rect 1555 15702 1613 15708
rect 2896 15699 2902 15751
rect 2954 15699 2960 15751
rect 5584 15699 5590 15751
rect 5642 15739 5648 15751
rect 7507 15742 7565 15748
rect 7507 15739 7519 15742
rect 5642 15711 7519 15739
rect 5642 15699 5648 15711
rect 7507 15708 7519 15711
rect 7553 15708 7565 15742
rect 7507 15702 7565 15708
rect 1843 15668 1901 15674
rect 1843 15634 1855 15668
rect 1889 15665 1901 15668
rect 2992 15665 2998 15677
rect 1889 15637 2998 15665
rect 1889 15634 1901 15637
rect 1843 15628 1901 15634
rect 2992 15625 2998 15637
rect 3050 15625 3056 15677
rect 3283 15668 3341 15674
rect 3283 15634 3295 15668
rect 3329 15665 3341 15668
rect 3664 15665 3670 15677
rect 3329 15637 3670 15665
rect 3329 15634 3341 15637
rect 3283 15628 3341 15634
rect 3664 15625 3670 15637
rect 3722 15625 3728 15677
rect 7888 15625 7894 15677
rect 7946 15625 7952 15677
rect 9808 15625 9814 15677
rect 9866 15625 9872 15677
rect 2800 15551 2806 15603
rect 2858 15591 2864 15603
rect 2858 15563 3120 15591
rect 2858 15551 2864 15563
rect 8752 15551 8758 15603
rect 8810 15551 8816 15603
rect 4915 15446 4973 15452
rect 4915 15412 4927 15446
rect 4961 15443 4973 15446
rect 5392 15443 5398 15455
rect 4961 15415 5398 15443
rect 4961 15412 4973 15415
rect 4915 15406 4973 15412
rect 5392 15403 5398 15415
rect 5450 15443 5456 15455
rect 5680 15443 5686 15455
rect 5450 15415 5686 15443
rect 5450 15403 5456 15415
rect 5680 15403 5686 15415
rect 5738 15403 5744 15455
rect 9523 15446 9581 15452
rect 9523 15412 9535 15446
rect 9569 15443 9581 15446
rect 9808 15443 9814 15455
rect 9569 15415 9814 15443
rect 9569 15412 9581 15415
rect 9523 15406 9581 15412
rect 9808 15403 9814 15415
rect 9866 15403 9872 15455
rect 10096 15403 10102 15455
rect 10154 15403 10160 15455
rect 1152 15344 10560 15366
rect 1152 15292 1966 15344
rect 2018 15292 2030 15344
rect 2082 15292 2094 15344
rect 2146 15292 2158 15344
rect 2210 15292 2222 15344
rect 2274 15292 2286 15344
rect 2338 15292 7966 15344
rect 8018 15292 8030 15344
rect 8082 15292 8094 15344
rect 8146 15292 8158 15344
rect 8210 15292 8222 15344
rect 8274 15292 8286 15344
rect 8338 15292 10560 15344
rect 1152 15270 10560 15292
rect 2800 15033 2806 15085
rect 2858 15033 2864 15085
rect 3280 14959 3286 15011
rect 3338 14959 3344 15011
rect 3664 14885 3670 14937
rect 3722 14885 3728 14937
rect 1651 14780 1709 14786
rect 1651 14746 1663 14780
rect 1697 14777 1709 14780
rect 2992 14777 2998 14789
rect 1697 14749 2998 14777
rect 1697 14746 1709 14749
rect 1651 14740 1709 14746
rect 2992 14737 2998 14749
rect 3050 14777 3056 14789
rect 3376 14777 3382 14789
rect 3050 14749 3382 14777
rect 3050 14737 3056 14749
rect 3376 14737 3382 14749
rect 3434 14737 3440 14789
rect 1152 14678 10560 14700
rect 1152 14626 4966 14678
rect 5018 14626 5030 14678
rect 5082 14626 5094 14678
rect 5146 14626 5158 14678
rect 5210 14626 5222 14678
rect 5274 14626 5286 14678
rect 5338 14626 10560 14678
rect 1152 14604 10560 14626
rect 2800 14441 2806 14493
rect 2858 14481 2864 14493
rect 2858 14453 4286 14481
rect 2858 14441 2864 14453
rect 4258 14407 4286 14453
rect 5392 14441 5398 14493
rect 5450 14481 5456 14493
rect 5450 14453 7550 14481
rect 5450 14441 5456 14453
rect 7522 14416 7550 14453
rect 7507 14410 7565 14416
rect 4258 14379 4670 14407
rect 1843 14336 1901 14342
rect 1843 14302 1855 14336
rect 1889 14333 1901 14336
rect 3664 14333 3670 14345
rect 1889 14305 3670 14333
rect 1889 14302 1901 14305
rect 1843 14296 1901 14302
rect 3664 14293 3670 14305
rect 3722 14293 3728 14345
rect 4240 14293 4246 14345
rect 4298 14333 4304 14345
rect 4531 14336 4589 14342
rect 4531 14333 4543 14336
rect 4298 14305 4543 14333
rect 4298 14293 4304 14305
rect 4531 14302 4543 14305
rect 4577 14302 4589 14336
rect 4531 14296 4589 14302
rect 4642 14271 4670 14379
rect 7507 14376 7519 14410
rect 7553 14376 7565 14410
rect 7507 14370 7565 14376
rect 7888 14293 7894 14345
rect 7946 14333 7952 14345
rect 8368 14333 8374 14345
rect 7946 14305 8374 14333
rect 7946 14293 7952 14305
rect 8368 14293 8374 14305
rect 8426 14293 8432 14345
rect 784 14219 790 14271
rect 842 14259 848 14271
rect 1555 14262 1613 14268
rect 1555 14259 1567 14262
rect 842 14231 1567 14259
rect 842 14219 848 14231
rect 1555 14228 1567 14231
rect 1601 14228 1613 14262
rect 1555 14222 1613 14228
rect 2896 14219 2902 14271
rect 2954 14259 2960 14271
rect 4147 14262 4205 14268
rect 4147 14259 4159 14262
rect 2954 14231 4159 14259
rect 2954 14219 2960 14231
rect 4147 14228 4159 14231
rect 4193 14228 4205 14262
rect 4147 14222 4205 14228
rect 4624 14219 4630 14271
rect 4682 14219 4688 14271
rect 8752 14219 8758 14271
rect 8810 14219 8816 14271
rect 6163 14114 6221 14120
rect 6163 14080 6175 14114
rect 6209 14111 6221 14114
rect 7024 14111 7030 14123
rect 6209 14083 7030 14111
rect 6209 14080 6221 14083
rect 6163 14074 6221 14080
rect 7024 14071 7030 14083
rect 7082 14071 7088 14123
rect 9520 14071 9526 14123
rect 9578 14071 9584 14123
rect 1152 14012 10560 14034
rect 1152 13960 1966 14012
rect 2018 13960 2030 14012
rect 2082 13960 2094 14012
rect 2146 13960 2158 14012
rect 2210 13960 2222 14012
rect 2274 13960 2286 14012
rect 2338 13960 7966 14012
rect 8018 13960 8030 14012
rect 8082 13960 8094 14012
rect 8146 13960 8158 14012
rect 8210 13960 8222 14012
rect 8274 13960 8286 14012
rect 8338 13960 10560 14012
rect 1152 13938 10560 13960
rect 7216 13815 7222 13827
rect 5314 13787 7222 13815
rect 4624 13701 4630 13753
rect 4682 13741 4688 13753
rect 5314 13741 5342 13787
rect 7216 13775 7222 13787
rect 7274 13775 7280 13827
rect 4682 13727 5342 13741
rect 4682 13713 5328 13727
rect 4682 13701 4688 13713
rect 4144 13627 4150 13679
rect 4202 13667 4208 13679
rect 5491 13670 5549 13676
rect 5491 13667 5503 13670
rect 4202 13639 5503 13667
rect 4202 13627 4208 13639
rect 5491 13636 5503 13639
rect 5537 13636 5549 13670
rect 5491 13630 5549 13636
rect 9712 13627 9718 13679
rect 9770 13667 9776 13679
rect 9811 13670 9869 13676
rect 9811 13667 9823 13670
rect 9770 13639 9823 13667
rect 9770 13627 9776 13639
rect 9811 13636 9823 13639
rect 9857 13636 9869 13670
rect 9811 13630 9869 13636
rect 2896 13553 2902 13605
rect 2954 13593 2960 13605
rect 5107 13596 5165 13602
rect 5107 13593 5119 13596
rect 2954 13565 5119 13593
rect 2954 13553 2960 13565
rect 5107 13562 5119 13565
rect 5153 13593 5165 13596
rect 6160 13593 6166 13605
rect 5153 13565 6166 13593
rect 5153 13562 5165 13565
rect 5107 13556 5165 13562
rect 6160 13553 6166 13565
rect 6218 13553 6224 13605
rect 7123 13448 7181 13454
rect 7123 13414 7135 13448
rect 7169 13445 7181 13448
rect 7504 13445 7510 13457
rect 7169 13417 7510 13445
rect 7169 13414 7181 13417
rect 7123 13408 7181 13414
rect 7504 13405 7510 13417
rect 7562 13405 7568 13457
rect 10096 13405 10102 13457
rect 10154 13405 10160 13457
rect 1152 13346 10560 13368
rect 1152 13294 4966 13346
rect 5018 13294 5030 13346
rect 5082 13294 5094 13346
rect 5146 13294 5158 13346
rect 5210 13294 5222 13346
rect 5274 13294 5286 13346
rect 5338 13294 10560 13346
rect 1152 13272 10560 13294
rect 2704 13109 2710 13161
rect 2762 13149 2768 13161
rect 4336 13149 4342 13161
rect 2762 13121 4342 13149
rect 2762 13109 2768 13121
rect 4336 13109 4342 13121
rect 4394 13149 4400 13161
rect 4394 13121 7838 13149
rect 4394 13109 4400 13121
rect 7810 13084 7838 13121
rect 7795 13078 7853 13084
rect 7795 13044 7807 13078
rect 7841 13044 7853 13078
rect 7795 13038 7853 13044
rect 1552 12961 1558 13013
rect 1610 12961 1616 13013
rect 1747 13004 1805 13010
rect 1747 12970 1759 13004
rect 1793 12970 1805 13004
rect 1747 12964 1805 12970
rect 1456 12887 1462 12939
rect 1514 12927 1520 12939
rect 1762 12927 1790 12964
rect 2896 12961 2902 13013
rect 2954 13001 2960 13013
rect 2995 13004 3053 13010
rect 2995 13001 3007 13004
rect 2954 12973 3007 13001
rect 2954 12961 2960 12973
rect 2995 12970 3007 12973
rect 3041 12970 3053 13004
rect 2995 12964 3053 12970
rect 3376 12961 3382 13013
rect 3434 12961 3440 13013
rect 5011 13004 5069 13010
rect 5011 12970 5023 13004
rect 5057 13001 5069 13004
rect 5488 13001 5494 13013
rect 5057 12973 5494 13001
rect 5057 12970 5069 12973
rect 5011 12964 5069 12970
rect 5488 12961 5494 12973
rect 5546 12961 5552 13013
rect 8179 13004 8237 13010
rect 8179 12970 8191 13004
rect 8225 13001 8237 13004
rect 8368 13001 8374 13013
rect 8225 12973 8374 13001
rect 8225 12970 8237 12973
rect 8179 12964 8237 12970
rect 8368 12961 8374 12973
rect 8426 12961 8432 13013
rect 8758 12939 8810 12945
rect 1514 12899 1790 12927
rect 1514 12887 1520 12899
rect 2800 12887 2806 12939
rect 2858 12927 2864 12939
rect 2858 12899 3216 12927
rect 2858 12887 2864 12899
rect 8758 12881 8810 12887
rect 9712 12739 9718 12791
rect 9770 12739 9776 12791
rect 1152 12680 10560 12702
rect 1152 12628 1966 12680
rect 2018 12628 2030 12680
rect 2082 12628 2094 12680
rect 2146 12628 2158 12680
rect 2210 12628 2222 12680
rect 2274 12628 2286 12680
rect 2338 12628 7966 12680
rect 8018 12628 8030 12680
rect 8082 12628 8094 12680
rect 8146 12628 8158 12680
rect 8210 12628 8222 12680
rect 8274 12628 8286 12680
rect 8338 12628 10560 12680
rect 1152 12606 10560 12628
rect 2800 12369 2806 12421
rect 2858 12369 2864 12421
rect 6160 12369 6166 12421
rect 6218 12369 6224 12421
rect 7216 12369 7222 12421
rect 7274 12369 7280 12421
rect 1840 12295 1846 12347
rect 1898 12335 1904 12347
rect 1939 12338 1997 12344
rect 1939 12335 1951 12338
rect 1898 12307 1951 12335
rect 1898 12295 1904 12307
rect 1939 12304 1951 12307
rect 1985 12335 1997 12338
rect 3280 12335 3286 12347
rect 1985 12307 3286 12335
rect 1985 12304 1997 12307
rect 1939 12298 1997 12304
rect 3280 12295 3286 12307
rect 3338 12295 3344 12347
rect 6544 12295 6550 12347
rect 6602 12295 6608 12347
rect 1456 12221 1462 12273
rect 1514 12261 1520 12273
rect 1555 12264 1613 12270
rect 1555 12261 1567 12264
rect 1514 12233 1567 12261
rect 1514 12221 1520 12233
rect 1555 12230 1567 12233
rect 1601 12230 1613 12264
rect 1555 12224 1613 12230
rect 3571 12116 3629 12122
rect 3571 12082 3583 12116
rect 3617 12113 3629 12116
rect 3664 12113 3670 12125
rect 3617 12085 3670 12113
rect 3617 12082 3629 12085
rect 3571 12076 3629 12082
rect 3664 12073 3670 12085
rect 3722 12113 3728 12125
rect 4240 12113 4246 12125
rect 3722 12085 4246 12113
rect 3722 12073 3728 12085
rect 4240 12073 4246 12085
rect 4298 12073 4304 12125
rect 8179 12116 8237 12122
rect 8179 12082 8191 12116
rect 8225 12113 8237 12116
rect 10192 12113 10198 12125
rect 8225 12085 10198 12113
rect 8225 12082 8237 12085
rect 8179 12076 8237 12082
rect 10192 12073 10198 12085
rect 10250 12073 10256 12125
rect 1152 12014 10560 12036
rect 1152 11962 4966 12014
rect 5018 11962 5030 12014
rect 5082 11962 5094 12014
rect 5146 11962 5158 12014
rect 5210 11962 5222 12014
rect 5274 11962 5286 12014
rect 5338 11962 10560 12014
rect 1152 11940 10560 11962
rect 3088 11851 3094 11903
rect 3146 11891 3152 11903
rect 4435 11894 4493 11900
rect 4435 11891 4447 11894
rect 3146 11863 4447 11891
rect 3146 11851 3152 11863
rect 4435 11860 4447 11863
rect 4481 11891 4493 11894
rect 7696 11891 7702 11903
rect 4481 11863 7702 11891
rect 4481 11860 4493 11863
rect 4435 11854 4493 11860
rect 7696 11851 7702 11863
rect 7754 11851 7760 11903
rect 1456 11703 1462 11755
rect 1514 11743 1520 11755
rect 1514 11715 2846 11743
rect 1514 11703 1520 11715
rect 1843 11672 1901 11678
rect 1843 11638 1855 11672
rect 1889 11669 1901 11672
rect 2704 11669 2710 11681
rect 1889 11641 2710 11669
rect 1889 11638 1901 11641
rect 1843 11632 1901 11638
rect 2704 11629 2710 11641
rect 2762 11629 2768 11681
rect 2818 11678 2846 11715
rect 2803 11672 2861 11678
rect 2803 11638 2815 11672
rect 2849 11638 2861 11672
rect 2803 11632 2861 11638
rect 5872 11629 5878 11681
rect 5930 11669 5936 11681
rect 6835 11672 6893 11678
rect 6835 11669 6847 11672
rect 5930 11641 6847 11669
rect 5930 11629 5936 11641
rect 6835 11638 6847 11641
rect 6881 11638 6893 11672
rect 6835 11632 6893 11638
rect 2419 11598 2477 11604
rect 2419 11564 2431 11598
rect 2465 11564 2477 11598
rect 2419 11558 2477 11564
rect 2434 11521 2462 11558
rect 2992 11521 2998 11533
rect 2434 11493 2998 11521
rect 2992 11481 2998 11493
rect 3050 11481 3056 11533
rect 1552 11407 1558 11459
rect 1610 11407 1616 11459
rect 2800 11407 2806 11459
rect 2858 11447 2864 11459
rect 3106 11447 3134 11581
rect 6160 11555 6166 11607
rect 6218 11595 6224 11607
rect 6451 11598 6509 11604
rect 6451 11595 6463 11598
rect 6218 11567 6463 11595
rect 6218 11555 6224 11567
rect 6451 11564 6463 11567
rect 6497 11564 6509 11598
rect 6451 11558 6509 11564
rect 7216 11555 7222 11607
rect 7274 11555 7280 11607
rect 8464 11555 8470 11607
rect 8522 11555 8528 11607
rect 2858 11419 3134 11447
rect 2858 11407 2864 11419
rect 1152 11348 10560 11370
rect 1152 11296 1966 11348
rect 2018 11296 2030 11348
rect 2082 11296 2094 11348
rect 2146 11296 2158 11348
rect 2210 11296 2222 11348
rect 2274 11296 2286 11348
rect 2338 11296 7966 11348
rect 8018 11296 8030 11348
rect 8082 11296 8094 11348
rect 8146 11296 8158 11348
rect 8210 11296 8222 11348
rect 8274 11296 8286 11348
rect 8338 11296 10560 11348
rect 1152 11274 10560 11296
rect 2512 11185 2518 11237
rect 2570 11225 2576 11237
rect 3475 11228 3533 11234
rect 3475 11225 3487 11228
rect 2570 11197 3487 11225
rect 2570 11185 2576 11197
rect 3475 11194 3487 11197
rect 3521 11225 3533 11228
rect 7792 11225 7798 11237
rect 3521 11197 7798 11225
rect 3521 11194 3533 11197
rect 3475 11188 3533 11194
rect 7792 11185 7798 11197
rect 7850 11185 7856 11237
rect 2992 11151 2998 11163
rect 1570 11123 2998 11151
rect 1570 11086 1598 11123
rect 2992 11111 2998 11123
rect 3050 11111 3056 11163
rect 7222 11089 7274 11095
rect 1555 11080 1613 11086
rect 1555 11046 1567 11080
rect 1601 11046 1613 11080
rect 1555 11040 1613 11046
rect 2800 11037 2806 11089
rect 2858 11037 2864 11089
rect 1936 10963 1942 11015
rect 1994 10963 2000 11015
rect 2818 11003 2846 11037
rect 4066 11003 4094 11063
rect 6160 11037 6166 11089
rect 6218 11077 6224 11089
rect 6259 11080 6317 11086
rect 6259 11077 6271 11080
rect 6218 11049 6271 11077
rect 6218 11037 6224 11049
rect 6259 11046 6271 11049
rect 6305 11046 6317 11080
rect 6259 11040 6317 11046
rect 7222 11031 7274 11037
rect 2818 10975 4094 11003
rect 4240 10963 4246 11015
rect 4298 10963 4304 11015
rect 6643 11006 6701 11012
rect 6643 10972 6655 11006
rect 6689 11003 6701 11006
rect 6736 11003 6742 11015
rect 6689 10975 6742 11003
rect 6689 10972 6701 10975
rect 6643 10966 6701 10972
rect 6736 10963 6742 10975
rect 6794 10963 6800 11015
rect 9808 10963 9814 11015
rect 9866 10963 9872 11015
rect 2896 10889 2902 10941
rect 2954 10929 2960 10941
rect 3859 10932 3917 10938
rect 3859 10929 3871 10932
rect 2954 10901 3871 10929
rect 2954 10889 2960 10901
rect 3859 10898 3871 10901
rect 3905 10898 3917 10932
rect 3859 10892 3917 10898
rect 4432 10741 4438 10793
rect 4490 10781 4496 10793
rect 5875 10784 5933 10790
rect 5875 10781 5887 10784
rect 4490 10753 5887 10781
rect 4490 10741 4496 10753
rect 5875 10750 5887 10753
rect 5921 10750 5933 10784
rect 5875 10744 5933 10750
rect 8275 10784 8333 10790
rect 8275 10750 8287 10784
rect 8321 10781 8333 10784
rect 9424 10781 9430 10793
rect 8321 10753 9430 10781
rect 8321 10750 8333 10753
rect 8275 10744 8333 10750
rect 9424 10741 9430 10753
rect 9482 10741 9488 10793
rect 10096 10741 10102 10793
rect 10154 10741 10160 10793
rect 1152 10682 10560 10704
rect 1152 10630 4966 10682
rect 5018 10630 5030 10682
rect 5082 10630 5094 10682
rect 5146 10630 5158 10682
rect 5210 10630 5222 10682
rect 5274 10630 5286 10682
rect 5338 10630 10560 10682
rect 1152 10608 10560 10630
rect 4336 10519 4342 10571
rect 4394 10519 4400 10571
rect 2323 10414 2381 10420
rect 2323 10380 2335 10414
rect 2369 10411 2381 10414
rect 2992 10411 2998 10423
rect 2369 10383 2998 10411
rect 2369 10380 2381 10383
rect 2323 10374 2381 10380
rect 2992 10371 2998 10383
rect 3050 10371 3056 10423
rect 7696 10371 7702 10423
rect 7754 10371 7760 10423
rect 1843 10340 1901 10346
rect 1843 10306 1855 10340
rect 1889 10337 1901 10340
rect 1936 10337 1942 10349
rect 1889 10309 1942 10337
rect 1889 10306 1901 10309
rect 1843 10300 1901 10306
rect 1936 10297 1942 10309
rect 1994 10297 2000 10349
rect 2704 10297 2710 10349
rect 2762 10337 2768 10349
rect 3664 10337 3670 10349
rect 2762 10309 3670 10337
rect 2762 10297 2768 10309
rect 3664 10297 3670 10309
rect 3722 10297 3728 10349
rect 8083 10340 8141 10346
rect 8083 10306 8095 10340
rect 8129 10337 8141 10340
rect 8368 10337 8374 10349
rect 8129 10309 8374 10337
rect 8129 10306 8141 10309
rect 8083 10300 8141 10306
rect 8368 10297 8374 10309
rect 8426 10297 8432 10349
rect 2722 10201 2750 10249
rect 8752 10223 8758 10275
rect 8810 10223 8816 10275
rect 2704 10149 2710 10201
rect 2762 10149 2768 10201
rect 1552 10075 1558 10127
rect 1610 10075 1616 10127
rect 9715 10118 9773 10124
rect 9715 10084 9727 10118
rect 9761 10115 9773 10118
rect 9808 10115 9814 10127
rect 9761 10087 9814 10115
rect 9761 10084 9773 10087
rect 9715 10078 9773 10084
rect 9808 10075 9814 10087
rect 9866 10075 9872 10127
rect 1152 10016 10560 10038
rect 1152 9964 1966 10016
rect 2018 9964 2030 10016
rect 2082 9964 2094 10016
rect 2146 9964 2158 10016
rect 2210 9964 2222 10016
rect 2274 9964 2286 10016
rect 2338 9964 7966 10016
rect 8018 9964 8030 10016
rect 8082 9964 8094 10016
rect 8146 9964 8158 10016
rect 8210 9964 8222 10016
rect 8274 9964 8286 10016
rect 8338 9964 10560 10016
rect 1152 9942 10560 9964
rect 1152 9350 10560 9372
rect 1152 9298 4966 9350
rect 5018 9298 5030 9350
rect 5082 9298 5094 9350
rect 5146 9298 5158 9350
rect 5210 9298 5222 9350
rect 5274 9298 5286 9350
rect 5338 9298 10560 9350
rect 1152 9276 10560 9298
rect 7792 9039 7798 9091
rect 7850 9039 7856 9091
rect 8179 9008 8237 9014
rect 8179 8974 8191 9008
rect 8225 9005 8237 9008
rect 8368 9005 8374 9017
rect 8225 8977 8374 9005
rect 8225 8974 8237 8977
rect 8179 8968 8237 8974
rect 8368 8965 8374 8977
rect 8426 8965 8432 9017
rect 8758 8943 8810 8949
rect 1648 8891 1654 8943
rect 1706 8891 1712 8943
rect 1747 8934 1805 8940
rect 1747 8900 1759 8934
rect 1793 8931 1805 8934
rect 2896 8931 2902 8943
rect 1793 8903 2902 8931
rect 1793 8900 1805 8903
rect 1747 8894 1805 8900
rect 2896 8891 2902 8903
rect 2954 8891 2960 8943
rect 8758 8885 8810 8891
rect 9811 8786 9869 8792
rect 9811 8752 9823 8786
rect 9857 8783 9869 8786
rect 10000 8783 10006 8795
rect 9857 8755 10006 8783
rect 9857 8752 9869 8755
rect 9811 8746 9869 8752
rect 10000 8743 10006 8755
rect 10058 8743 10064 8795
rect 1152 8684 10560 8706
rect 1152 8632 1966 8684
rect 2018 8632 2030 8684
rect 2082 8632 2094 8684
rect 2146 8632 2158 8684
rect 2210 8632 2222 8684
rect 2274 8632 2286 8684
rect 2338 8632 7966 8684
rect 8018 8632 8030 8684
rect 8082 8632 8094 8684
rect 8146 8632 8158 8684
rect 8210 8632 8222 8684
rect 8274 8632 8286 8684
rect 8338 8632 10560 8684
rect 1152 8610 10560 8632
rect 1744 8521 1750 8573
rect 1802 8521 1808 8573
rect 6256 8373 6262 8425
rect 6314 8373 6320 8425
rect 7696 8299 7702 8351
rect 7754 8299 7760 8351
rect 9520 8299 9526 8351
rect 9578 8339 9584 8351
rect 9811 8342 9869 8348
rect 9811 8339 9823 8342
rect 9578 8311 9823 8339
rect 9578 8299 9584 8311
rect 9811 8308 9823 8311
rect 9857 8308 9869 8342
rect 9811 8302 9869 8308
rect 10096 8299 10102 8351
rect 10154 8299 10160 8351
rect 1648 8225 1654 8277
rect 1706 8225 1712 8277
rect 1152 8018 10560 8040
rect 1152 7966 4966 8018
rect 5018 7966 5030 8018
rect 5082 7966 5094 8018
rect 5146 7966 5158 8018
rect 5210 7966 5222 8018
rect 5274 7966 5286 8018
rect 5338 7966 10560 8018
rect 1152 7944 10560 7966
rect 3664 7855 3670 7907
rect 3722 7855 3728 7907
rect 6352 7855 6358 7907
rect 6410 7895 6416 7907
rect 8179 7898 8237 7904
rect 8179 7895 8191 7898
rect 6410 7867 8191 7895
rect 6410 7855 6416 7867
rect 8179 7864 8191 7867
rect 8225 7864 8237 7898
rect 8179 7858 8237 7864
rect 1552 7707 1558 7759
rect 1610 7747 1616 7759
rect 1651 7750 1709 7756
rect 1651 7747 1663 7750
rect 1610 7719 1663 7747
rect 1610 7707 1616 7719
rect 1651 7716 1663 7719
rect 1697 7747 1709 7750
rect 1840 7747 1846 7759
rect 1697 7719 1846 7747
rect 1697 7716 1709 7719
rect 1651 7710 1709 7716
rect 1840 7707 1846 7719
rect 1898 7707 1904 7759
rect 8083 7750 8141 7756
rect 8083 7716 8095 7750
rect 8129 7747 8141 7750
rect 8368 7747 8374 7759
rect 8129 7719 8374 7747
rect 8129 7716 8141 7719
rect 8083 7710 8141 7716
rect 8368 7707 8374 7719
rect 8426 7707 8432 7759
rect 1744 7633 1750 7685
rect 1802 7673 1808 7685
rect 2035 7676 2093 7682
rect 2035 7673 2047 7676
rect 1802 7645 2047 7673
rect 1802 7633 1808 7645
rect 2035 7642 2047 7645
rect 2081 7673 2093 7676
rect 2800 7673 2806 7685
rect 2081 7645 2806 7673
rect 2081 7642 2093 7645
rect 2035 7636 2093 7642
rect 2800 7633 2806 7645
rect 2858 7633 2864 7685
rect 7123 7676 7181 7682
rect 7123 7642 7135 7676
rect 7169 7642 7181 7676
rect 7123 7636 7181 7642
rect 2704 7559 2710 7611
rect 2762 7559 2768 7611
rect 7138 7599 7166 7636
rect 7891 7602 7949 7608
rect 7891 7599 7903 7602
rect 7138 7571 7903 7599
rect 7891 7568 7903 7571
rect 7937 7568 7949 7602
rect 7891 7562 7949 7568
rect 1456 7485 1462 7537
rect 1514 7525 1520 7537
rect 1744 7525 1750 7537
rect 1514 7497 1750 7525
rect 1514 7485 1520 7497
rect 1744 7485 1750 7497
rect 1802 7485 1808 7537
rect 6832 7411 6838 7463
rect 6890 7411 6896 7463
rect 1152 7352 10560 7374
rect 1152 7300 1966 7352
rect 2018 7300 2030 7352
rect 2082 7300 2094 7352
rect 2146 7300 2158 7352
rect 2210 7300 2222 7352
rect 2274 7300 2286 7352
rect 2338 7300 7966 7352
rect 8018 7300 8030 7352
rect 8082 7300 8094 7352
rect 8146 7300 8158 7352
rect 8210 7300 8222 7352
rect 8274 7300 8286 7352
rect 8338 7300 10560 7352
rect 1152 7278 10560 7300
rect 1552 7189 1558 7241
rect 1610 7229 1616 7241
rect 1651 7232 1709 7238
rect 1651 7229 1663 7232
rect 1610 7201 1663 7229
rect 1610 7189 1616 7201
rect 1651 7198 1663 7201
rect 1697 7198 1709 7232
rect 1651 7192 1709 7198
rect 8179 7232 8237 7238
rect 8179 7198 8191 7232
rect 8225 7229 8237 7232
rect 8368 7229 8374 7241
rect 8225 7201 8374 7229
rect 8225 7198 8237 7201
rect 8179 7192 8237 7198
rect 8368 7189 8374 7201
rect 8426 7189 8432 7241
rect 6643 7084 6701 7090
rect 2800 6967 2806 7019
rect 2858 7007 2864 7019
rect 3283 7010 3341 7016
rect 3283 7007 3295 7010
rect 2858 6979 3295 7007
rect 2858 6967 2864 6979
rect 3283 6976 3295 6979
rect 3329 6976 3341 7010
rect 3283 6970 3341 6976
rect 2704 6893 2710 6945
rect 2762 6933 2768 6945
rect 3490 6933 3518 7067
rect 6643 7050 6655 7084
rect 6689 7081 6701 7084
rect 6832 7081 6838 7093
rect 6689 7053 6838 7081
rect 6689 7050 6701 7053
rect 6643 7044 6701 7050
rect 6832 7041 6838 7053
rect 6890 7041 6896 7093
rect 6256 6967 6262 7019
rect 6314 7007 6320 7019
rect 6448 7007 6454 7019
rect 6314 6979 6454 7007
rect 6314 6967 6320 6979
rect 6448 6967 6454 6979
rect 6506 6967 6512 7019
rect 8563 7010 8621 7016
rect 8563 6976 8575 7010
rect 8609 7007 8621 7010
rect 9520 7007 9526 7019
rect 8609 6979 9526 7007
rect 8609 6976 8621 6979
rect 8563 6970 8621 6976
rect 9520 6967 9526 6979
rect 9578 6967 9584 7019
rect 3667 6936 3725 6942
rect 3667 6933 3679 6936
rect 2762 6905 3679 6933
rect 2762 6893 2768 6905
rect 3667 6902 3679 6905
rect 3713 6902 3725 6936
rect 8761 6936 8819 6942
rect 8761 6933 8773 6936
rect 3667 6896 3725 6902
rect 7810 6905 8773 6933
rect 7810 6868 7838 6905
rect 8761 6902 8773 6905
rect 8807 6933 8819 6936
rect 8848 6933 8854 6945
rect 8807 6905 8854 6933
rect 8807 6902 8819 6905
rect 8761 6896 8819 6902
rect 8848 6893 8854 6905
rect 8906 6893 8912 6945
rect 7795 6862 7853 6868
rect 7795 6828 7807 6862
rect 7841 6828 7853 6862
rect 7795 6822 7853 6828
rect 1152 6686 10560 6708
rect 1152 6634 4966 6686
rect 5018 6634 5030 6686
rect 5082 6634 5094 6686
rect 5146 6634 5158 6686
rect 5210 6634 5222 6686
rect 5274 6634 5286 6686
rect 5338 6634 10560 6686
rect 1152 6612 10560 6634
rect 1744 6523 1750 6575
rect 1802 6523 1808 6575
rect 5872 6523 5878 6575
rect 5930 6563 5936 6575
rect 6259 6566 6317 6572
rect 6259 6563 6271 6566
rect 5930 6535 6271 6563
rect 5930 6523 5936 6535
rect 6259 6532 6271 6535
rect 6305 6563 6317 6566
rect 6352 6563 6358 6575
rect 6305 6535 6358 6563
rect 6305 6532 6317 6535
rect 6259 6526 6317 6532
rect 6352 6523 6358 6535
rect 6410 6523 6416 6575
rect 6064 6449 6070 6501
rect 6122 6489 6128 6501
rect 8179 6492 8237 6498
rect 8179 6489 8191 6492
rect 6122 6461 8191 6489
rect 6122 6449 6128 6461
rect 8179 6458 8191 6461
rect 8225 6458 8237 6492
rect 8179 6452 8237 6458
rect 2800 6375 2806 6427
rect 2858 6415 2864 6427
rect 5779 6418 5837 6424
rect 2858 6387 3422 6415
rect 2858 6375 2864 6387
rect 3394 6350 3422 6387
rect 5779 6384 5791 6418
rect 5825 6415 5837 6418
rect 5968 6415 5974 6427
rect 5825 6387 5974 6415
rect 5825 6384 5837 6387
rect 5779 6378 5837 6384
rect 5968 6375 5974 6387
rect 6026 6375 6032 6427
rect 8848 6375 8854 6427
rect 8906 6375 8912 6427
rect 3379 6344 3437 6350
rect 3379 6310 3391 6344
rect 3425 6310 3437 6344
rect 3379 6304 3437 6310
rect 5299 6344 5357 6350
rect 5299 6310 5311 6344
rect 5345 6310 5357 6344
rect 5299 6304 5357 6310
rect 2704 6153 2710 6205
rect 2762 6193 2768 6205
rect 3586 6193 3614 6253
rect 3760 6227 3766 6279
rect 3818 6227 3824 6279
rect 5314 6267 5342 6304
rect 5680 6301 5686 6353
rect 5738 6341 5744 6353
rect 6067 6344 6125 6350
rect 6067 6341 6079 6344
rect 5738 6313 6079 6341
rect 5738 6301 5744 6313
rect 6067 6310 6079 6313
rect 6113 6310 6125 6344
rect 6067 6304 6125 6310
rect 6448 6301 6454 6353
rect 6506 6341 6512 6353
rect 6547 6344 6605 6350
rect 6547 6341 6559 6344
rect 6506 6313 6559 6341
rect 6506 6301 6512 6313
rect 6547 6310 6559 6313
rect 6593 6310 6605 6344
rect 6547 6304 6605 6310
rect 7792 6301 7798 6353
rect 7850 6341 7856 6353
rect 8272 6341 8278 6353
rect 7850 6313 8278 6341
rect 7850 6301 7856 6313
rect 8272 6301 8278 6313
rect 8330 6301 8336 6353
rect 8371 6344 8429 6350
rect 8371 6310 8383 6344
rect 8417 6341 8429 6344
rect 8464 6341 8470 6353
rect 8417 6313 8470 6341
rect 8417 6310 8429 6313
rect 8371 6304 8429 6310
rect 8464 6301 8470 6313
rect 8522 6301 8528 6353
rect 9040 6341 9046 6353
rect 8962 6313 9046 6341
rect 5587 6270 5645 6276
rect 5587 6267 5599 6270
rect 5314 6239 5599 6267
rect 5587 6236 5599 6239
rect 5633 6236 5645 6270
rect 5587 6230 5645 6236
rect 6931 6270 6989 6276
rect 6931 6236 6943 6270
rect 6977 6267 6989 6270
rect 8962 6267 8990 6313
rect 9040 6301 9046 6313
rect 9098 6301 9104 6353
rect 9328 6301 9334 6353
rect 9386 6301 9392 6353
rect 9808 6301 9814 6353
rect 9866 6301 9872 6353
rect 6977 6239 7214 6267
rect 6977 6236 6989 6239
rect 6931 6230 6989 6236
rect 5680 6193 5686 6205
rect 2762 6165 5686 6193
rect 2762 6153 2768 6165
rect 5680 6153 5686 6165
rect 5738 6153 5744 6205
rect 5491 6122 5549 6128
rect 5491 6088 5503 6122
rect 5537 6119 5549 6122
rect 6832 6119 6838 6131
rect 5537 6091 6838 6119
rect 5537 6088 5549 6091
rect 5491 6082 5549 6088
rect 6832 6079 6838 6091
rect 6890 6079 6896 6131
rect 7186 6119 7214 6239
rect 8098 6239 8990 6267
rect 8098 6202 8126 6239
rect 8083 6196 8141 6202
rect 8083 6162 8095 6196
rect 8129 6162 8141 6196
rect 8083 6156 8141 6162
rect 8272 6153 8278 6205
rect 8330 6193 8336 6205
rect 8467 6196 8525 6202
rect 8467 6193 8479 6196
rect 8330 6165 8479 6193
rect 8330 6153 8336 6165
rect 8467 6162 8479 6165
rect 8513 6162 8525 6196
rect 8467 6156 8525 6162
rect 8368 6119 8374 6131
rect 7186 6091 8374 6119
rect 8368 6079 8374 6091
rect 8426 6079 8432 6131
rect 8560 6079 8566 6131
rect 8618 6119 8624 6131
rect 9139 6122 9197 6128
rect 9139 6119 9151 6122
rect 8618 6091 9151 6119
rect 8618 6079 8624 6091
rect 9139 6088 9151 6091
rect 9185 6088 9197 6122
rect 9139 6082 9197 6088
rect 10096 6079 10102 6131
rect 10154 6079 10160 6131
rect 1152 6020 10560 6042
rect 1152 5968 1966 6020
rect 2018 5968 2030 6020
rect 2082 5968 2094 6020
rect 2146 5968 2158 6020
rect 2210 5968 2222 6020
rect 2274 5968 2286 6020
rect 2338 5968 7966 6020
rect 8018 5968 8030 6020
rect 8082 5968 8094 6020
rect 8146 5968 8158 6020
rect 8210 5968 8222 6020
rect 8274 5968 8286 6020
rect 8338 5968 10560 6020
rect 1152 5946 10560 5968
rect 9619 5826 9677 5832
rect 9619 5823 9631 5826
rect 9442 5795 9631 5823
rect 1552 5709 1558 5761
rect 1610 5709 1616 5761
rect 2704 5709 2710 5761
rect 2762 5709 2768 5761
rect 7696 5709 7702 5761
rect 7754 5709 7760 5761
rect 8368 5709 8374 5761
rect 8426 5749 8432 5761
rect 9442 5749 9470 5795
rect 9619 5792 9631 5795
rect 9665 5792 9677 5826
rect 9619 5786 9677 5792
rect 8426 5721 9470 5749
rect 8426 5709 8432 5721
rect 9520 5709 9526 5761
rect 9578 5749 9584 5761
rect 9578 5721 9758 5749
rect 9578 5709 9584 5721
rect 1570 5675 1598 5709
rect 1939 5678 1997 5684
rect 1939 5675 1951 5678
rect 1570 5647 1951 5675
rect 1939 5644 1951 5647
rect 1985 5644 1997 5678
rect 5587 5678 5645 5684
rect 5587 5675 5599 5678
rect 1939 5638 1997 5644
rect 5026 5647 5599 5675
rect 1555 5604 1613 5610
rect 1555 5570 1567 5604
rect 1601 5601 1613 5604
rect 1648 5601 1654 5613
rect 1601 5573 1654 5601
rect 1601 5570 1613 5573
rect 1555 5564 1613 5570
rect 1648 5561 1654 5573
rect 1706 5601 1712 5613
rect 2896 5601 2902 5613
rect 1706 5573 2902 5601
rect 1706 5561 1712 5573
rect 2896 5561 2902 5573
rect 2954 5561 2960 5613
rect 4816 5561 4822 5613
rect 4874 5561 4880 5613
rect 5026 5610 5054 5647
rect 5587 5644 5599 5647
rect 5633 5675 5645 5678
rect 6064 5675 6070 5687
rect 5633 5647 6070 5675
rect 5633 5644 5645 5647
rect 5587 5638 5645 5644
rect 6064 5635 6070 5647
rect 6122 5635 6128 5687
rect 6352 5635 6358 5687
rect 6410 5635 6416 5687
rect 6658 5647 8606 5675
rect 5011 5604 5069 5610
rect 5011 5570 5023 5604
rect 5057 5570 5069 5604
rect 5011 5564 5069 5570
rect 5104 5561 5110 5613
rect 5162 5561 5168 5613
rect 5491 5604 5549 5610
rect 5491 5570 5503 5604
rect 5537 5601 5549 5604
rect 5680 5601 5686 5613
rect 5537 5573 5686 5601
rect 5537 5570 5549 5573
rect 5491 5564 5549 5570
rect 5680 5561 5686 5573
rect 5738 5561 5744 5613
rect 4915 5530 4973 5536
rect 4915 5496 4927 5530
rect 4961 5527 4973 5530
rect 6064 5527 6070 5539
rect 4961 5499 6070 5527
rect 4961 5496 4973 5499
rect 4915 5490 4973 5496
rect 6064 5487 6070 5499
rect 6122 5527 6128 5539
rect 6658 5527 6686 5647
rect 6122 5499 6686 5527
rect 8578 5527 8606 5647
rect 9040 5635 9046 5687
rect 9098 5675 9104 5687
rect 9331 5678 9389 5684
rect 9331 5675 9343 5678
rect 9098 5647 9343 5675
rect 9098 5635 9104 5647
rect 9331 5644 9343 5647
rect 9377 5644 9389 5678
rect 9331 5638 9389 5644
rect 9616 5635 9622 5687
rect 9674 5635 9680 5687
rect 9730 5684 9758 5721
rect 9715 5678 9773 5684
rect 9715 5644 9727 5678
rect 9761 5644 9773 5678
rect 9715 5638 9773 5644
rect 9136 5561 9142 5613
rect 9194 5601 9200 5613
rect 9235 5604 9293 5610
rect 9235 5601 9247 5604
rect 9194 5573 9247 5601
rect 9194 5561 9200 5573
rect 9235 5570 9247 5573
rect 9281 5570 9293 5604
rect 9235 5564 9293 5570
rect 9907 5604 9965 5610
rect 9907 5570 9919 5604
rect 9953 5570 9965 5604
rect 9907 5564 9965 5570
rect 9922 5527 9950 5564
rect 8578 5499 9950 5527
rect 6122 5487 6128 5499
rect 2896 5413 2902 5465
rect 2954 5453 2960 5465
rect 3571 5456 3629 5462
rect 3571 5453 3583 5456
rect 2954 5425 3583 5453
rect 2954 5413 2960 5425
rect 3571 5422 3583 5425
rect 3617 5422 3629 5456
rect 3571 5416 3629 5422
rect 5779 5456 5837 5462
rect 5779 5422 5791 5456
rect 5825 5453 5837 5456
rect 5968 5453 5974 5465
rect 5825 5425 5974 5453
rect 5825 5422 5837 5425
rect 5779 5416 5837 5422
rect 5968 5413 5974 5425
rect 6026 5413 6032 5465
rect 8368 5413 8374 5465
rect 8426 5453 8432 5465
rect 9139 5456 9197 5462
rect 9139 5453 9151 5456
rect 8426 5425 9151 5453
rect 8426 5413 8432 5425
rect 9139 5422 9151 5425
rect 9185 5422 9197 5456
rect 9139 5416 9197 5422
rect 1152 5354 10560 5376
rect 1152 5302 4966 5354
rect 5018 5302 5030 5354
rect 5082 5302 5094 5354
rect 5146 5302 5158 5354
rect 5210 5302 5222 5354
rect 5274 5302 5286 5354
rect 5338 5302 10560 5354
rect 1152 5280 10560 5302
rect 5680 5191 5686 5243
rect 5738 5231 5744 5243
rect 7987 5234 8045 5240
rect 7987 5231 7999 5234
rect 5738 5203 7999 5231
rect 5738 5191 5744 5203
rect 7987 5200 7999 5203
rect 8033 5200 8045 5234
rect 7987 5194 8045 5200
rect 9040 5191 9046 5243
rect 9098 5191 9104 5243
rect 9331 5234 9389 5240
rect 9331 5200 9343 5234
rect 9377 5231 9389 5234
rect 9616 5231 9622 5243
rect 9377 5203 9622 5231
rect 9377 5200 9389 5203
rect 9331 5194 9389 5200
rect 9616 5191 9622 5203
rect 9674 5191 9680 5243
rect 9058 5157 9086 5191
rect 9058 5129 9470 5157
rect 1648 5043 1654 5095
rect 1706 5043 1712 5095
rect 1840 5043 1846 5095
rect 1898 5043 1904 5095
rect 6832 5043 6838 5095
rect 6890 5043 6896 5095
rect 8368 5043 8374 5095
rect 8426 5083 8432 5095
rect 9043 5086 9101 5092
rect 9043 5083 9055 5086
rect 8426 5055 9055 5083
rect 8426 5043 8432 5055
rect 9043 5052 9055 5055
rect 9089 5052 9101 5086
rect 9043 5046 9101 5052
rect 1858 5009 1886 5043
rect 2035 5012 2093 5018
rect 2035 5009 2047 5012
rect 1858 4981 2047 5009
rect 2035 4978 2047 4981
rect 2081 4978 2093 5012
rect 2035 4972 2093 4978
rect 6163 5012 6221 5018
rect 6163 4978 6175 5012
rect 6209 4978 6221 5012
rect 6163 4972 6221 4978
rect 2704 4895 2710 4947
rect 2762 4895 2768 4947
rect 5776 4895 5782 4947
rect 5834 4895 5840 4947
rect 6178 4935 6206 4972
rect 6448 4969 6454 5021
rect 6506 4969 6512 5021
rect 7792 4969 7798 5021
rect 7850 5009 7856 5021
rect 8563 5012 8621 5018
rect 8563 5009 8575 5012
rect 7850 4981 8575 5009
rect 7850 4969 7856 4981
rect 8563 4978 8575 4981
rect 8609 4978 8621 5012
rect 9058 5009 9086 5046
rect 9136 5043 9142 5095
rect 9194 5083 9200 5095
rect 9442 5092 9470 5129
rect 9427 5086 9485 5092
rect 9194 5055 9374 5083
rect 9194 5043 9200 5055
rect 9235 5012 9293 5018
rect 9235 5009 9247 5012
rect 9058 4981 9247 5009
rect 8563 4972 8621 4978
rect 9235 4978 9247 4981
rect 9281 4978 9293 5012
rect 9235 4972 9293 4978
rect 6544 4935 6550 4947
rect 6178 4907 6550 4935
rect 6544 4895 6550 4907
rect 6602 4895 6608 4947
rect 8578 4935 8606 4972
rect 9346 4935 9374 5055
rect 9427 5052 9439 5086
rect 9473 5052 9485 5086
rect 9427 5046 9485 5052
rect 8578 4907 9374 4935
rect 3280 4747 3286 4799
rect 3338 4787 3344 4799
rect 3571 4790 3629 4796
rect 3571 4787 3583 4790
rect 3338 4759 3583 4787
rect 3338 4747 3344 4759
rect 3571 4756 3583 4759
rect 3617 4756 3629 4790
rect 3571 4750 3629 4756
rect 4624 4747 4630 4799
rect 4682 4747 4688 4799
rect 8371 4790 8429 4796
rect 8371 4756 8383 4790
rect 8417 4787 8429 4790
rect 8464 4787 8470 4799
rect 8417 4759 8470 4787
rect 8417 4756 8429 4759
rect 8371 4750 8429 4756
rect 8464 4747 8470 4759
rect 8522 4747 8528 4799
rect 1152 4688 10560 4710
rect 1152 4636 1966 4688
rect 2018 4636 2030 4688
rect 2082 4636 2094 4688
rect 2146 4636 2158 4688
rect 2210 4636 2222 4688
rect 2274 4636 2286 4688
rect 2338 4636 7966 4688
rect 8018 4636 8030 4688
rect 8082 4636 8094 4688
rect 8146 4636 8158 4688
rect 8210 4636 8222 4688
rect 8274 4636 8286 4688
rect 8338 4636 10560 4688
rect 1152 4614 10560 4636
rect 5776 4525 5782 4577
rect 5834 4565 5840 4577
rect 6163 4568 6221 4574
rect 6163 4565 6175 4568
rect 5834 4537 6175 4565
rect 5834 4525 5840 4537
rect 6163 4534 6175 4537
rect 6209 4534 6221 4568
rect 6163 4528 6221 4534
rect 8179 4568 8237 4574
rect 8179 4534 8191 4568
rect 8225 4565 8237 4568
rect 8368 4565 8374 4577
rect 8225 4537 8374 4565
rect 8225 4534 8237 4537
rect 8179 4528 8237 4534
rect 8368 4525 8374 4537
rect 8426 4525 8432 4577
rect 2710 4429 2762 4435
rect 6064 4417 6070 4429
rect 2710 4371 2762 4377
rect 5794 4389 6070 4417
rect 3283 4346 3341 4352
rect 3283 4312 3295 4346
rect 3329 4343 3341 4346
rect 3760 4343 3766 4355
rect 3329 4315 3766 4343
rect 3329 4312 3341 4315
rect 3283 4306 3341 4312
rect 3760 4303 3766 4315
rect 3818 4303 3824 4355
rect 4624 4303 4630 4355
rect 4682 4343 4688 4355
rect 5794 4352 5822 4389
rect 6064 4377 6070 4389
rect 6122 4417 6128 4429
rect 7027 4420 7085 4426
rect 6122 4389 6302 4417
rect 6122 4377 6128 4389
rect 5683 4346 5741 4352
rect 5683 4343 5695 4346
rect 4682 4315 5695 4343
rect 4682 4303 4688 4315
rect 5683 4312 5695 4315
rect 5729 4312 5741 4346
rect 5683 4306 5741 4312
rect 5779 4346 5837 4352
rect 5779 4312 5791 4346
rect 5825 4312 5837 4346
rect 5779 4306 5837 4312
rect 5968 4303 5974 4355
rect 6026 4303 6032 4355
rect 6274 4352 6302 4389
rect 7027 4386 7039 4420
rect 7073 4417 7085 4420
rect 8560 4417 8566 4429
rect 7073 4389 8566 4417
rect 7073 4386 7085 4389
rect 7027 4380 7085 4386
rect 8560 4377 8566 4389
rect 8618 4377 8624 4429
rect 6259 4346 6317 4352
rect 6259 4312 6271 4346
rect 6305 4312 6317 4346
rect 6259 4306 6317 4312
rect 6451 4346 6509 4352
rect 6451 4312 6463 4346
rect 6497 4312 6509 4346
rect 6451 4306 6509 4312
rect 2992 4229 2998 4281
rect 3050 4269 3056 4281
rect 3667 4272 3725 4278
rect 3667 4269 3679 4272
rect 3050 4241 3679 4269
rect 3050 4229 3056 4241
rect 3667 4238 3679 4241
rect 3713 4238 3725 4272
rect 3667 4232 3725 4238
rect 6466 4195 6494 4306
rect 6544 4303 6550 4355
rect 6602 4343 6608 4355
rect 6643 4346 6701 4352
rect 6643 4343 6655 4346
rect 6602 4315 6655 4343
rect 6602 4303 6608 4315
rect 6643 4312 6655 4315
rect 6689 4312 6701 4346
rect 6643 4306 6701 4312
rect 7120 4303 7126 4355
rect 7178 4343 7184 4355
rect 7696 4343 7702 4355
rect 7178 4315 7702 4343
rect 7178 4303 7184 4315
rect 7696 4303 7702 4315
rect 7754 4303 7760 4355
rect 8464 4229 8470 4281
rect 8522 4229 8528 4281
rect 7792 4195 7798 4207
rect 6466 4167 7798 4195
rect 7792 4155 7798 4167
rect 7850 4195 7856 4207
rect 8080 4195 8086 4207
rect 7850 4167 8086 4195
rect 7850 4155 7856 4167
rect 8080 4155 8086 4167
rect 8138 4155 8144 4207
rect 8659 4198 8717 4204
rect 8659 4164 8671 4198
rect 8705 4195 8717 4198
rect 9328 4195 9334 4207
rect 8705 4167 9334 4195
rect 8705 4164 8717 4167
rect 8659 4158 8717 4164
rect 9328 4155 9334 4167
rect 9386 4155 9392 4207
rect 1648 4081 1654 4133
rect 1706 4081 1712 4133
rect 6352 4081 6358 4133
rect 6410 4081 6416 4133
rect 8371 4124 8429 4130
rect 8371 4090 8383 4124
rect 8417 4121 8429 4124
rect 8752 4121 8758 4133
rect 8417 4093 8758 4121
rect 8417 4090 8429 4093
rect 8371 4084 8429 4090
rect 8752 4081 8758 4093
rect 8810 4081 8816 4133
rect 1152 4022 10560 4044
rect 1152 3970 4966 4022
rect 5018 3970 5030 4022
rect 5082 3970 5094 4022
rect 5146 3970 5158 4022
rect 5210 3970 5222 4022
rect 5274 3970 5286 4022
rect 5338 3970 10560 4022
rect 1152 3948 10560 3970
rect 5872 3859 5878 3911
rect 5930 3859 5936 3911
rect 6163 3902 6221 3908
rect 6163 3868 6175 3902
rect 6209 3868 6221 3902
rect 6163 3862 6221 3868
rect 2515 3828 2573 3834
rect 2515 3794 2527 3828
rect 2561 3825 2573 3828
rect 4816 3825 4822 3837
rect 2561 3797 4822 3825
rect 2561 3794 2573 3797
rect 2515 3788 2573 3794
rect 4816 3785 4822 3797
rect 4874 3825 4880 3837
rect 6178 3825 6206 3862
rect 8080 3859 8086 3911
rect 8138 3859 8144 3911
rect 8752 3825 8758 3837
rect 4874 3797 8758 3825
rect 4874 3785 4880 3797
rect 8752 3785 8758 3797
rect 8810 3785 8816 3837
rect 6067 3754 6125 3760
rect 6067 3720 6079 3754
rect 6113 3751 6125 3754
rect 6160 3751 6166 3763
rect 6113 3723 6166 3751
rect 6113 3720 6125 3723
rect 6067 3714 6125 3720
rect 6160 3711 6166 3723
rect 6218 3711 6224 3763
rect 6352 3711 6358 3763
rect 6410 3751 6416 3763
rect 6931 3754 6989 3760
rect 6931 3751 6943 3754
rect 6410 3723 6943 3751
rect 6410 3711 6416 3723
rect 6931 3720 6943 3723
rect 6977 3720 6989 3754
rect 6931 3714 6989 3720
rect 880 3637 886 3689
rect 938 3677 944 3689
rect 1555 3680 1613 3686
rect 1555 3677 1567 3680
rect 938 3649 1567 3677
rect 938 3637 944 3649
rect 1555 3646 1567 3649
rect 1601 3646 1613 3680
rect 1555 3640 1613 3646
rect 6544 3637 6550 3689
rect 6602 3637 6608 3689
rect 7504 3637 7510 3689
rect 7562 3677 7568 3689
rect 8371 3680 8429 3686
rect 8371 3677 8383 3680
rect 7562 3649 8383 3677
rect 7562 3637 7568 3649
rect 8371 3646 8383 3649
rect 8417 3646 8429 3680
rect 8371 3640 8429 3646
rect 9424 3637 9430 3689
rect 9482 3637 9488 3689
rect 9712 3637 9718 3689
rect 9770 3677 9776 3689
rect 9811 3680 9869 3686
rect 9811 3677 9823 3680
rect 9770 3649 9823 3677
rect 9770 3637 9776 3649
rect 9811 3646 9823 3649
rect 9857 3646 9869 3680
rect 9811 3640 9869 3646
rect 10096 3563 10102 3615
rect 10154 3563 10160 3615
rect 7504 3489 7510 3541
rect 7562 3529 7568 3541
rect 8179 3532 8237 3538
rect 8179 3529 8191 3532
rect 7562 3501 8191 3529
rect 7562 3489 7568 3501
rect 8179 3498 8191 3501
rect 8225 3498 8237 3532
rect 8179 3492 8237 3498
rect 9715 3458 9773 3464
rect 9715 3424 9727 3458
rect 9761 3455 9773 3458
rect 10960 3455 10966 3467
rect 9761 3427 10966 3455
rect 9761 3424 9773 3427
rect 9715 3418 9773 3424
rect 10960 3415 10966 3427
rect 11018 3415 11024 3467
rect 1152 3356 10560 3378
rect 1152 3304 1966 3356
rect 2018 3304 2030 3356
rect 2082 3304 2094 3356
rect 2146 3304 2158 3356
rect 2210 3304 2222 3356
rect 2274 3304 2286 3356
rect 2338 3304 7966 3356
rect 8018 3304 8030 3356
rect 8082 3304 8094 3356
rect 8146 3304 8158 3356
rect 8210 3304 8222 3356
rect 8274 3304 8286 3356
rect 8338 3304 10560 3356
rect 1152 3282 10560 3304
rect 7888 3193 7894 3245
rect 7946 3233 7952 3245
rect 7946 3205 9278 3233
rect 7946 3193 7952 3205
rect 592 3045 598 3097
rect 650 3085 656 3097
rect 2611 3088 2669 3094
rect 2611 3085 2623 3088
rect 650 3057 2623 3085
rect 650 3045 656 3057
rect 2611 3054 2623 3057
rect 2657 3054 2669 3088
rect 4624 3085 4630 3097
rect 2611 3048 2669 3054
rect 2818 3057 4630 3085
rect 1648 2971 1654 3023
rect 1706 3011 1712 3023
rect 2035 3014 2093 3020
rect 2035 3011 2047 3014
rect 1706 2983 2047 3011
rect 1706 2971 1712 2983
rect 2035 2980 2047 2983
rect 2081 2980 2093 3014
rect 2035 2974 2093 2980
rect 2515 3014 2573 3020
rect 2515 2980 2527 3014
rect 2561 3011 2573 3014
rect 2818 3011 2846 3057
rect 4624 3045 4630 3057
rect 4682 3045 4688 3097
rect 6544 3045 6550 3097
rect 6602 3085 6608 3097
rect 6602 3057 7440 3085
rect 6602 3045 6608 3057
rect 2561 2983 2846 3011
rect 2561 2980 2573 2983
rect 2515 2974 2573 2980
rect 2896 2971 2902 3023
rect 2954 2971 2960 3023
rect 3280 2971 3286 3023
rect 3338 2971 3344 3023
rect 4432 2971 4438 3023
rect 4490 2971 4496 3023
rect 5488 2971 5494 3023
rect 5546 2971 5552 3023
rect 6739 3014 6797 3020
rect 6739 2980 6751 3014
rect 6785 3011 6797 3014
rect 7024 3011 7030 3023
rect 6785 2983 7030 3011
rect 6785 2980 6797 2983
rect 6739 2974 6797 2980
rect 7024 2971 7030 2983
rect 7082 2971 7088 3023
rect 7120 2971 7126 3023
rect 7178 2971 7184 3023
rect 9250 3020 9278 3205
rect 9235 3014 9293 3020
rect 9235 2980 9247 3014
rect 9281 2980 9293 3014
rect 9235 2974 9293 2980
rect 9523 3014 9581 3020
rect 9523 2980 9535 3014
rect 9569 3011 9581 3014
rect 10000 3011 10006 3023
rect 9569 2983 10006 3011
rect 9569 2980 9581 2983
rect 9523 2974 9581 2980
rect 10000 2971 10006 2983
rect 10058 2971 10064 3023
rect 10099 3014 10157 3020
rect 10099 2980 10111 3014
rect 10145 3011 10157 3014
rect 10192 3011 10198 3023
rect 10145 2983 10198 3011
rect 10145 2980 10157 2983
rect 10099 2974 10157 2980
rect 10192 2971 10198 2983
rect 10250 2971 10256 3023
rect 1840 2897 1846 2949
rect 1898 2897 1904 2949
rect 2992 2897 2998 2949
rect 3050 2897 3056 2949
rect 4144 2897 4150 2949
rect 4202 2897 4208 2949
rect 5299 2940 5357 2946
rect 5299 2906 5311 2940
rect 5345 2937 5357 2940
rect 5392 2937 5398 2949
rect 5345 2909 5398 2937
rect 5345 2906 5357 2909
rect 5299 2900 5357 2906
rect 5392 2897 5398 2909
rect 5450 2897 5456 2949
rect 6448 2897 6454 2949
rect 6506 2897 6512 2949
rect 8848 2897 8854 2949
rect 8906 2937 8912 2949
rect 9043 2940 9101 2946
rect 9043 2937 9055 2940
rect 8906 2909 9055 2937
rect 8906 2897 8912 2909
rect 9043 2906 9055 2909
rect 9089 2906 9101 2940
rect 9043 2900 9101 2906
rect 9712 2897 9718 2949
rect 9770 2897 9776 2949
rect 9808 2897 9814 2949
rect 9866 2897 9872 2949
rect 2224 2749 2230 2801
rect 2282 2749 2288 2801
rect 1152 2690 10560 2712
rect 1152 2638 4966 2690
rect 5018 2638 5030 2690
rect 5082 2638 5094 2690
rect 5146 2638 5158 2690
rect 5210 2638 5222 2690
rect 5274 2638 5286 2690
rect 5338 2638 10560 2690
rect 1152 2616 10560 2638
<< via1 >>
rect 1966 25948 2018 26000
rect 2030 25948 2082 26000
rect 2094 25948 2146 26000
rect 2158 25948 2210 26000
rect 2222 25948 2274 26000
rect 2286 25948 2338 26000
rect 7966 25948 8018 26000
rect 8030 25948 8082 26000
rect 8094 25948 8146 26000
rect 8158 25948 8210 26000
rect 8222 25948 8274 26000
rect 8286 25948 8338 26000
rect 1750 25837 1802 25889
rect 2998 25880 3050 25889
rect 2998 25846 3007 25880
rect 3007 25846 3041 25880
rect 3041 25846 3050 25880
rect 2998 25837 3050 25846
rect 4150 25880 4202 25889
rect 4150 25846 4159 25880
rect 4159 25846 4193 25880
rect 4193 25846 4202 25880
rect 4150 25837 4202 25846
rect 5302 25880 5354 25889
rect 5302 25846 5311 25880
rect 5311 25846 5345 25880
rect 5345 25846 5354 25880
rect 5302 25837 5354 25846
rect 6454 25880 6506 25889
rect 6454 25846 6463 25880
rect 6463 25846 6497 25880
rect 6497 25846 6506 25880
rect 6454 25837 6506 25846
rect 7606 25880 7658 25889
rect 7606 25846 7615 25880
rect 7615 25846 7649 25880
rect 7649 25846 7658 25880
rect 7606 25837 7658 25846
rect 8662 25837 8714 25889
rect 9718 25880 9770 25889
rect 9718 25846 9727 25880
rect 9727 25846 9761 25880
rect 9761 25846 9770 25880
rect 9718 25837 9770 25846
rect 9814 25880 9866 25889
rect 9814 25846 9823 25880
rect 9823 25846 9857 25880
rect 9857 25846 9866 25880
rect 9814 25837 9866 25846
rect 1654 25763 1706 25815
rect 2422 25658 2474 25667
rect 2422 25624 2431 25658
rect 2431 25624 2465 25658
rect 2465 25624 2474 25658
rect 2422 25615 2474 25624
rect 3190 25658 3242 25667
rect 3190 25624 3199 25658
rect 3199 25624 3233 25658
rect 3233 25624 3242 25658
rect 3190 25615 3242 25624
rect 2710 25541 2762 25593
rect 5494 25658 5546 25667
rect 5494 25624 5503 25658
rect 5503 25624 5537 25658
rect 5537 25624 5546 25658
rect 5494 25615 5546 25624
rect 6454 25615 6506 25667
rect 7798 25658 7850 25667
rect 7798 25624 7807 25658
rect 7807 25624 7841 25658
rect 7841 25624 7850 25658
rect 7798 25615 7850 25624
rect 7894 25615 7946 25667
rect 9430 25658 9482 25667
rect 9430 25624 9439 25658
rect 9439 25624 9473 25658
rect 9473 25624 9482 25658
rect 9430 25615 9482 25624
rect 5686 25541 5738 25593
rect 7606 25541 7658 25593
rect 4966 25282 5018 25334
rect 5030 25282 5082 25334
rect 5094 25282 5146 25334
rect 5158 25282 5210 25334
rect 5222 25282 5274 25334
rect 5286 25282 5338 25334
rect 598 25171 650 25223
rect 10966 25171 11018 25223
rect 2518 24949 2570 25001
rect 8470 24949 8522 25001
rect 886 24875 938 24927
rect 5590 24875 5642 24927
rect 1966 24616 2018 24668
rect 2030 24616 2082 24668
rect 2094 24616 2146 24668
rect 2158 24616 2210 24668
rect 2222 24616 2274 24668
rect 2286 24616 2338 24668
rect 7966 24616 8018 24668
rect 8030 24616 8082 24668
rect 8094 24616 8146 24668
rect 8158 24616 8210 24668
rect 8222 24616 8274 24668
rect 8286 24616 8338 24668
rect 4966 23950 5018 24002
rect 5030 23950 5082 24002
rect 5094 23950 5146 24002
rect 5158 23950 5210 24002
rect 5222 23950 5274 24002
rect 5286 23950 5338 24002
rect 8470 23882 8522 23891
rect 8470 23848 8479 23882
rect 8479 23848 8513 23882
rect 8513 23848 8522 23882
rect 8470 23839 8522 23848
rect 9430 23839 9482 23891
rect 3862 23617 3914 23669
rect 6742 23617 6794 23669
rect 8758 23660 8810 23669
rect 8758 23626 8767 23660
rect 8767 23626 8801 23660
rect 8801 23626 8810 23660
rect 8758 23617 8810 23626
rect 5590 23543 5642 23595
rect 6070 23469 6122 23521
rect 790 23395 842 23447
rect 1966 23284 2018 23336
rect 2030 23284 2082 23336
rect 2094 23284 2146 23336
rect 2158 23284 2210 23336
rect 2222 23284 2274 23336
rect 2286 23284 2338 23336
rect 7966 23284 8018 23336
rect 8030 23284 8082 23336
rect 8094 23284 8146 23336
rect 8158 23284 8210 23336
rect 8222 23284 8274 23336
rect 8286 23284 8338 23336
rect 3862 23099 3914 23151
rect 6742 23099 6794 23151
rect 6070 23025 6122 23077
rect 5590 22994 5642 23003
rect 5590 22960 5599 22994
rect 5599 22960 5633 22994
rect 5633 22960 5642 22994
rect 5590 22951 5642 22960
rect 7606 22994 7658 23003
rect 7606 22960 7615 22994
rect 7615 22960 7649 22994
rect 7649 22960 7658 22994
rect 7606 22951 7658 22960
rect 9814 22994 9866 23003
rect 9814 22960 9823 22994
rect 9823 22960 9857 22994
rect 9857 22960 9866 22994
rect 9814 22951 9866 22960
rect 6550 22877 6602 22929
rect 8374 22877 8426 22929
rect 6070 22729 6122 22781
rect 8758 22803 8810 22855
rect 10102 22772 10154 22781
rect 10102 22738 10111 22772
rect 10111 22738 10145 22772
rect 10145 22738 10154 22772
rect 10102 22729 10154 22738
rect 4966 22618 5018 22670
rect 5030 22618 5082 22670
rect 5094 22618 5146 22670
rect 5158 22618 5210 22670
rect 5222 22618 5274 22670
rect 5286 22618 5338 22670
rect 9814 22550 9866 22559
rect 9814 22516 9823 22550
rect 9823 22516 9857 22550
rect 9857 22516 9866 22550
rect 9814 22507 9866 22516
rect 8470 22359 8522 22411
rect 1846 22328 1898 22337
rect 1846 22294 1855 22328
rect 1855 22294 1889 22328
rect 1889 22294 1898 22328
rect 1846 22285 1898 22294
rect 6550 22285 6602 22337
rect 8374 22285 8426 22337
rect 8662 22211 8714 22263
rect 886 22063 938 22115
rect 1966 21952 2018 22004
rect 2030 21952 2082 22004
rect 2094 21952 2146 22004
rect 2158 21952 2210 22004
rect 2222 21952 2274 22004
rect 2286 21952 2338 22004
rect 7966 21952 8018 22004
rect 8030 21952 8082 22004
rect 8094 21952 8146 22004
rect 8158 21952 8210 22004
rect 8222 21952 8274 22004
rect 8286 21952 8338 22004
rect 2422 21693 2474 21745
rect 3862 21736 3914 21745
rect 3862 21702 3871 21736
rect 3871 21702 3905 21736
rect 3905 21702 3914 21736
rect 3862 21693 3914 21702
rect 3286 21619 3338 21671
rect 8374 21619 8426 21671
rect 1846 21545 1898 21597
rect 4966 21286 5018 21338
rect 5030 21286 5082 21338
rect 5094 21286 5146 21338
rect 5158 21286 5210 21338
rect 5222 21286 5274 21338
rect 5286 21286 5338 21338
rect 7606 21027 7658 21079
rect 8374 20953 8426 21005
rect 8662 20879 8714 20931
rect 9814 20774 9866 20783
rect 9814 20740 9823 20774
rect 9823 20740 9857 20774
rect 9857 20740 9866 20774
rect 9814 20731 9866 20740
rect 1966 20620 2018 20672
rect 2030 20620 2082 20672
rect 2094 20620 2146 20672
rect 2158 20620 2210 20672
rect 2222 20620 2274 20672
rect 2286 20620 2338 20672
rect 7966 20620 8018 20672
rect 8030 20620 8082 20672
rect 8094 20620 8146 20672
rect 8158 20620 8210 20672
rect 8222 20620 8274 20672
rect 8286 20620 8338 20672
rect 1846 20509 1898 20561
rect 5590 20509 5642 20561
rect 7894 20509 7946 20561
rect 2422 20361 2474 20413
rect 5398 20404 5450 20413
rect 5398 20370 5407 20404
rect 5407 20370 5441 20404
rect 5441 20370 5450 20404
rect 5398 20361 5450 20370
rect 6070 20361 6122 20413
rect 3286 20330 3338 20339
rect 3286 20296 3295 20330
rect 3295 20296 3329 20330
rect 3329 20296 3338 20330
rect 3286 20287 3338 20296
rect 3670 20330 3722 20339
rect 3670 20296 3679 20330
rect 3679 20296 3713 20330
rect 3713 20296 3722 20330
rect 3670 20287 3722 20296
rect 5878 20287 5930 20339
rect 9814 20330 9866 20339
rect 9814 20296 9823 20330
rect 9823 20296 9857 20330
rect 9857 20296 9866 20330
rect 9814 20287 9866 20296
rect 10102 20182 10154 20191
rect 10102 20148 10111 20182
rect 10111 20148 10145 20182
rect 10145 20148 10154 20182
rect 10102 20139 10154 20148
rect 4966 19954 5018 20006
rect 5030 19954 5082 20006
rect 5094 19954 5146 20006
rect 5158 19954 5210 20006
rect 5222 19954 5274 20006
rect 5286 19954 5338 20006
rect 1558 19886 1610 19895
rect 1558 19852 1567 19886
rect 1567 19852 1601 19886
rect 1601 19852 1610 19886
rect 1558 19843 1610 19852
rect 7894 19695 7946 19747
rect 1750 19621 1802 19673
rect 3670 19621 3722 19673
rect 8374 19621 8426 19673
rect 7894 19547 7946 19599
rect 8662 19547 8714 19599
rect 9814 19442 9866 19451
rect 9814 19408 9823 19442
rect 9823 19408 9857 19442
rect 9857 19408 9866 19442
rect 9814 19399 9866 19408
rect 1966 19288 2018 19340
rect 2030 19288 2082 19340
rect 2094 19288 2146 19340
rect 2158 19288 2210 19340
rect 2222 19288 2274 19340
rect 2286 19288 2338 19340
rect 7966 19288 8018 19340
rect 8030 19288 8082 19340
rect 8094 19288 8146 19340
rect 8158 19288 8210 19340
rect 8222 19288 8274 19340
rect 8286 19288 8338 19340
rect 1750 19220 1802 19229
rect 1750 19186 1759 19220
rect 1759 19186 1793 19220
rect 1793 19186 1802 19220
rect 1750 19177 1802 19186
rect 2422 19029 2474 19081
rect 4438 19029 4490 19081
rect 5398 19103 5450 19155
rect 6070 19103 6122 19155
rect 5590 19029 5642 19081
rect 3286 18998 3338 19007
rect 3286 18964 3295 18998
rect 3295 18964 3329 18998
rect 3329 18964 3338 18998
rect 3286 18955 3338 18964
rect 4150 18955 4202 19007
rect 7798 18733 7850 18785
rect 4966 18622 5018 18674
rect 5030 18622 5082 18674
rect 5094 18622 5146 18674
rect 5158 18622 5210 18674
rect 5222 18622 5274 18674
rect 5286 18622 5338 18674
rect 1558 18554 1610 18563
rect 1558 18520 1567 18554
rect 1567 18520 1601 18554
rect 1601 18520 1610 18554
rect 1558 18511 1610 18520
rect 6454 18363 6506 18415
rect 1750 18289 1802 18341
rect 4150 18289 4202 18341
rect 7894 18289 7946 18341
rect 8662 18215 8714 18267
rect 9718 18110 9770 18119
rect 9718 18076 9727 18110
rect 9727 18076 9761 18110
rect 9761 18076 9770 18110
rect 9718 18067 9770 18076
rect 1966 17956 2018 18008
rect 2030 17956 2082 18008
rect 2094 17956 2146 18008
rect 2158 17956 2210 18008
rect 2222 17956 2274 18008
rect 2286 17956 2338 18008
rect 7966 17956 8018 18008
rect 8030 17956 8082 18008
rect 8094 17956 8146 18008
rect 8158 17956 8210 18008
rect 8222 17956 8274 18008
rect 8286 17956 8338 18008
rect 1750 17888 1802 17897
rect 1750 17854 1759 17888
rect 1759 17854 1793 17888
rect 1793 17854 1802 17888
rect 1750 17845 1802 17854
rect 6454 17888 6506 17897
rect 6454 17854 6463 17888
rect 6463 17854 6497 17888
rect 6497 17854 6506 17888
rect 6454 17845 6506 17854
rect 2422 17697 2474 17749
rect 4438 17740 4490 17749
rect 4438 17706 4447 17740
rect 4447 17706 4481 17740
rect 4481 17706 4490 17740
rect 4438 17697 4490 17706
rect 5590 17771 5642 17823
rect 10102 17814 10154 17823
rect 10102 17780 10111 17814
rect 10111 17780 10145 17814
rect 10145 17780 10154 17814
rect 10102 17771 10154 17780
rect 2806 17623 2858 17675
rect 3286 17666 3338 17675
rect 3286 17632 3295 17666
rect 3295 17632 3329 17666
rect 3329 17632 3338 17666
rect 3286 17623 3338 17632
rect 4246 17623 4298 17675
rect 9814 17666 9866 17675
rect 9814 17632 9823 17666
rect 9823 17632 9857 17666
rect 9857 17632 9866 17666
rect 9814 17623 9866 17632
rect 4966 17290 5018 17342
rect 5030 17290 5082 17342
rect 5094 17290 5146 17342
rect 5158 17290 5210 17342
rect 5222 17290 5274 17342
rect 5286 17290 5338 17342
rect 1270 17179 1322 17231
rect 1750 16957 1802 17009
rect 4246 17031 4298 17083
rect 7798 17074 7850 17083
rect 7798 17040 7807 17074
rect 7807 17040 7841 17074
rect 7841 17040 7850 17074
rect 7798 17031 7850 17040
rect 3958 17000 4010 17009
rect 3958 16966 3967 17000
rect 3967 16966 4001 17000
rect 4001 16966 4010 17000
rect 3958 16957 4010 16966
rect 7894 16957 7946 17009
rect 2902 16809 2954 16861
rect 5590 16883 5642 16935
rect 8758 16883 8810 16935
rect 4438 16809 4490 16861
rect 5590 16778 5642 16787
rect 5590 16744 5599 16778
rect 5599 16744 5633 16778
rect 5633 16744 5642 16778
rect 5590 16735 5642 16744
rect 9814 16778 9866 16787
rect 9814 16744 9823 16778
rect 9823 16744 9857 16778
rect 9857 16744 9866 16778
rect 9814 16735 9866 16744
rect 1966 16624 2018 16676
rect 2030 16624 2082 16676
rect 2094 16624 2146 16676
rect 2158 16624 2210 16676
rect 2222 16624 2274 16676
rect 2286 16624 2338 16676
rect 7966 16624 8018 16676
rect 8030 16624 8082 16676
rect 8094 16624 8146 16676
rect 8158 16624 8210 16676
rect 8222 16624 8274 16676
rect 8286 16624 8338 16676
rect 1750 16556 1802 16565
rect 1750 16522 1759 16556
rect 1759 16522 1793 16556
rect 1793 16522 1802 16556
rect 1750 16513 1802 16522
rect 2806 16365 2858 16417
rect 3286 16334 3338 16343
rect 3286 16300 3295 16334
rect 3295 16300 3329 16334
rect 3329 16300 3338 16334
rect 3286 16291 3338 16300
rect 2998 16217 3050 16269
rect 3958 16217 4010 16269
rect 4966 15958 5018 16010
rect 5030 15958 5082 16010
rect 5094 15958 5146 16010
rect 5158 15958 5210 16010
rect 5222 15958 5274 16010
rect 5286 15958 5338 16010
rect 790 15699 842 15751
rect 2902 15742 2954 15751
rect 2902 15708 2911 15742
rect 2911 15708 2945 15742
rect 2945 15708 2954 15742
rect 2902 15699 2954 15708
rect 5590 15699 5642 15751
rect 2998 15625 3050 15677
rect 3670 15625 3722 15677
rect 7894 15668 7946 15677
rect 7894 15634 7903 15668
rect 7903 15634 7937 15668
rect 7937 15634 7946 15668
rect 7894 15625 7946 15634
rect 9814 15668 9866 15677
rect 9814 15634 9823 15668
rect 9823 15634 9857 15668
rect 9857 15634 9866 15668
rect 9814 15625 9866 15634
rect 2806 15551 2858 15603
rect 8758 15551 8810 15603
rect 5398 15403 5450 15455
rect 5686 15403 5738 15455
rect 9814 15403 9866 15455
rect 10102 15446 10154 15455
rect 10102 15412 10111 15446
rect 10111 15412 10145 15446
rect 10145 15412 10154 15446
rect 10102 15403 10154 15412
rect 1966 15292 2018 15344
rect 2030 15292 2082 15344
rect 2094 15292 2146 15344
rect 2158 15292 2210 15344
rect 2222 15292 2274 15344
rect 2286 15292 2338 15344
rect 7966 15292 8018 15344
rect 8030 15292 8082 15344
rect 8094 15292 8146 15344
rect 8158 15292 8210 15344
rect 8222 15292 8274 15344
rect 8286 15292 8338 15344
rect 2806 15033 2858 15085
rect 3286 15002 3338 15011
rect 3286 14968 3295 15002
rect 3295 14968 3329 15002
rect 3329 14968 3338 15002
rect 3286 14959 3338 14968
rect 3670 14928 3722 14937
rect 3670 14894 3679 14928
rect 3679 14894 3713 14928
rect 3713 14894 3722 14928
rect 3670 14885 3722 14894
rect 2998 14737 3050 14789
rect 3382 14737 3434 14789
rect 4966 14626 5018 14678
rect 5030 14626 5082 14678
rect 5094 14626 5146 14678
rect 5158 14626 5210 14678
rect 5222 14626 5274 14678
rect 5286 14626 5338 14678
rect 2806 14441 2858 14493
rect 5398 14441 5450 14493
rect 3670 14293 3722 14345
rect 4246 14293 4298 14345
rect 7894 14336 7946 14345
rect 7894 14302 7903 14336
rect 7903 14302 7937 14336
rect 7937 14302 7946 14336
rect 7894 14293 7946 14302
rect 8374 14293 8426 14345
rect 790 14219 842 14271
rect 2902 14219 2954 14271
rect 4630 14219 4682 14271
rect 8758 14219 8810 14271
rect 7030 14071 7082 14123
rect 9526 14114 9578 14123
rect 9526 14080 9535 14114
rect 9535 14080 9569 14114
rect 9569 14080 9578 14114
rect 9526 14071 9578 14080
rect 1966 13960 2018 14012
rect 2030 13960 2082 14012
rect 2094 13960 2146 14012
rect 2158 13960 2210 14012
rect 2222 13960 2274 14012
rect 2286 13960 2338 14012
rect 7966 13960 8018 14012
rect 8030 13960 8082 14012
rect 8094 13960 8146 14012
rect 8158 13960 8210 14012
rect 8222 13960 8274 14012
rect 8286 13960 8338 14012
rect 4630 13701 4682 13753
rect 7222 13775 7274 13827
rect 4150 13627 4202 13679
rect 9718 13627 9770 13679
rect 2902 13553 2954 13605
rect 6166 13553 6218 13605
rect 7510 13405 7562 13457
rect 10102 13448 10154 13457
rect 10102 13414 10111 13448
rect 10111 13414 10145 13448
rect 10145 13414 10154 13448
rect 10102 13405 10154 13414
rect 4966 13294 5018 13346
rect 5030 13294 5082 13346
rect 5094 13294 5146 13346
rect 5158 13294 5210 13346
rect 5222 13294 5274 13346
rect 5286 13294 5338 13346
rect 2710 13109 2762 13161
rect 4342 13109 4394 13161
rect 1558 13004 1610 13013
rect 1558 12970 1567 13004
rect 1567 12970 1601 13004
rect 1601 12970 1610 13004
rect 1558 12961 1610 12970
rect 1462 12887 1514 12939
rect 2902 12961 2954 13013
rect 3382 13004 3434 13013
rect 3382 12970 3391 13004
rect 3391 12970 3425 13004
rect 3425 12970 3434 13004
rect 3382 12961 3434 12970
rect 5494 12961 5546 13013
rect 8374 12961 8426 13013
rect 2806 12887 2858 12939
rect 8758 12887 8810 12939
rect 9718 12782 9770 12791
rect 9718 12748 9727 12782
rect 9727 12748 9761 12782
rect 9761 12748 9770 12782
rect 9718 12739 9770 12748
rect 1966 12628 2018 12680
rect 2030 12628 2082 12680
rect 2094 12628 2146 12680
rect 2158 12628 2210 12680
rect 2222 12628 2274 12680
rect 2286 12628 2338 12680
rect 7966 12628 8018 12680
rect 8030 12628 8082 12680
rect 8094 12628 8146 12680
rect 8158 12628 8210 12680
rect 8222 12628 8274 12680
rect 8286 12628 8338 12680
rect 2806 12369 2858 12421
rect 6166 12412 6218 12421
rect 6166 12378 6175 12412
rect 6175 12378 6209 12412
rect 6209 12378 6218 12412
rect 6166 12369 6218 12378
rect 7222 12369 7274 12421
rect 1846 12295 1898 12347
rect 3286 12295 3338 12347
rect 6550 12338 6602 12347
rect 6550 12304 6559 12338
rect 6559 12304 6593 12338
rect 6593 12304 6602 12338
rect 6550 12295 6602 12304
rect 1462 12221 1514 12273
rect 3670 12073 3722 12125
rect 4246 12073 4298 12125
rect 10198 12073 10250 12125
rect 4966 11962 5018 12014
rect 5030 11962 5082 12014
rect 5094 11962 5146 12014
rect 5158 11962 5210 12014
rect 5222 11962 5274 12014
rect 5286 11962 5338 12014
rect 3094 11851 3146 11903
rect 7702 11851 7754 11903
rect 1462 11703 1514 11755
rect 2710 11629 2762 11681
rect 5878 11629 5930 11681
rect 2998 11481 3050 11533
rect 1558 11450 1610 11459
rect 1558 11416 1567 11450
rect 1567 11416 1601 11450
rect 1601 11416 1610 11450
rect 1558 11407 1610 11416
rect 2806 11407 2858 11459
rect 6166 11555 6218 11607
rect 7222 11555 7274 11607
rect 8470 11598 8522 11607
rect 8470 11564 8479 11598
rect 8479 11564 8513 11598
rect 8513 11564 8522 11598
rect 8470 11555 8522 11564
rect 1966 11296 2018 11348
rect 2030 11296 2082 11348
rect 2094 11296 2146 11348
rect 2158 11296 2210 11348
rect 2222 11296 2274 11348
rect 2286 11296 2338 11348
rect 7966 11296 8018 11348
rect 8030 11296 8082 11348
rect 8094 11296 8146 11348
rect 8158 11296 8210 11348
rect 8222 11296 8274 11348
rect 8286 11296 8338 11348
rect 2518 11185 2570 11237
rect 7798 11185 7850 11237
rect 2998 11111 3050 11163
rect 2806 11037 2858 11089
rect 1942 11006 1994 11015
rect 1942 10972 1951 11006
rect 1951 10972 1985 11006
rect 1985 10972 1994 11006
rect 1942 10963 1994 10972
rect 6166 11037 6218 11089
rect 7222 11037 7274 11089
rect 4246 11006 4298 11015
rect 4246 10972 4255 11006
rect 4255 10972 4289 11006
rect 4289 10972 4298 11006
rect 4246 10963 4298 10972
rect 6742 10963 6794 11015
rect 9814 11006 9866 11015
rect 9814 10972 9823 11006
rect 9823 10972 9857 11006
rect 9857 10972 9866 11006
rect 9814 10963 9866 10972
rect 2902 10889 2954 10941
rect 4438 10741 4490 10793
rect 9430 10741 9482 10793
rect 10102 10784 10154 10793
rect 10102 10750 10111 10784
rect 10111 10750 10145 10784
rect 10145 10750 10154 10784
rect 10102 10741 10154 10750
rect 4966 10630 5018 10682
rect 5030 10630 5082 10682
rect 5094 10630 5146 10682
rect 5158 10630 5210 10682
rect 5222 10630 5274 10682
rect 5286 10630 5338 10682
rect 4342 10562 4394 10571
rect 4342 10528 4351 10562
rect 4351 10528 4385 10562
rect 4385 10528 4394 10562
rect 4342 10519 4394 10528
rect 2998 10371 3050 10423
rect 7702 10414 7754 10423
rect 7702 10380 7711 10414
rect 7711 10380 7745 10414
rect 7745 10380 7754 10414
rect 7702 10371 7754 10380
rect 1942 10297 1994 10349
rect 2710 10340 2762 10349
rect 2710 10306 2719 10340
rect 2719 10306 2753 10340
rect 2753 10306 2762 10340
rect 2710 10297 2762 10306
rect 3670 10297 3722 10349
rect 8374 10297 8426 10349
rect 8758 10223 8810 10275
rect 2710 10149 2762 10201
rect 1558 10118 1610 10127
rect 1558 10084 1567 10118
rect 1567 10084 1601 10118
rect 1601 10084 1610 10118
rect 1558 10075 1610 10084
rect 9814 10075 9866 10127
rect 1966 9964 2018 10016
rect 2030 9964 2082 10016
rect 2094 9964 2146 10016
rect 2158 9964 2210 10016
rect 2222 9964 2274 10016
rect 2286 9964 2338 10016
rect 7966 9964 8018 10016
rect 8030 9964 8082 10016
rect 8094 9964 8146 10016
rect 8158 9964 8210 10016
rect 8222 9964 8274 10016
rect 8286 9964 8338 10016
rect 4966 9298 5018 9350
rect 5030 9298 5082 9350
rect 5094 9298 5146 9350
rect 5158 9298 5210 9350
rect 5222 9298 5274 9350
rect 5286 9298 5338 9350
rect 7798 9082 7850 9091
rect 7798 9048 7807 9082
rect 7807 9048 7841 9082
rect 7841 9048 7850 9082
rect 7798 9039 7850 9048
rect 8374 8965 8426 9017
rect 1654 8934 1706 8943
rect 1654 8900 1663 8934
rect 1663 8900 1697 8934
rect 1697 8900 1706 8934
rect 1654 8891 1706 8900
rect 2902 8891 2954 8943
rect 8758 8891 8810 8943
rect 10006 8743 10058 8795
rect 1966 8632 2018 8684
rect 2030 8632 2082 8684
rect 2094 8632 2146 8684
rect 2158 8632 2210 8684
rect 2222 8632 2274 8684
rect 2286 8632 2338 8684
rect 7966 8632 8018 8684
rect 8030 8632 8082 8684
rect 8094 8632 8146 8684
rect 8158 8632 8210 8684
rect 8222 8632 8274 8684
rect 8286 8632 8338 8684
rect 1750 8564 1802 8573
rect 1750 8530 1759 8564
rect 1759 8530 1793 8564
rect 1793 8530 1802 8564
rect 1750 8521 1802 8530
rect 6262 8373 6314 8425
rect 7702 8342 7754 8351
rect 7702 8308 7711 8342
rect 7711 8308 7745 8342
rect 7745 8308 7754 8342
rect 7702 8299 7754 8308
rect 9526 8299 9578 8351
rect 10102 8342 10154 8351
rect 10102 8308 10111 8342
rect 10111 8308 10145 8342
rect 10145 8308 10154 8342
rect 10102 8299 10154 8308
rect 1654 8268 1706 8277
rect 1654 8234 1663 8268
rect 1663 8234 1697 8268
rect 1697 8234 1706 8268
rect 1654 8225 1706 8234
rect 4966 7966 5018 8018
rect 5030 7966 5082 8018
rect 5094 7966 5146 8018
rect 5158 7966 5210 8018
rect 5222 7966 5274 8018
rect 5286 7966 5338 8018
rect 3670 7898 3722 7907
rect 3670 7864 3679 7898
rect 3679 7864 3713 7898
rect 3713 7864 3722 7898
rect 3670 7855 3722 7864
rect 6358 7855 6410 7907
rect 1558 7707 1610 7759
rect 1846 7707 1898 7759
rect 8374 7707 8426 7759
rect 1750 7633 1802 7685
rect 2806 7633 2858 7685
rect 2710 7559 2762 7611
rect 1462 7485 1514 7537
rect 1750 7485 1802 7537
rect 6838 7454 6890 7463
rect 6838 7420 6847 7454
rect 6847 7420 6881 7454
rect 6881 7420 6890 7454
rect 6838 7411 6890 7420
rect 1966 7300 2018 7352
rect 2030 7300 2082 7352
rect 2094 7300 2146 7352
rect 2158 7300 2210 7352
rect 2222 7300 2274 7352
rect 2286 7300 2338 7352
rect 7966 7300 8018 7352
rect 8030 7300 8082 7352
rect 8094 7300 8146 7352
rect 8158 7300 8210 7352
rect 8222 7300 8274 7352
rect 8286 7300 8338 7352
rect 1558 7189 1610 7241
rect 8374 7189 8426 7241
rect 2806 6967 2858 7019
rect 2710 6893 2762 6945
rect 6838 7041 6890 7093
rect 6262 7010 6314 7019
rect 6262 6976 6271 7010
rect 6271 6976 6305 7010
rect 6305 6976 6314 7010
rect 6262 6967 6314 6976
rect 6454 6967 6506 7019
rect 9526 6967 9578 7019
rect 8854 6893 8906 6945
rect 4966 6634 5018 6686
rect 5030 6634 5082 6686
rect 5094 6634 5146 6686
rect 5158 6634 5210 6686
rect 5222 6634 5274 6686
rect 5286 6634 5338 6686
rect 1750 6566 1802 6575
rect 1750 6532 1759 6566
rect 1759 6532 1793 6566
rect 1793 6532 1802 6566
rect 1750 6523 1802 6532
rect 5878 6523 5930 6575
rect 6358 6523 6410 6575
rect 6070 6449 6122 6501
rect 2806 6375 2858 6427
rect 5974 6375 6026 6427
rect 8854 6418 8906 6427
rect 8854 6384 8863 6418
rect 8863 6384 8897 6418
rect 8897 6384 8906 6418
rect 8854 6375 8906 6384
rect 2710 6153 2762 6205
rect 3766 6270 3818 6279
rect 3766 6236 3775 6270
rect 3775 6236 3809 6270
rect 3809 6236 3818 6270
rect 3766 6227 3818 6236
rect 5686 6301 5738 6353
rect 6454 6301 6506 6353
rect 7798 6301 7850 6353
rect 8278 6301 8330 6353
rect 8470 6301 8522 6353
rect 9046 6344 9098 6353
rect 9046 6310 9055 6344
rect 9055 6310 9089 6344
rect 9089 6310 9098 6344
rect 9046 6301 9098 6310
rect 9334 6344 9386 6353
rect 9334 6310 9343 6344
rect 9343 6310 9377 6344
rect 9377 6310 9386 6344
rect 9334 6301 9386 6310
rect 9814 6344 9866 6353
rect 9814 6310 9823 6344
rect 9823 6310 9857 6344
rect 9857 6310 9866 6344
rect 9814 6301 9866 6310
rect 5686 6153 5738 6205
rect 6838 6079 6890 6131
rect 8278 6153 8330 6205
rect 8374 6079 8426 6131
rect 8566 6079 8618 6131
rect 10102 6122 10154 6131
rect 10102 6088 10111 6122
rect 10111 6088 10145 6122
rect 10145 6088 10154 6122
rect 10102 6079 10154 6088
rect 1966 5968 2018 6020
rect 2030 5968 2082 6020
rect 2094 5968 2146 6020
rect 2158 5968 2210 6020
rect 2222 5968 2274 6020
rect 2286 5968 2338 6020
rect 7966 5968 8018 6020
rect 8030 5968 8082 6020
rect 8094 5968 8146 6020
rect 8158 5968 8210 6020
rect 8222 5968 8274 6020
rect 8286 5968 8338 6020
rect 1558 5709 1610 5761
rect 2710 5709 2762 5761
rect 7702 5709 7754 5761
rect 8374 5709 8426 5761
rect 9526 5752 9578 5761
rect 9526 5718 9535 5752
rect 9535 5718 9569 5752
rect 9569 5718 9578 5752
rect 9526 5709 9578 5718
rect 1654 5561 1706 5613
rect 2902 5561 2954 5613
rect 4822 5604 4874 5613
rect 4822 5570 4831 5604
rect 4831 5570 4865 5604
rect 4865 5570 4874 5604
rect 4822 5561 4874 5570
rect 6070 5635 6122 5687
rect 6358 5678 6410 5687
rect 6358 5644 6367 5678
rect 6367 5644 6401 5678
rect 6401 5644 6410 5678
rect 6358 5635 6410 5644
rect 5110 5604 5162 5613
rect 5110 5570 5119 5604
rect 5119 5570 5153 5604
rect 5153 5570 5162 5604
rect 5110 5561 5162 5570
rect 5686 5561 5738 5613
rect 6070 5487 6122 5539
rect 9046 5635 9098 5687
rect 9622 5678 9674 5687
rect 9622 5644 9631 5678
rect 9631 5644 9665 5678
rect 9665 5644 9674 5678
rect 9622 5635 9674 5644
rect 9142 5561 9194 5613
rect 2902 5413 2954 5465
rect 5974 5413 6026 5465
rect 8374 5413 8426 5465
rect 4966 5302 5018 5354
rect 5030 5302 5082 5354
rect 5094 5302 5146 5354
rect 5158 5302 5210 5354
rect 5222 5302 5274 5354
rect 5286 5302 5338 5354
rect 5686 5191 5738 5243
rect 9046 5191 9098 5243
rect 9622 5191 9674 5243
rect 1654 5086 1706 5095
rect 1654 5052 1663 5086
rect 1663 5052 1697 5086
rect 1697 5052 1706 5086
rect 1654 5043 1706 5052
rect 1846 5043 1898 5095
rect 6838 5086 6890 5095
rect 6838 5052 6847 5086
rect 6847 5052 6881 5086
rect 6881 5052 6890 5086
rect 6838 5043 6890 5052
rect 8374 5043 8426 5095
rect 2710 4895 2762 4947
rect 5782 4938 5834 4947
rect 5782 4904 5791 4938
rect 5791 4904 5825 4938
rect 5825 4904 5834 4938
rect 5782 4895 5834 4904
rect 6454 5012 6506 5021
rect 6454 4978 6463 5012
rect 6463 4978 6497 5012
rect 6497 4978 6506 5012
rect 6454 4969 6506 4978
rect 7798 4969 7850 5021
rect 9142 5086 9194 5095
rect 9142 5052 9151 5086
rect 9151 5052 9185 5086
rect 9185 5052 9194 5086
rect 9142 5043 9194 5052
rect 6550 4895 6602 4947
rect 3286 4747 3338 4799
rect 4630 4790 4682 4799
rect 4630 4756 4639 4790
rect 4639 4756 4673 4790
rect 4673 4756 4682 4790
rect 4630 4747 4682 4756
rect 8470 4747 8522 4799
rect 1966 4636 2018 4688
rect 2030 4636 2082 4688
rect 2094 4636 2146 4688
rect 2158 4636 2210 4688
rect 2222 4636 2274 4688
rect 2286 4636 2338 4688
rect 7966 4636 8018 4688
rect 8030 4636 8082 4688
rect 8094 4636 8146 4688
rect 8158 4636 8210 4688
rect 8222 4636 8274 4688
rect 8286 4636 8338 4688
rect 5782 4525 5834 4577
rect 8374 4525 8426 4577
rect 2710 4377 2762 4429
rect 3766 4303 3818 4355
rect 4630 4303 4682 4355
rect 6070 4377 6122 4429
rect 5974 4346 6026 4355
rect 5974 4312 5983 4346
rect 5983 4312 6017 4346
rect 6017 4312 6026 4346
rect 5974 4303 6026 4312
rect 8566 4377 8618 4429
rect 2998 4229 3050 4281
rect 6550 4303 6602 4355
rect 7126 4303 7178 4355
rect 7702 4303 7754 4355
rect 8470 4272 8522 4281
rect 8470 4238 8479 4272
rect 8479 4238 8513 4272
rect 8513 4238 8522 4272
rect 8470 4229 8522 4238
rect 7798 4155 7850 4207
rect 8086 4155 8138 4207
rect 9334 4155 9386 4207
rect 1654 4124 1706 4133
rect 1654 4090 1663 4124
rect 1663 4090 1697 4124
rect 1697 4090 1706 4124
rect 1654 4081 1706 4090
rect 6358 4124 6410 4133
rect 6358 4090 6367 4124
rect 6367 4090 6401 4124
rect 6401 4090 6410 4124
rect 6358 4081 6410 4090
rect 8758 4081 8810 4133
rect 4966 3970 5018 4022
rect 5030 3970 5082 4022
rect 5094 3970 5146 4022
rect 5158 3970 5210 4022
rect 5222 3970 5274 4022
rect 5286 3970 5338 4022
rect 5878 3902 5930 3911
rect 5878 3868 5887 3902
rect 5887 3868 5921 3902
rect 5921 3868 5930 3902
rect 5878 3859 5930 3868
rect 4822 3785 4874 3837
rect 8086 3902 8138 3911
rect 8086 3868 8095 3902
rect 8095 3868 8129 3902
rect 8129 3868 8138 3902
rect 8086 3859 8138 3868
rect 8758 3785 8810 3837
rect 6166 3711 6218 3763
rect 6358 3711 6410 3763
rect 886 3637 938 3689
rect 6550 3680 6602 3689
rect 6550 3646 6559 3680
rect 6559 3646 6593 3680
rect 6593 3646 6602 3680
rect 6550 3637 6602 3646
rect 7510 3637 7562 3689
rect 9430 3680 9482 3689
rect 9430 3646 9439 3680
rect 9439 3646 9473 3680
rect 9473 3646 9482 3680
rect 9430 3637 9482 3646
rect 9718 3637 9770 3689
rect 10102 3606 10154 3615
rect 10102 3572 10111 3606
rect 10111 3572 10145 3606
rect 10145 3572 10154 3606
rect 10102 3563 10154 3572
rect 7510 3489 7562 3541
rect 10966 3415 11018 3467
rect 1966 3304 2018 3356
rect 2030 3304 2082 3356
rect 2094 3304 2146 3356
rect 2158 3304 2210 3356
rect 2222 3304 2274 3356
rect 2286 3304 2338 3356
rect 7966 3304 8018 3356
rect 8030 3304 8082 3356
rect 8094 3304 8146 3356
rect 8158 3304 8210 3356
rect 8222 3304 8274 3356
rect 8286 3304 8338 3356
rect 7894 3193 7946 3245
rect 598 3045 650 3097
rect 1654 2971 1706 3023
rect 4630 3045 4682 3097
rect 6550 3045 6602 3097
rect 2902 3014 2954 3023
rect 2902 2980 2911 3014
rect 2911 2980 2945 3014
rect 2945 2980 2954 3014
rect 2902 2971 2954 2980
rect 3286 3014 3338 3023
rect 3286 2980 3295 3014
rect 3295 2980 3329 3014
rect 3329 2980 3338 3014
rect 3286 2971 3338 2980
rect 4438 3014 4490 3023
rect 4438 2980 4447 3014
rect 4447 2980 4481 3014
rect 4481 2980 4490 3014
rect 4438 2971 4490 2980
rect 5494 3014 5546 3023
rect 5494 2980 5503 3014
rect 5503 2980 5537 3014
rect 5537 2980 5546 3014
rect 5494 2971 5546 2980
rect 7030 2971 7082 3023
rect 7126 3014 7178 3023
rect 7126 2980 7135 3014
rect 7135 2980 7169 3014
rect 7169 2980 7178 3014
rect 7126 2971 7178 2980
rect 10006 2971 10058 3023
rect 10198 2971 10250 3023
rect 1846 2940 1898 2949
rect 1846 2906 1855 2940
rect 1855 2906 1889 2940
rect 1889 2906 1898 2940
rect 1846 2897 1898 2906
rect 2998 2940 3050 2949
rect 2998 2906 3007 2940
rect 3007 2906 3041 2940
rect 3041 2906 3050 2940
rect 2998 2897 3050 2906
rect 4150 2940 4202 2949
rect 4150 2906 4159 2940
rect 4159 2906 4193 2940
rect 4193 2906 4202 2940
rect 4150 2897 4202 2906
rect 5398 2897 5450 2949
rect 6454 2940 6506 2949
rect 6454 2906 6463 2940
rect 6463 2906 6497 2940
rect 6497 2906 6506 2940
rect 6454 2897 6506 2906
rect 8854 2897 8906 2949
rect 9718 2940 9770 2949
rect 9718 2906 9727 2940
rect 9727 2906 9761 2940
rect 9761 2906 9770 2940
rect 9718 2897 9770 2906
rect 9814 2940 9866 2949
rect 9814 2906 9823 2940
rect 9823 2906 9857 2940
rect 9857 2906 9866 2940
rect 9814 2897 9866 2906
rect 2230 2792 2282 2801
rect 2230 2758 2239 2792
rect 2239 2758 2273 2792
rect 2273 2758 2282 2792
rect 2230 2749 2282 2758
rect 4966 2638 5018 2690
rect 5030 2638 5082 2690
rect 5094 2638 5146 2690
rect 5158 2638 5210 2690
rect 5222 2638 5274 2690
rect 5286 2638 5338 2690
<< metal2 >>
rect 596 28074 652 28874
rect 1748 28074 1804 28874
rect 2900 28208 2956 28874
rect 4052 28208 4108 28874
rect 5204 28208 5260 28874
rect 6356 28208 6412 28874
rect 7508 28208 7564 28874
rect 2900 28180 3038 28208
rect 2900 28074 2956 28180
rect 610 25229 638 28074
rect 1652 26150 1708 26159
rect 1652 26085 1708 26094
rect 1666 25821 1694 26085
rect 1762 25895 1790 28074
rect 1964 26002 2340 26011
rect 2020 26000 2044 26002
rect 2100 26000 2124 26002
rect 2180 26000 2204 26002
rect 2260 26000 2284 26002
rect 2020 25948 2030 26000
rect 2274 25948 2284 26000
rect 2020 25946 2044 25948
rect 2100 25946 2124 25948
rect 2180 25946 2204 25948
rect 2260 25946 2284 25948
rect 1964 25937 2340 25946
rect 3010 25895 3038 28180
rect 4052 28180 4190 28208
rect 4052 28074 4108 28180
rect 4162 25895 4190 28180
rect 5204 28180 5342 28208
rect 5204 28074 5260 28180
rect 5314 25895 5342 28180
rect 6356 28180 6494 28208
rect 6356 28074 6412 28180
rect 6466 25895 6494 28180
rect 7508 28180 7646 28208
rect 7508 28074 7564 28180
rect 7618 25895 7646 28180
rect 8660 28074 8716 28874
rect 9812 28074 9868 28874
rect 10964 28074 11020 28874
rect 7964 26002 8340 26011
rect 8020 26000 8044 26002
rect 8100 26000 8124 26002
rect 8180 26000 8204 26002
rect 8260 26000 8284 26002
rect 8020 25948 8030 26000
rect 8274 25948 8284 26000
rect 8020 25946 8044 25948
rect 8100 25946 8124 25948
rect 8180 25946 8204 25948
rect 8260 25946 8284 25948
rect 7964 25937 8340 25946
rect 8674 25895 8702 28074
rect 9716 27334 9772 27343
rect 9716 27269 9772 27278
rect 9730 25895 9758 27269
rect 9826 25895 9854 28074
rect 1750 25889 1802 25895
rect 1750 25831 1802 25837
rect 2998 25889 3050 25895
rect 2998 25831 3050 25837
rect 4150 25889 4202 25895
rect 4150 25831 4202 25837
rect 5302 25889 5354 25895
rect 5302 25831 5354 25837
rect 6454 25889 6506 25895
rect 6454 25831 6506 25837
rect 7606 25889 7658 25895
rect 7606 25831 7658 25837
rect 8662 25889 8714 25895
rect 8662 25831 8714 25837
rect 9718 25889 9770 25895
rect 9718 25831 9770 25837
rect 9814 25889 9866 25895
rect 9814 25831 9866 25837
rect 1654 25815 1706 25821
rect 1654 25757 1706 25763
rect 2422 25667 2474 25673
rect 2422 25609 2474 25615
rect 3190 25667 3242 25673
rect 3190 25609 3242 25615
rect 5494 25667 5546 25673
rect 5494 25609 5546 25615
rect 6454 25667 6506 25673
rect 6454 25609 6506 25615
rect 7798 25667 7850 25673
rect 7798 25609 7850 25615
rect 7894 25667 7946 25673
rect 7894 25609 7946 25615
rect 9430 25667 9482 25673
rect 9430 25609 9482 25615
rect 598 25223 650 25229
rect 598 25165 650 25171
rect 886 24927 938 24933
rect 886 24869 938 24875
rect 898 24679 926 24869
rect 884 24670 940 24679
rect 884 24605 940 24614
rect 1964 24670 2340 24679
rect 2020 24668 2044 24670
rect 2100 24668 2124 24670
rect 2180 24668 2204 24670
rect 2260 24668 2284 24670
rect 2020 24616 2030 24668
rect 2274 24616 2284 24668
rect 2020 24614 2044 24616
rect 2100 24614 2124 24616
rect 2180 24614 2204 24616
rect 2260 24614 2284 24616
rect 1964 24605 2340 24614
rect 790 23447 842 23453
rect 790 23389 842 23395
rect 802 23199 830 23389
rect 1964 23338 2340 23347
rect 2020 23336 2044 23338
rect 2100 23336 2124 23338
rect 2180 23336 2204 23338
rect 2260 23336 2284 23338
rect 2020 23284 2030 23336
rect 2274 23284 2284 23336
rect 2020 23282 2044 23284
rect 2100 23282 2124 23284
rect 2180 23282 2204 23284
rect 2260 23282 2284 23284
rect 1964 23273 2340 23282
rect 788 23190 844 23199
rect 788 23125 844 23134
rect 1846 22337 1898 22343
rect 1846 22279 1898 22285
rect 886 22115 938 22121
rect 886 22057 938 22063
rect 898 21719 926 22057
rect 884 21710 940 21719
rect 884 21645 940 21654
rect 1858 21603 1886 22279
rect 1964 22006 2340 22015
rect 2020 22004 2044 22006
rect 2100 22004 2124 22006
rect 2180 22004 2204 22006
rect 2260 22004 2284 22006
rect 2020 21952 2030 22004
rect 2274 21952 2284 22004
rect 2020 21950 2044 21952
rect 2100 21950 2124 21952
rect 2180 21950 2204 21952
rect 2260 21950 2284 21952
rect 1964 21941 2340 21950
rect 2434 21751 2462 25609
rect 2710 25593 2762 25599
rect 2710 25535 2762 25541
rect 2518 25001 2570 25007
rect 2518 24943 2570 24949
rect 2422 21745 2474 21751
rect 2422 21687 2474 21693
rect 1846 21597 1898 21603
rect 1846 21539 1898 21545
rect 1858 20567 1886 21539
rect 1964 20674 2340 20683
rect 2020 20672 2044 20674
rect 2100 20672 2124 20674
rect 2180 20672 2204 20674
rect 2260 20672 2284 20674
rect 2020 20620 2030 20672
rect 2274 20620 2284 20672
rect 2020 20618 2044 20620
rect 2100 20618 2124 20620
rect 2180 20618 2204 20620
rect 2260 20618 2284 20620
rect 1964 20609 2340 20618
rect 1846 20561 1898 20567
rect 1846 20503 1898 20509
rect 2434 20419 2462 21687
rect 2422 20413 2474 20419
rect 2422 20355 2474 20361
rect 1556 20230 1612 20239
rect 1556 20165 1612 20174
rect 1570 19901 1598 20165
rect 1558 19895 1610 19901
rect 1558 19837 1610 19843
rect 1750 19673 1802 19679
rect 1750 19615 1802 19621
rect 1762 19235 1790 19615
rect 1964 19342 2340 19351
rect 2020 19340 2044 19342
rect 2100 19340 2124 19342
rect 2180 19340 2204 19342
rect 2260 19340 2284 19342
rect 2020 19288 2030 19340
rect 2274 19288 2284 19340
rect 2020 19286 2044 19288
rect 2100 19286 2124 19288
rect 2180 19286 2204 19288
rect 2260 19286 2284 19288
rect 1964 19277 2340 19286
rect 1750 19229 1802 19235
rect 1750 19171 1802 19177
rect 2434 19087 2462 20355
rect 2422 19081 2474 19087
rect 2422 19023 2474 19029
rect 1556 18750 1612 18759
rect 1556 18685 1612 18694
rect 1570 18569 1598 18685
rect 1558 18563 1610 18569
rect 1558 18505 1610 18511
rect 1750 18341 1802 18347
rect 1750 18283 1802 18289
rect 1762 17903 1790 18283
rect 1964 18010 2340 18019
rect 2020 18008 2044 18010
rect 2100 18008 2124 18010
rect 2180 18008 2204 18010
rect 2260 18008 2284 18010
rect 2020 17956 2030 18008
rect 2274 17956 2284 18008
rect 2020 17954 2044 17956
rect 2100 17954 2124 17956
rect 2180 17954 2204 17956
rect 2260 17954 2284 17956
rect 1964 17945 2340 17954
rect 1750 17897 1802 17903
rect 1750 17839 1802 17845
rect 2434 17755 2462 19023
rect 2422 17749 2474 17755
rect 2422 17691 2474 17697
rect 1268 17270 1324 17279
rect 1268 17205 1270 17214
rect 1322 17205 1324 17214
rect 1270 17173 1322 17179
rect 1750 17009 1802 17015
rect 1750 16951 1802 16957
rect 1762 16571 1790 16951
rect 1964 16678 2340 16687
rect 2020 16676 2044 16678
rect 2100 16676 2124 16678
rect 2180 16676 2204 16678
rect 2260 16676 2284 16678
rect 2020 16624 2030 16676
rect 2274 16624 2284 16676
rect 2020 16622 2044 16624
rect 2100 16622 2124 16624
rect 2180 16622 2204 16624
rect 2260 16622 2284 16624
rect 1964 16613 2340 16622
rect 1750 16565 1802 16571
rect 1750 16507 1802 16513
rect 788 15790 844 15799
rect 788 15725 790 15734
rect 842 15725 844 15734
rect 790 15693 842 15699
rect 1964 15346 2340 15355
rect 2020 15344 2044 15346
rect 2100 15344 2124 15346
rect 2180 15344 2204 15346
rect 2260 15344 2284 15346
rect 2020 15292 2030 15344
rect 2274 15292 2284 15344
rect 2020 15290 2044 15292
rect 2100 15290 2124 15292
rect 2180 15290 2204 15292
rect 2260 15290 2284 15292
rect 1964 15281 2340 15290
rect 788 14310 844 14319
rect 788 14245 790 14254
rect 842 14245 844 14254
rect 790 14213 842 14219
rect 1964 14014 2340 14023
rect 2020 14012 2044 14014
rect 2100 14012 2124 14014
rect 2180 14012 2204 14014
rect 2260 14012 2284 14014
rect 2020 13960 2030 14012
rect 2274 13960 2284 14012
rect 2020 13958 2044 13960
rect 2100 13958 2124 13960
rect 2180 13958 2204 13960
rect 2260 13958 2284 13960
rect 1964 13949 2340 13958
rect 1558 13013 1610 13019
rect 1558 12955 1610 12961
rect 1462 12939 1514 12945
rect 1462 12881 1514 12887
rect 1474 12279 1502 12881
rect 1570 12839 1598 12955
rect 1556 12830 1612 12839
rect 1556 12765 1612 12774
rect 1964 12682 2340 12691
rect 2020 12680 2044 12682
rect 2100 12680 2124 12682
rect 2180 12680 2204 12682
rect 2260 12680 2284 12682
rect 2020 12628 2030 12680
rect 2274 12628 2284 12680
rect 2020 12626 2044 12628
rect 2100 12626 2124 12628
rect 2180 12626 2204 12628
rect 2260 12626 2284 12628
rect 1964 12617 2340 12626
rect 1846 12347 1898 12353
rect 1846 12289 1898 12295
rect 1462 12273 1514 12279
rect 1462 12215 1514 12221
rect 1474 11761 1502 12215
rect 1462 11755 1514 11761
rect 1462 11697 1514 11703
rect 1474 7543 1502 11697
rect 1558 11459 1610 11465
rect 1558 11401 1610 11407
rect 1570 11359 1598 11401
rect 1556 11350 1612 11359
rect 1556 11285 1612 11294
rect 1858 10892 1886 12289
rect 1964 11350 2340 11359
rect 2020 11348 2044 11350
rect 2100 11348 2124 11350
rect 2180 11348 2204 11350
rect 2260 11348 2284 11350
rect 2020 11296 2030 11348
rect 2274 11296 2284 11348
rect 2020 11294 2044 11296
rect 2100 11294 2124 11296
rect 2180 11294 2204 11296
rect 2260 11294 2284 11296
rect 1964 11285 2340 11294
rect 2530 11243 2558 24943
rect 2722 13167 2750 25535
rect 2806 17675 2858 17681
rect 2806 17617 2858 17623
rect 2818 16423 2846 17617
rect 2902 16861 2954 16867
rect 2902 16803 2954 16809
rect 2806 16417 2858 16423
rect 2806 16359 2858 16365
rect 2818 15609 2846 16359
rect 2914 15757 2942 16803
rect 2998 16269 3050 16275
rect 2998 16211 3050 16217
rect 2902 15751 2954 15757
rect 2902 15693 2954 15699
rect 2806 15603 2858 15609
rect 2806 15545 2858 15551
rect 2818 15091 2846 15545
rect 2806 15085 2858 15091
rect 2806 15027 2858 15033
rect 2818 14499 2846 15027
rect 2806 14493 2858 14499
rect 2806 14435 2858 14441
rect 2914 14444 2942 15693
rect 3010 15683 3038 16211
rect 2998 15677 3050 15683
rect 2998 15619 3050 15625
rect 3010 14795 3038 15619
rect 2998 14789 3050 14795
rect 2998 14731 3050 14737
rect 2710 13161 2762 13167
rect 2710 13103 2762 13109
rect 2818 12945 2846 14435
rect 2914 14416 3038 14444
rect 2902 14271 2954 14277
rect 2902 14213 2954 14219
rect 2914 13611 2942 14213
rect 2902 13605 2954 13611
rect 2902 13547 2954 13553
rect 2914 13019 2942 13547
rect 2902 13013 2954 13019
rect 2902 12955 2954 12961
rect 2806 12939 2858 12945
rect 2806 12881 2858 12887
rect 2818 12427 2846 12881
rect 2806 12421 2858 12427
rect 2806 12363 2858 12369
rect 2710 11681 2762 11687
rect 2710 11623 2762 11629
rect 2518 11237 2570 11243
rect 2518 11179 2570 11185
rect 1942 11015 1994 11021
rect 1942 10957 1994 10963
rect 1762 10864 1886 10892
rect 1558 10127 1610 10133
rect 1558 10069 1610 10075
rect 1570 9879 1598 10069
rect 1556 9870 1612 9879
rect 1556 9805 1612 9814
rect 1654 8943 1706 8949
rect 1654 8885 1706 8891
rect 1666 8399 1694 8885
rect 1762 8579 1790 10864
rect 1954 10355 1982 10957
rect 2722 10355 2750 11623
rect 2818 11465 2846 12363
rect 2806 11459 2858 11465
rect 2806 11401 2858 11407
rect 2818 11095 2846 11401
rect 2806 11089 2858 11095
rect 2806 11031 2858 11037
rect 1942 10349 1994 10355
rect 1942 10291 1994 10297
rect 2710 10349 2762 10355
rect 2710 10291 2762 10297
rect 1954 10152 1982 10291
rect 1858 10124 1982 10152
rect 2710 10201 2762 10207
rect 2818 10152 2846 11031
rect 2914 10947 2942 12955
rect 3010 11539 3038 14416
rect 3202 13112 3230 25609
rect 4964 25336 5340 25345
rect 5020 25334 5044 25336
rect 5100 25334 5124 25336
rect 5180 25334 5204 25336
rect 5260 25334 5284 25336
rect 5020 25282 5030 25334
rect 5274 25282 5284 25334
rect 5020 25280 5044 25282
rect 5100 25280 5124 25282
rect 5180 25280 5204 25282
rect 5260 25280 5284 25282
rect 4964 25271 5340 25280
rect 4964 24004 5340 24013
rect 5020 24002 5044 24004
rect 5100 24002 5124 24004
rect 5180 24002 5204 24004
rect 5260 24002 5284 24004
rect 5020 23950 5030 24002
rect 5274 23950 5284 24002
rect 5020 23948 5044 23950
rect 5100 23948 5124 23950
rect 5180 23948 5204 23950
rect 5260 23948 5284 23950
rect 4964 23939 5340 23948
rect 3862 23669 3914 23675
rect 3862 23611 3914 23617
rect 3874 23157 3902 23611
rect 3862 23151 3914 23157
rect 3862 23093 3914 23099
rect 3874 21751 3902 23093
rect 4964 22672 5340 22681
rect 5020 22670 5044 22672
rect 5100 22670 5124 22672
rect 5180 22670 5204 22672
rect 5260 22670 5284 22672
rect 5020 22618 5030 22670
rect 5274 22618 5284 22670
rect 5020 22616 5044 22618
rect 5100 22616 5124 22618
rect 5180 22616 5204 22618
rect 5260 22616 5284 22618
rect 4964 22607 5340 22616
rect 3862 21745 3914 21751
rect 3862 21687 3914 21693
rect 3286 21671 3338 21677
rect 3286 21613 3338 21619
rect 3298 20345 3326 21613
rect 4964 21340 5340 21349
rect 5020 21338 5044 21340
rect 5100 21338 5124 21340
rect 5180 21338 5204 21340
rect 5260 21338 5284 21340
rect 5020 21286 5030 21338
rect 5274 21286 5284 21338
rect 5020 21284 5044 21286
rect 5100 21284 5124 21286
rect 5180 21284 5204 21286
rect 5260 21284 5284 21286
rect 4964 21275 5340 21284
rect 5398 20413 5450 20419
rect 5398 20355 5450 20361
rect 3286 20339 3338 20345
rect 3286 20281 3338 20287
rect 3670 20339 3722 20345
rect 3670 20281 3722 20287
rect 3298 19013 3326 20281
rect 3682 19679 3710 20281
rect 4964 20008 5340 20017
rect 5020 20006 5044 20008
rect 5100 20006 5124 20008
rect 5180 20006 5204 20008
rect 5260 20006 5284 20008
rect 5020 19954 5030 20006
rect 5274 19954 5284 20006
rect 5020 19952 5044 19954
rect 5100 19952 5124 19954
rect 5180 19952 5204 19954
rect 5260 19952 5284 19954
rect 4964 19943 5340 19952
rect 3670 19673 3722 19679
rect 3670 19615 3722 19621
rect 5410 19161 5438 20355
rect 5398 19155 5450 19161
rect 5398 19097 5450 19103
rect 4438 19081 4490 19087
rect 4438 19023 4490 19029
rect 3286 19007 3338 19013
rect 3286 18949 3338 18955
rect 4150 19007 4202 19013
rect 4150 18949 4202 18955
rect 3298 17681 3326 18949
rect 4162 18347 4190 18949
rect 4150 18341 4202 18347
rect 4150 18283 4202 18289
rect 3286 17675 3338 17681
rect 3286 17617 3338 17623
rect 3298 16349 3326 17617
rect 3958 17009 4010 17015
rect 3958 16951 4010 16957
rect 3286 16343 3338 16349
rect 3286 16285 3338 16291
rect 3298 15017 3326 16285
rect 3970 16275 3998 16951
rect 3958 16269 4010 16275
rect 3958 16211 4010 16217
rect 3670 15677 3722 15683
rect 3670 15619 3722 15625
rect 3286 15011 3338 15017
rect 3286 14953 3338 14959
rect 3106 13084 3230 13112
rect 3106 11909 3134 13084
rect 3298 12353 3326 14953
rect 3682 14943 3710 15619
rect 3670 14937 3722 14943
rect 3670 14879 3722 14885
rect 3382 14789 3434 14795
rect 3382 14731 3434 14737
rect 3394 13019 3422 14731
rect 3682 14351 3710 14879
rect 3670 14345 3722 14351
rect 3670 14287 3722 14293
rect 3382 13013 3434 13019
rect 3382 12955 3434 12961
rect 3286 12347 3338 12353
rect 3286 12289 3338 12295
rect 3682 12131 3710 14287
rect 4162 13685 4190 18283
rect 4450 17755 4478 19023
rect 4964 18676 5340 18685
rect 5020 18674 5044 18676
rect 5100 18674 5124 18676
rect 5180 18674 5204 18676
rect 5260 18674 5284 18676
rect 5020 18622 5030 18674
rect 5274 18622 5284 18674
rect 5020 18620 5044 18622
rect 5100 18620 5124 18622
rect 5180 18620 5204 18622
rect 5260 18620 5284 18622
rect 4964 18611 5340 18620
rect 4438 17749 4490 17755
rect 4438 17691 4490 17697
rect 4246 17675 4298 17681
rect 4246 17617 4298 17623
rect 4258 17089 4286 17617
rect 4246 17083 4298 17089
rect 4246 17025 4298 17031
rect 4258 14351 4286 17025
rect 4450 16867 4478 17691
rect 4964 17344 5340 17353
rect 5020 17342 5044 17344
rect 5100 17342 5124 17344
rect 5180 17342 5204 17344
rect 5260 17342 5284 17344
rect 5020 17290 5030 17342
rect 5274 17290 5284 17342
rect 5020 17288 5044 17290
rect 5100 17288 5124 17290
rect 5180 17288 5204 17290
rect 5260 17288 5284 17290
rect 4964 17279 5340 17288
rect 4438 16861 4490 16867
rect 4438 16803 4490 16809
rect 5506 16812 5534 25609
rect 5686 25593 5738 25599
rect 5686 25535 5738 25541
rect 5590 24927 5642 24933
rect 5590 24869 5642 24875
rect 5602 23601 5630 24869
rect 5590 23595 5642 23601
rect 5590 23537 5642 23543
rect 5602 23009 5630 23537
rect 5590 23003 5642 23009
rect 5590 22945 5642 22951
rect 5602 20567 5630 22945
rect 5590 20561 5642 20567
rect 5590 20503 5642 20509
rect 5590 19081 5642 19087
rect 5590 19023 5642 19029
rect 5602 17829 5630 19023
rect 5590 17823 5642 17829
rect 5590 17765 5642 17771
rect 5602 16941 5630 17765
rect 5590 16935 5642 16941
rect 5590 16877 5642 16883
rect 5506 16793 5630 16812
rect 5506 16787 5642 16793
rect 5506 16784 5590 16787
rect 5590 16729 5642 16735
rect 4964 16012 5340 16021
rect 5020 16010 5044 16012
rect 5100 16010 5124 16012
rect 5180 16010 5204 16012
rect 5260 16010 5284 16012
rect 5020 15958 5030 16010
rect 5274 15958 5284 16010
rect 5020 15956 5044 15958
rect 5100 15956 5124 15958
rect 5180 15956 5204 15958
rect 5260 15956 5284 15958
rect 4964 15947 5340 15956
rect 5602 15757 5630 16729
rect 5590 15751 5642 15757
rect 5590 15693 5642 15699
rect 5698 15461 5726 25535
rect 6070 23521 6122 23527
rect 6070 23463 6122 23469
rect 6082 23083 6110 23463
rect 6070 23077 6122 23083
rect 6070 23019 6122 23025
rect 6082 22787 6110 23019
rect 6070 22781 6122 22787
rect 6070 22723 6122 22729
rect 6082 20419 6110 22723
rect 6070 20413 6122 20419
rect 6070 20355 6122 20361
rect 5878 20339 5930 20345
rect 5878 20281 5930 20287
rect 5398 15455 5450 15461
rect 5398 15397 5450 15403
rect 5686 15455 5738 15461
rect 5686 15397 5738 15403
rect 4964 14680 5340 14689
rect 5020 14678 5044 14680
rect 5100 14678 5124 14680
rect 5180 14678 5204 14680
rect 5260 14678 5284 14680
rect 5020 14626 5030 14678
rect 5274 14626 5284 14678
rect 5020 14624 5044 14626
rect 5100 14624 5124 14626
rect 5180 14624 5204 14626
rect 5260 14624 5284 14626
rect 4964 14615 5340 14624
rect 5410 14499 5438 15397
rect 5398 14493 5450 14499
rect 5398 14435 5450 14441
rect 4246 14345 4298 14351
rect 4246 14287 4298 14293
rect 4630 14271 4682 14277
rect 4630 14213 4682 14219
rect 4642 13759 4670 14213
rect 4630 13753 4682 13759
rect 4630 13695 4682 13701
rect 4150 13679 4202 13685
rect 4150 13621 4202 13627
rect 4964 13348 5340 13357
rect 5020 13346 5044 13348
rect 5100 13346 5124 13348
rect 5180 13346 5204 13348
rect 5260 13346 5284 13348
rect 5020 13294 5030 13346
rect 5274 13294 5284 13346
rect 5020 13292 5044 13294
rect 5100 13292 5124 13294
rect 5180 13292 5204 13294
rect 5260 13292 5284 13294
rect 4964 13283 5340 13292
rect 4342 13161 4394 13167
rect 4342 13103 4394 13109
rect 3670 12125 3722 12131
rect 3670 12067 3722 12073
rect 4246 12125 4298 12131
rect 4246 12067 4298 12073
rect 3094 11903 3146 11909
rect 3094 11845 3146 11851
rect 2998 11533 3050 11539
rect 2998 11475 3050 11481
rect 3010 11169 3038 11475
rect 2998 11163 3050 11169
rect 2998 11105 3050 11111
rect 2902 10941 2954 10947
rect 2902 10883 2954 10889
rect 2762 10149 2846 10152
rect 2710 10143 2846 10149
rect 2722 10124 2846 10143
rect 1750 8573 1802 8579
rect 1750 8515 1802 8521
rect 1652 8390 1708 8399
rect 1652 8325 1708 8334
rect 1654 8277 1706 8283
rect 1654 8219 1706 8225
rect 1558 7759 1610 7765
rect 1558 7701 1610 7707
rect 1462 7537 1514 7543
rect 1462 7479 1514 7485
rect 1570 7247 1598 7701
rect 1558 7241 1610 7247
rect 1558 7183 1610 7189
rect 1570 5767 1598 7183
rect 1666 6919 1694 8219
rect 1762 7691 1790 8515
rect 1858 7765 1886 10124
rect 1964 10018 2340 10027
rect 2020 10016 2044 10018
rect 2100 10016 2124 10018
rect 2180 10016 2204 10018
rect 2260 10016 2284 10018
rect 2020 9964 2030 10016
rect 2274 9964 2284 10016
rect 2020 9962 2044 9964
rect 2100 9962 2124 9964
rect 2180 9962 2204 9964
rect 2260 9962 2284 9964
rect 1964 9953 2340 9962
rect 1964 8686 2340 8695
rect 2020 8684 2044 8686
rect 2100 8684 2124 8686
rect 2180 8684 2204 8686
rect 2260 8684 2284 8686
rect 2020 8632 2030 8684
rect 2274 8632 2284 8684
rect 2020 8630 2044 8632
rect 2100 8630 2124 8632
rect 2180 8630 2204 8632
rect 2260 8630 2284 8632
rect 1964 8621 2340 8630
rect 1846 7759 1898 7765
rect 1846 7701 1898 7707
rect 1750 7685 1802 7691
rect 1750 7627 1802 7633
rect 2722 7617 2750 10124
rect 2914 8949 2942 10883
rect 3010 10429 3038 11105
rect 4258 11021 4286 12067
rect 4246 11015 4298 11021
rect 4246 10957 4298 10963
rect 4354 10577 4382 13103
rect 5494 13013 5546 13019
rect 5494 12955 5546 12961
rect 4964 12016 5340 12025
rect 5020 12014 5044 12016
rect 5100 12014 5124 12016
rect 5180 12014 5204 12016
rect 5260 12014 5284 12016
rect 5020 11962 5030 12014
rect 5274 11962 5284 12014
rect 5020 11960 5044 11962
rect 5100 11960 5124 11962
rect 5180 11960 5204 11962
rect 5260 11960 5284 11962
rect 4964 11951 5340 11960
rect 4438 10793 4490 10799
rect 4438 10735 4490 10741
rect 4342 10571 4394 10577
rect 4342 10513 4394 10519
rect 2998 10423 3050 10429
rect 2998 10365 3050 10371
rect 3670 10349 3722 10355
rect 3670 10291 3722 10297
rect 2902 8943 2954 8949
rect 2902 8885 2954 8891
rect 2806 7685 2858 7691
rect 2806 7627 2858 7633
rect 2710 7611 2762 7617
rect 2710 7553 2762 7559
rect 1750 7537 1802 7543
rect 1750 7479 1802 7485
rect 1652 6910 1708 6919
rect 1652 6845 1708 6854
rect 1762 6581 1790 7479
rect 1964 7354 2340 7363
rect 2020 7352 2044 7354
rect 2100 7352 2124 7354
rect 2180 7352 2204 7354
rect 2260 7352 2284 7354
rect 2020 7300 2030 7352
rect 2274 7300 2284 7352
rect 2020 7298 2044 7300
rect 2100 7298 2124 7300
rect 2180 7298 2204 7300
rect 2260 7298 2284 7300
rect 1964 7289 2340 7298
rect 2722 6951 2750 7553
rect 2818 7025 2846 7627
rect 2806 7019 2858 7025
rect 2806 6961 2858 6967
rect 2710 6945 2762 6951
rect 2710 6887 2762 6893
rect 1750 6575 1802 6581
rect 1750 6517 1802 6523
rect 1762 5860 1790 6517
rect 2722 6211 2750 6887
rect 2818 6433 2846 6961
rect 2806 6427 2858 6433
rect 2806 6369 2858 6375
rect 2710 6205 2762 6211
rect 2710 6147 2762 6153
rect 1964 6022 2340 6031
rect 2020 6020 2044 6022
rect 2100 6020 2124 6022
rect 2180 6020 2204 6022
rect 2260 6020 2284 6022
rect 2020 5968 2030 6020
rect 2274 5968 2284 6020
rect 2020 5966 2044 5968
rect 2100 5966 2124 5968
rect 2180 5966 2204 5968
rect 2260 5966 2284 5968
rect 1964 5957 2340 5966
rect 1762 5832 1886 5860
rect 1558 5761 1610 5767
rect 1558 5703 1610 5709
rect 1654 5613 1706 5619
rect 1654 5555 1706 5561
rect 1666 5101 1694 5555
rect 1858 5101 1886 5832
rect 2722 5767 2750 6147
rect 2710 5761 2762 5767
rect 2710 5703 2762 5709
rect 1654 5095 1706 5101
rect 1654 5037 1706 5043
rect 1846 5095 1898 5101
rect 1846 5037 1898 5043
rect 2722 4953 2750 5703
rect 2914 5619 2942 8885
rect 3682 7913 3710 10291
rect 3670 7907 3722 7913
rect 3670 7849 3722 7855
rect 3682 7214 3710 7849
rect 3682 7186 3806 7214
rect 3778 6285 3806 7186
rect 3766 6279 3818 6285
rect 3766 6221 3818 6227
rect 2902 5613 2954 5619
rect 2954 5561 3038 5564
rect 2902 5555 3038 5561
rect 2914 5536 3038 5555
rect 2902 5465 2954 5471
rect 2902 5407 2954 5413
rect 2710 4947 2762 4953
rect 2710 4889 2762 4895
rect 1964 4690 2340 4699
rect 2020 4688 2044 4690
rect 2100 4688 2124 4690
rect 2180 4688 2204 4690
rect 2260 4688 2284 4690
rect 2020 4636 2030 4688
rect 2274 4636 2284 4688
rect 2020 4634 2044 4636
rect 2100 4634 2124 4636
rect 2180 4634 2204 4636
rect 2260 4634 2284 4636
rect 1964 4625 2340 4634
rect 2722 4435 2750 4889
rect 2710 4429 2762 4435
rect 2710 4371 2762 4377
rect 1654 4133 1706 4139
rect 1654 4075 1706 4081
rect 884 3950 940 3959
rect 884 3885 940 3894
rect 898 3695 926 3885
rect 886 3689 938 3695
rect 886 3631 938 3637
rect 598 3097 650 3103
rect 598 3039 650 3045
rect 610 800 638 3039
rect 1666 3029 1694 4075
rect 1964 3358 2340 3367
rect 2020 3356 2044 3358
rect 2100 3356 2124 3358
rect 2180 3356 2204 3358
rect 2260 3356 2284 3358
rect 2020 3304 2030 3356
rect 2274 3304 2284 3356
rect 2020 3302 2044 3304
rect 2100 3302 2124 3304
rect 2180 3302 2204 3304
rect 2260 3302 2284 3304
rect 1964 3293 2340 3302
rect 2914 3029 2942 5407
rect 3010 4287 3038 5536
rect 3286 4799 3338 4805
rect 3286 4741 3338 4747
rect 2998 4281 3050 4287
rect 2998 4223 3050 4229
rect 3298 3029 3326 4741
rect 3778 4361 3806 6221
rect 3766 4355 3818 4361
rect 3766 4297 3818 4303
rect 4450 3029 4478 10735
rect 4964 10684 5340 10693
rect 5020 10682 5044 10684
rect 5100 10682 5124 10684
rect 5180 10682 5204 10684
rect 5260 10682 5284 10684
rect 5020 10630 5030 10682
rect 5274 10630 5284 10682
rect 5020 10628 5044 10630
rect 5100 10628 5124 10630
rect 5180 10628 5204 10630
rect 5260 10628 5284 10630
rect 4964 10619 5340 10628
rect 4964 9352 5340 9361
rect 5020 9350 5044 9352
rect 5100 9350 5124 9352
rect 5180 9350 5204 9352
rect 5260 9350 5284 9352
rect 5020 9298 5030 9350
rect 5274 9298 5284 9350
rect 5020 9296 5044 9298
rect 5100 9296 5124 9298
rect 5180 9296 5204 9298
rect 5260 9296 5284 9298
rect 4964 9287 5340 9296
rect 4964 8020 5340 8029
rect 5020 8018 5044 8020
rect 5100 8018 5124 8020
rect 5180 8018 5204 8020
rect 5260 8018 5284 8020
rect 5020 7966 5030 8018
rect 5274 7966 5284 8018
rect 5020 7964 5044 7966
rect 5100 7964 5124 7966
rect 5180 7964 5204 7966
rect 5260 7964 5284 7966
rect 4964 7955 5340 7964
rect 4964 6688 5340 6697
rect 5020 6686 5044 6688
rect 5100 6686 5124 6688
rect 5180 6686 5204 6688
rect 5260 6686 5284 6688
rect 5020 6634 5030 6686
rect 5274 6634 5284 6686
rect 5020 6632 5044 6634
rect 5100 6632 5124 6634
rect 5180 6632 5204 6634
rect 5260 6632 5284 6634
rect 4964 6623 5340 6632
rect 4822 5613 4874 5619
rect 5110 5613 5162 5619
rect 4874 5561 5110 5564
rect 4822 5555 5162 5561
rect 4834 5536 5150 5555
rect 4630 4799 4682 4805
rect 4630 4741 4682 4747
rect 4642 4361 4670 4741
rect 4630 4355 4682 4361
rect 4630 4297 4682 4303
rect 4642 3103 4670 4297
rect 4834 3843 4862 5536
rect 4964 5356 5340 5365
rect 5020 5354 5044 5356
rect 5100 5354 5124 5356
rect 5180 5354 5204 5356
rect 5260 5354 5284 5356
rect 5020 5302 5030 5354
rect 5274 5302 5284 5354
rect 5020 5300 5044 5302
rect 5100 5300 5124 5302
rect 5180 5300 5204 5302
rect 5260 5300 5284 5302
rect 4964 5291 5340 5300
rect 4964 4024 5340 4033
rect 5020 4022 5044 4024
rect 5100 4022 5124 4024
rect 5180 4022 5204 4024
rect 5260 4022 5284 4024
rect 5020 3970 5030 4022
rect 5274 3970 5284 4022
rect 5020 3968 5044 3970
rect 5100 3968 5124 3970
rect 5180 3968 5204 3970
rect 5260 3968 5284 3970
rect 4964 3959 5340 3968
rect 4822 3837 4874 3843
rect 4822 3779 4874 3785
rect 4630 3097 4682 3103
rect 4630 3039 4682 3045
rect 5506 3029 5534 12955
rect 5890 11687 5918 20281
rect 6082 19161 6110 20355
rect 6070 19155 6122 19161
rect 6070 19097 6122 19103
rect 6466 18421 6494 25609
rect 7606 25593 7658 25599
rect 7606 25535 7658 25541
rect 6742 23669 6794 23675
rect 6742 23611 6794 23617
rect 6754 23157 6782 23611
rect 6742 23151 6794 23157
rect 6742 23093 6794 23099
rect 6550 22929 6602 22935
rect 6550 22871 6602 22877
rect 6562 22343 6590 22871
rect 6550 22337 6602 22343
rect 6550 22279 6602 22285
rect 6454 18415 6506 18421
rect 6454 18357 6506 18363
rect 6466 17903 6494 18357
rect 6454 17897 6506 17903
rect 6454 17839 6506 17845
rect 6166 13605 6218 13611
rect 6166 13547 6218 13553
rect 6178 12427 6206 13547
rect 6166 12421 6218 12427
rect 6166 12363 6218 12369
rect 5878 11681 5930 11687
rect 5878 11623 5930 11629
rect 6178 11613 6206 12363
rect 6562 12353 6590 22279
rect 6550 12347 6602 12353
rect 6550 12289 6602 12295
rect 6166 11607 6218 11613
rect 6166 11549 6218 11555
rect 6178 11095 6206 11549
rect 6166 11089 6218 11095
rect 6166 11031 6218 11037
rect 6754 11021 6782 23093
rect 7618 23009 7646 25535
rect 7606 23003 7658 23009
rect 7606 22945 7658 22951
rect 7618 21085 7646 22945
rect 7606 21079 7658 21085
rect 7606 21021 7658 21027
rect 7810 18791 7838 25609
rect 7906 20567 7934 25609
rect 8470 25001 8522 25007
rect 8470 24943 8522 24949
rect 7964 24670 8340 24679
rect 8020 24668 8044 24670
rect 8100 24668 8124 24670
rect 8180 24668 8204 24670
rect 8260 24668 8284 24670
rect 8020 24616 8030 24668
rect 8274 24616 8284 24668
rect 8020 24614 8044 24616
rect 8100 24614 8124 24616
rect 8180 24614 8204 24616
rect 8260 24614 8284 24616
rect 7964 24605 8340 24614
rect 8482 23897 8510 24943
rect 9442 23897 9470 25609
rect 10978 25229 11006 28074
rect 10966 25223 11018 25229
rect 10966 25165 11018 25171
rect 8470 23891 8522 23897
rect 8470 23833 8522 23839
rect 9430 23891 9482 23897
rect 9430 23833 9482 23839
rect 7964 23338 8340 23347
rect 8020 23336 8044 23338
rect 8100 23336 8124 23338
rect 8180 23336 8204 23338
rect 8260 23336 8284 23338
rect 8020 23284 8030 23336
rect 8274 23284 8284 23336
rect 8020 23282 8044 23284
rect 8100 23282 8124 23284
rect 8180 23282 8204 23284
rect 8260 23282 8284 23284
rect 7964 23273 8340 23282
rect 8374 22929 8426 22935
rect 8374 22871 8426 22877
rect 8386 22343 8414 22871
rect 8482 22417 8510 23833
rect 8758 23669 8810 23675
rect 8758 23611 8810 23617
rect 8770 22861 8798 23611
rect 9814 23003 9866 23009
rect 9814 22945 9866 22951
rect 8758 22855 8810 22861
rect 8758 22797 8810 22803
rect 9826 22565 9854 22945
rect 10102 22781 10154 22787
rect 10102 22723 10154 22729
rect 10114 22607 10142 22723
rect 10100 22598 10156 22607
rect 9814 22559 9866 22565
rect 10100 22533 10156 22542
rect 9814 22501 9866 22507
rect 8470 22411 8522 22417
rect 8470 22353 8522 22359
rect 8374 22337 8426 22343
rect 8374 22279 8426 22285
rect 7964 22006 8340 22015
rect 8020 22004 8044 22006
rect 8100 22004 8124 22006
rect 8180 22004 8204 22006
rect 8260 22004 8284 22006
rect 8020 21952 8030 22004
rect 8274 21952 8284 22004
rect 8020 21950 8044 21952
rect 8100 21950 8124 21952
rect 8180 21950 8204 21952
rect 8260 21950 8284 21952
rect 7964 21941 8340 21950
rect 8386 21677 8414 22279
rect 8662 22263 8714 22269
rect 8662 22205 8714 22211
rect 8374 21671 8426 21677
rect 8374 21613 8426 21619
rect 8386 21011 8414 21613
rect 8374 21005 8426 21011
rect 8374 20947 8426 20953
rect 7964 20674 8340 20683
rect 8020 20672 8044 20674
rect 8100 20672 8124 20674
rect 8180 20672 8204 20674
rect 8260 20672 8284 20674
rect 8020 20620 8030 20672
rect 8274 20620 8284 20672
rect 8020 20618 8044 20620
rect 8100 20618 8124 20620
rect 8180 20618 8204 20620
rect 8260 20618 8284 20620
rect 7964 20609 8340 20618
rect 7894 20561 7946 20567
rect 7894 20503 7946 20509
rect 7906 19753 7934 20503
rect 7894 19747 7946 19753
rect 7894 19689 7946 19695
rect 8386 19679 8414 20947
rect 8674 20937 8702 22205
rect 8662 20931 8714 20937
rect 8662 20873 8714 20879
rect 8374 19673 8426 19679
rect 8374 19615 8426 19621
rect 8674 19605 8702 20873
rect 9814 20783 9866 20789
rect 9814 20725 9866 20731
rect 9826 20345 9854 20725
rect 9814 20339 9866 20345
rect 9814 20281 9866 20287
rect 10100 20230 10156 20239
rect 10100 20165 10102 20174
rect 10154 20165 10156 20174
rect 10102 20133 10154 20139
rect 7894 19599 7946 19605
rect 7894 19541 7946 19547
rect 8662 19599 8714 19605
rect 8662 19541 8714 19547
rect 7798 18785 7850 18791
rect 7798 18727 7850 18733
rect 7810 17089 7838 18727
rect 7906 18347 7934 19541
rect 7964 19342 8340 19351
rect 8020 19340 8044 19342
rect 8100 19340 8124 19342
rect 8180 19340 8204 19342
rect 8260 19340 8284 19342
rect 8020 19288 8030 19340
rect 8274 19288 8284 19340
rect 8020 19286 8044 19288
rect 8100 19286 8124 19288
rect 8180 19286 8204 19288
rect 8260 19286 8284 19288
rect 7964 19277 8340 19286
rect 7894 18341 7946 18347
rect 7894 18283 7946 18289
rect 7798 17083 7850 17089
rect 7798 17025 7850 17031
rect 7906 17015 7934 18283
rect 8674 18273 8702 19541
rect 9814 19451 9866 19457
rect 9814 19393 9866 19399
rect 8662 18267 8714 18273
rect 8662 18209 8714 18215
rect 7964 18010 8340 18019
rect 8020 18008 8044 18010
rect 8100 18008 8124 18010
rect 8180 18008 8204 18010
rect 8260 18008 8284 18010
rect 8020 17956 8030 18008
rect 8274 17956 8284 18008
rect 8020 17954 8044 17956
rect 8100 17954 8124 17956
rect 8180 17954 8204 17956
rect 8260 17954 8284 17956
rect 7964 17945 8340 17954
rect 8674 17294 8702 18209
rect 9718 18119 9770 18125
rect 9718 18061 9770 18067
rect 8674 17266 8798 17294
rect 7894 17009 7946 17015
rect 7894 16951 7946 16957
rect 7906 15683 7934 16951
rect 8770 16941 8798 17266
rect 8758 16935 8810 16941
rect 8758 16877 8810 16883
rect 7964 16678 8340 16687
rect 8020 16676 8044 16678
rect 8100 16676 8124 16678
rect 8180 16676 8204 16678
rect 8260 16676 8284 16678
rect 8020 16624 8030 16676
rect 8274 16624 8284 16676
rect 8020 16622 8044 16624
rect 8100 16622 8124 16624
rect 8180 16622 8204 16624
rect 8260 16622 8284 16624
rect 7964 16613 8340 16622
rect 7894 15677 7946 15683
rect 7894 15619 7946 15625
rect 7906 14351 7934 15619
rect 8770 15609 8798 16877
rect 8758 15603 8810 15609
rect 8758 15545 8810 15551
rect 7964 15346 8340 15355
rect 8020 15344 8044 15346
rect 8100 15344 8124 15346
rect 8180 15344 8204 15346
rect 8260 15344 8284 15346
rect 8020 15292 8030 15344
rect 8274 15292 8284 15344
rect 8020 15290 8044 15292
rect 8100 15290 8124 15292
rect 8180 15290 8204 15292
rect 8260 15290 8284 15292
rect 7964 15281 8340 15290
rect 7894 14345 7946 14351
rect 7894 14287 7946 14293
rect 8374 14345 8426 14351
rect 8374 14287 8426 14293
rect 7030 14123 7082 14129
rect 7030 14065 7082 14071
rect 6742 11015 6794 11021
rect 6742 10957 6794 10963
rect 6262 8425 6314 8431
rect 6262 8367 6314 8373
rect 6274 7025 6302 8367
rect 6358 7907 6410 7913
rect 6358 7849 6410 7855
rect 6262 7019 6314 7025
rect 6262 6961 6314 6967
rect 6370 6581 6398 7849
rect 6838 7463 6890 7469
rect 6838 7405 6890 7411
rect 6850 7099 6878 7405
rect 6838 7093 6890 7099
rect 6838 7035 6890 7041
rect 6454 7019 6506 7025
rect 6454 6961 6506 6967
rect 5878 6575 5930 6581
rect 5878 6517 5930 6523
rect 6358 6575 6410 6581
rect 6358 6517 6410 6523
rect 5686 6353 5738 6359
rect 5686 6295 5738 6301
rect 5698 6211 5726 6295
rect 5686 6205 5738 6211
rect 5686 6147 5738 6153
rect 5698 5619 5726 6147
rect 5686 5613 5738 5619
rect 5686 5555 5738 5561
rect 5698 5249 5726 5555
rect 5686 5243 5738 5249
rect 5686 5185 5738 5191
rect 5782 4947 5834 4953
rect 5782 4889 5834 4895
rect 5794 4583 5822 4889
rect 5782 4577 5834 4583
rect 5782 4519 5834 4525
rect 5890 3917 5918 6517
rect 6070 6501 6122 6507
rect 6070 6443 6122 6449
rect 5974 6427 6026 6433
rect 5974 6369 6026 6375
rect 5986 5471 6014 6369
rect 6082 5712 6110 6443
rect 6466 6359 6494 6961
rect 6454 6353 6506 6359
rect 6454 6295 6506 6301
rect 6082 5693 6206 5712
rect 6070 5687 6206 5693
rect 6122 5684 6206 5687
rect 6070 5629 6122 5635
rect 6070 5539 6122 5545
rect 6070 5481 6122 5487
rect 5974 5465 6026 5471
rect 5974 5407 6026 5413
rect 5986 4361 6014 5407
rect 6082 4435 6110 5481
rect 6070 4429 6122 4435
rect 6070 4371 6122 4377
rect 5974 4355 6026 4361
rect 5974 4297 6026 4303
rect 5878 3911 5930 3917
rect 5878 3853 5930 3859
rect 6178 3769 6206 5684
rect 6358 5687 6410 5693
rect 6358 5629 6410 5635
rect 6370 5587 6398 5629
rect 6356 5578 6412 5587
rect 6356 5513 6412 5522
rect 6466 5027 6494 6295
rect 6838 6131 6890 6137
rect 6838 6073 6890 6079
rect 6850 5101 6878 6073
rect 6838 5095 6890 5101
rect 6838 5037 6890 5043
rect 6454 5021 6506 5027
rect 6454 4963 6506 4969
rect 6550 4947 6602 4953
rect 6550 4889 6602 4895
rect 6562 4361 6590 4889
rect 6550 4355 6602 4361
rect 6550 4297 6602 4303
rect 6358 4133 6410 4139
rect 6358 4075 6410 4081
rect 6370 3769 6398 4075
rect 6166 3763 6218 3769
rect 6166 3705 6218 3711
rect 6358 3763 6410 3769
rect 6358 3705 6410 3711
rect 6562 3695 6590 4297
rect 6550 3689 6602 3695
rect 6550 3631 6602 3637
rect 6562 3103 6590 3631
rect 6550 3097 6602 3103
rect 6550 3039 6602 3045
rect 7042 3029 7070 14065
rect 7964 14014 8340 14023
rect 8020 14012 8044 14014
rect 8100 14012 8124 14014
rect 8180 14012 8204 14014
rect 8260 14012 8284 14014
rect 8020 13960 8030 14012
rect 8274 13960 8284 14012
rect 8020 13958 8044 13960
rect 8100 13958 8124 13960
rect 8180 13958 8204 13960
rect 8260 13958 8284 13960
rect 7964 13949 8340 13958
rect 7222 13827 7274 13833
rect 7222 13769 7274 13775
rect 7234 12427 7262 13769
rect 7510 13457 7562 13463
rect 7510 13399 7562 13405
rect 7222 12421 7274 12427
rect 7222 12363 7274 12369
rect 7234 11613 7262 12363
rect 7222 11607 7274 11613
rect 7222 11549 7274 11555
rect 7234 11095 7262 11549
rect 7222 11089 7274 11095
rect 7222 11031 7274 11037
rect 7126 4355 7178 4361
rect 7126 4297 7178 4303
rect 7138 3029 7166 4297
rect 7522 3695 7550 13399
rect 8386 13019 8414 14287
rect 8770 14277 8798 15545
rect 8758 14271 8810 14277
rect 8758 14213 8810 14219
rect 8374 13013 8426 13019
rect 8374 12955 8426 12961
rect 7964 12682 8340 12691
rect 8020 12680 8044 12682
rect 8100 12680 8124 12682
rect 8180 12680 8204 12682
rect 8260 12680 8284 12682
rect 8020 12628 8030 12680
rect 8274 12628 8284 12680
rect 8020 12626 8044 12628
rect 8100 12626 8124 12628
rect 8180 12626 8204 12628
rect 8260 12626 8284 12628
rect 7964 12617 8340 12626
rect 7702 11903 7754 11909
rect 7702 11845 7754 11851
rect 7714 10429 7742 11845
rect 7964 11350 8340 11359
rect 8020 11348 8044 11350
rect 8100 11348 8124 11350
rect 8180 11348 8204 11350
rect 8260 11348 8284 11350
rect 8020 11296 8030 11348
rect 8274 11296 8284 11348
rect 8020 11294 8044 11296
rect 8100 11294 8124 11296
rect 8180 11294 8204 11296
rect 8260 11294 8284 11296
rect 7964 11285 8340 11294
rect 7798 11237 7850 11243
rect 7798 11179 7850 11185
rect 7702 10423 7754 10429
rect 7702 10365 7754 10371
rect 7810 9097 7838 11179
rect 8386 10355 8414 12955
rect 8770 12945 8798 14213
rect 9526 14123 9578 14129
rect 9526 14065 9578 14071
rect 8758 12939 8810 12945
rect 8758 12881 8810 12887
rect 8470 11607 8522 11613
rect 8470 11549 8522 11555
rect 8374 10349 8426 10355
rect 8374 10291 8426 10297
rect 7964 10018 8340 10027
rect 8020 10016 8044 10018
rect 8100 10016 8124 10018
rect 8180 10016 8204 10018
rect 8260 10016 8284 10018
rect 8020 9964 8030 10016
rect 8274 9964 8284 10016
rect 8020 9962 8044 9964
rect 8100 9962 8124 9964
rect 8180 9962 8204 9964
rect 8260 9962 8284 9964
rect 7964 9953 8340 9962
rect 7798 9091 7850 9097
rect 7798 9033 7850 9039
rect 8386 9023 8414 10291
rect 8374 9017 8426 9023
rect 8374 8959 8426 8965
rect 7964 8686 8340 8695
rect 8020 8684 8044 8686
rect 8100 8684 8124 8686
rect 8180 8684 8204 8686
rect 8260 8684 8284 8686
rect 8020 8632 8030 8684
rect 8274 8632 8284 8684
rect 8020 8630 8044 8632
rect 8100 8630 8124 8632
rect 8180 8630 8204 8632
rect 8260 8630 8284 8632
rect 7964 8621 8340 8630
rect 7702 8351 7754 8357
rect 7702 8293 7754 8299
rect 7714 5767 7742 8293
rect 8374 7759 8426 7765
rect 8374 7701 8426 7707
rect 7964 7354 8340 7363
rect 8020 7352 8044 7354
rect 8100 7352 8124 7354
rect 8180 7352 8204 7354
rect 8260 7352 8284 7354
rect 8020 7300 8030 7352
rect 8274 7300 8284 7352
rect 8020 7298 8044 7300
rect 8100 7298 8124 7300
rect 8180 7298 8204 7300
rect 8260 7298 8284 7300
rect 7964 7289 8340 7298
rect 8386 7247 8414 7701
rect 8374 7241 8426 7247
rect 8374 7183 8426 7189
rect 8482 6452 8510 11549
rect 8770 10281 8798 12881
rect 9430 10793 9482 10799
rect 9430 10735 9482 10741
rect 8758 10275 8810 10281
rect 8758 10217 8810 10223
rect 8770 8949 8798 10217
rect 8758 8943 8810 8949
rect 8758 8885 8810 8891
rect 7906 6424 8510 6452
rect 7798 6353 7850 6359
rect 7798 6295 7850 6301
rect 7702 5761 7754 5767
rect 7702 5703 7754 5709
rect 7714 4361 7742 5703
rect 7810 5027 7838 6295
rect 7798 5021 7850 5027
rect 7798 4963 7850 4969
rect 7702 4355 7754 4361
rect 7702 4297 7754 4303
rect 7810 4213 7838 4963
rect 7798 4207 7850 4213
rect 7798 4149 7850 4155
rect 7510 3689 7562 3695
rect 7510 3631 7562 3637
rect 7510 3541 7562 3547
rect 7510 3483 7562 3489
rect 1654 3023 1706 3029
rect 1654 2965 1706 2971
rect 2902 3023 2954 3029
rect 2902 2965 2954 2971
rect 3286 3023 3338 3029
rect 3286 2965 3338 2971
rect 4438 3023 4490 3029
rect 4438 2965 4490 2971
rect 5494 3023 5546 3029
rect 5494 2965 5546 2971
rect 7030 3023 7082 3029
rect 7030 2965 7082 2971
rect 7126 3023 7178 3029
rect 7126 2965 7178 2971
rect 1846 2949 1898 2955
rect 1846 2891 1898 2897
rect 2998 2949 3050 2955
rect 2998 2891 3050 2897
rect 4150 2949 4202 2955
rect 4150 2891 4202 2897
rect 5398 2949 5450 2955
rect 5398 2891 5450 2897
rect 6454 2949 6506 2955
rect 6454 2891 6506 2897
rect 596 0 652 800
rect 1748 680 1804 800
rect 1858 680 1886 2891
rect 2230 2801 2282 2807
rect 2230 2743 2282 2749
rect 2242 2479 2270 2743
rect 2228 2470 2284 2479
rect 2228 2405 2284 2414
rect 1748 652 1886 680
rect 2900 680 2956 800
rect 3010 680 3038 2891
rect 2900 652 3038 680
rect 4052 680 4108 800
rect 4162 680 4190 2891
rect 4964 2692 5340 2701
rect 5020 2690 5044 2692
rect 5100 2690 5124 2692
rect 5180 2690 5204 2692
rect 5260 2690 5284 2692
rect 5020 2638 5030 2690
rect 5274 2638 5284 2690
rect 5020 2636 5044 2638
rect 5100 2636 5124 2638
rect 5180 2636 5204 2638
rect 5260 2636 5284 2638
rect 4964 2627 5340 2636
rect 4052 652 4190 680
rect 5204 680 5260 800
rect 5410 680 5438 2891
rect 5204 652 5438 680
rect 6356 680 6412 800
rect 6466 680 6494 2891
rect 7522 800 7550 3483
rect 7906 3251 7934 6424
rect 8278 6353 8330 6359
rect 8278 6295 8330 6301
rect 8470 6353 8522 6359
rect 8470 6295 8522 6301
rect 8290 6211 8318 6295
rect 8278 6205 8330 6211
rect 8278 6147 8330 6153
rect 8374 6131 8426 6137
rect 8374 6073 8426 6079
rect 7964 6022 8340 6031
rect 8020 6020 8044 6022
rect 8100 6020 8124 6022
rect 8180 6020 8204 6022
rect 8260 6020 8284 6022
rect 8020 5968 8030 6020
rect 8274 5968 8284 6020
rect 8020 5966 8044 5968
rect 8100 5966 8124 5968
rect 8180 5966 8204 5968
rect 8260 5966 8284 5968
rect 7964 5957 8340 5966
rect 8386 5767 8414 6073
rect 8374 5761 8426 5767
rect 8374 5703 8426 5709
rect 8482 5564 8510 6295
rect 8566 6131 8618 6137
rect 8566 6073 8618 6079
rect 8386 5536 8510 5564
rect 8386 5471 8414 5536
rect 8374 5465 8426 5471
rect 8374 5407 8426 5413
rect 8386 5101 8414 5407
rect 8374 5095 8426 5101
rect 8374 5037 8426 5043
rect 7964 4690 8340 4699
rect 8020 4688 8044 4690
rect 8100 4688 8124 4690
rect 8180 4688 8204 4690
rect 8260 4688 8284 4690
rect 8020 4636 8030 4688
rect 8274 4636 8284 4688
rect 8020 4634 8044 4636
rect 8100 4634 8124 4636
rect 8180 4634 8204 4636
rect 8260 4634 8284 4636
rect 7964 4625 8340 4634
rect 8386 4583 8414 5037
rect 8470 4799 8522 4805
rect 8470 4741 8522 4747
rect 8374 4577 8426 4583
rect 8374 4519 8426 4525
rect 8482 4287 8510 4741
rect 8578 4435 8606 6073
rect 8566 4429 8618 4435
rect 8566 4371 8618 4377
rect 8470 4281 8522 4287
rect 8470 4223 8522 4229
rect 8086 4207 8138 4213
rect 8086 4149 8138 4155
rect 8098 3917 8126 4149
rect 8770 4139 8798 8885
rect 8854 6945 8906 6951
rect 8854 6887 8906 6893
rect 8866 6433 8894 6887
rect 8854 6427 8906 6433
rect 8854 6369 8906 6375
rect 9046 6353 9098 6359
rect 9046 6295 9098 6301
rect 9334 6353 9386 6359
rect 9334 6295 9386 6301
rect 9058 5693 9086 6295
rect 9046 5687 9098 5693
rect 9046 5629 9098 5635
rect 9058 5249 9086 5629
rect 9142 5613 9194 5619
rect 9142 5555 9194 5561
rect 9046 5243 9098 5249
rect 9046 5185 9098 5191
rect 9154 5101 9182 5555
rect 9142 5095 9194 5101
rect 9142 5037 9194 5043
rect 9346 4213 9374 6295
rect 9334 4207 9386 4213
rect 9334 4149 9386 4155
rect 8758 4133 8810 4139
rect 8758 4075 8810 4081
rect 8086 3911 8138 3917
rect 8086 3853 8138 3859
rect 8770 3843 8798 4075
rect 8758 3837 8810 3843
rect 8758 3779 8810 3785
rect 9442 3695 9470 10735
rect 9538 8357 9566 14065
rect 9730 13685 9758 18061
rect 9826 17681 9854 19393
rect 10100 17862 10156 17871
rect 10100 17797 10102 17806
rect 10154 17797 10156 17806
rect 10102 17765 10154 17771
rect 9814 17675 9866 17681
rect 9814 17617 9866 17623
rect 9814 16787 9866 16793
rect 9814 16729 9866 16735
rect 9826 15683 9854 16729
rect 9814 15677 9866 15683
rect 9814 15619 9866 15625
rect 10100 15494 10156 15503
rect 9814 15455 9866 15461
rect 10100 15429 10102 15438
rect 9814 15397 9866 15403
rect 10154 15429 10156 15438
rect 10102 15397 10154 15403
rect 9718 13679 9770 13685
rect 9718 13621 9770 13627
rect 9718 12791 9770 12797
rect 9718 12733 9770 12739
rect 9526 8351 9578 8357
rect 9526 8293 9578 8299
rect 9526 7019 9578 7025
rect 9526 6961 9578 6967
rect 9538 5767 9566 6961
rect 9526 5761 9578 5767
rect 9526 5703 9578 5709
rect 9622 5687 9674 5693
rect 9622 5629 9674 5635
rect 9634 5249 9662 5629
rect 9622 5243 9674 5249
rect 9622 5185 9674 5191
rect 9730 3695 9758 12733
rect 9826 11021 9854 15397
rect 10102 13457 10154 13463
rect 10102 13399 10154 13405
rect 10114 13135 10142 13399
rect 10100 13126 10156 13135
rect 10100 13061 10156 13070
rect 10198 12125 10250 12131
rect 10198 12067 10250 12073
rect 9814 11015 9866 11021
rect 9814 10957 9866 10963
rect 10102 10793 10154 10799
rect 10100 10758 10102 10767
rect 10154 10758 10156 10767
rect 10100 10693 10156 10702
rect 9814 10127 9866 10133
rect 9814 10069 9866 10075
rect 9826 6359 9854 10069
rect 10006 8795 10058 8801
rect 10006 8737 10058 8743
rect 9814 6353 9866 6359
rect 9814 6295 9866 6301
rect 9430 3689 9482 3695
rect 9430 3631 9482 3637
rect 9718 3689 9770 3695
rect 9718 3631 9770 3637
rect 7964 3358 8340 3367
rect 8020 3356 8044 3358
rect 8100 3356 8124 3358
rect 8180 3356 8204 3358
rect 8260 3356 8284 3358
rect 8020 3304 8030 3356
rect 8274 3304 8284 3356
rect 8020 3302 8044 3304
rect 8100 3302 8124 3304
rect 8180 3302 8204 3304
rect 8260 3302 8284 3304
rect 7964 3293 8340 3302
rect 7894 3245 7946 3251
rect 7894 3187 7946 3193
rect 10018 3029 10046 8737
rect 10100 8390 10156 8399
rect 10100 8325 10102 8334
rect 10154 8325 10156 8334
rect 10102 8293 10154 8299
rect 10102 6131 10154 6137
rect 10102 6073 10154 6079
rect 10114 6031 10142 6073
rect 10100 6022 10156 6031
rect 10100 5957 10156 5966
rect 10100 3654 10156 3663
rect 10100 3589 10102 3598
rect 10154 3589 10156 3598
rect 10102 3557 10154 3563
rect 10210 3029 10238 12067
rect 10966 3467 11018 3473
rect 10966 3409 11018 3415
rect 10006 3023 10058 3029
rect 10006 2965 10058 2971
rect 10198 3023 10250 3029
rect 10198 2965 10250 2971
rect 8854 2949 8906 2955
rect 8854 2891 8906 2897
rect 9718 2949 9770 2955
rect 9718 2891 9770 2897
rect 9814 2949 9866 2955
rect 9814 2891 9866 2897
rect 6356 652 6494 680
rect 1748 0 1804 652
rect 2900 0 2956 652
rect 4052 0 4108 652
rect 5204 0 5260 652
rect 6356 0 6412 652
rect 7508 0 7564 800
rect 8660 680 8716 800
rect 8866 680 8894 2891
rect 9730 1295 9758 2891
rect 9716 1286 9772 1295
rect 9716 1221 9772 1230
rect 9826 800 9854 2891
rect 10978 800 11006 3409
rect 8660 652 8894 680
rect 8660 0 8716 652
rect 9812 0 9868 800
rect 10964 0 11020 800
<< via2 >>
rect 1652 26094 1708 26150
rect 1964 26000 2020 26002
rect 2044 26000 2100 26002
rect 2124 26000 2180 26002
rect 2204 26000 2260 26002
rect 2284 26000 2340 26002
rect 1964 25948 1966 26000
rect 1966 25948 2018 26000
rect 2018 25948 2020 26000
rect 2044 25948 2082 26000
rect 2082 25948 2094 26000
rect 2094 25948 2100 26000
rect 2124 25948 2146 26000
rect 2146 25948 2158 26000
rect 2158 25948 2180 26000
rect 2204 25948 2210 26000
rect 2210 25948 2222 26000
rect 2222 25948 2260 26000
rect 2284 25948 2286 26000
rect 2286 25948 2338 26000
rect 2338 25948 2340 26000
rect 1964 25946 2020 25948
rect 2044 25946 2100 25948
rect 2124 25946 2180 25948
rect 2204 25946 2260 25948
rect 2284 25946 2340 25948
rect 7964 26000 8020 26002
rect 8044 26000 8100 26002
rect 8124 26000 8180 26002
rect 8204 26000 8260 26002
rect 8284 26000 8340 26002
rect 7964 25948 7966 26000
rect 7966 25948 8018 26000
rect 8018 25948 8020 26000
rect 8044 25948 8082 26000
rect 8082 25948 8094 26000
rect 8094 25948 8100 26000
rect 8124 25948 8146 26000
rect 8146 25948 8158 26000
rect 8158 25948 8180 26000
rect 8204 25948 8210 26000
rect 8210 25948 8222 26000
rect 8222 25948 8260 26000
rect 8284 25948 8286 26000
rect 8286 25948 8338 26000
rect 8338 25948 8340 26000
rect 7964 25946 8020 25948
rect 8044 25946 8100 25948
rect 8124 25946 8180 25948
rect 8204 25946 8260 25948
rect 8284 25946 8340 25948
rect 9716 27278 9772 27334
rect 884 24614 940 24670
rect 1964 24668 2020 24670
rect 2044 24668 2100 24670
rect 2124 24668 2180 24670
rect 2204 24668 2260 24670
rect 2284 24668 2340 24670
rect 1964 24616 1966 24668
rect 1966 24616 2018 24668
rect 2018 24616 2020 24668
rect 2044 24616 2082 24668
rect 2082 24616 2094 24668
rect 2094 24616 2100 24668
rect 2124 24616 2146 24668
rect 2146 24616 2158 24668
rect 2158 24616 2180 24668
rect 2204 24616 2210 24668
rect 2210 24616 2222 24668
rect 2222 24616 2260 24668
rect 2284 24616 2286 24668
rect 2286 24616 2338 24668
rect 2338 24616 2340 24668
rect 1964 24614 2020 24616
rect 2044 24614 2100 24616
rect 2124 24614 2180 24616
rect 2204 24614 2260 24616
rect 2284 24614 2340 24616
rect 1964 23336 2020 23338
rect 2044 23336 2100 23338
rect 2124 23336 2180 23338
rect 2204 23336 2260 23338
rect 2284 23336 2340 23338
rect 1964 23284 1966 23336
rect 1966 23284 2018 23336
rect 2018 23284 2020 23336
rect 2044 23284 2082 23336
rect 2082 23284 2094 23336
rect 2094 23284 2100 23336
rect 2124 23284 2146 23336
rect 2146 23284 2158 23336
rect 2158 23284 2180 23336
rect 2204 23284 2210 23336
rect 2210 23284 2222 23336
rect 2222 23284 2260 23336
rect 2284 23284 2286 23336
rect 2286 23284 2338 23336
rect 2338 23284 2340 23336
rect 1964 23282 2020 23284
rect 2044 23282 2100 23284
rect 2124 23282 2180 23284
rect 2204 23282 2260 23284
rect 2284 23282 2340 23284
rect 788 23134 844 23190
rect 884 21654 940 21710
rect 1964 22004 2020 22006
rect 2044 22004 2100 22006
rect 2124 22004 2180 22006
rect 2204 22004 2260 22006
rect 2284 22004 2340 22006
rect 1964 21952 1966 22004
rect 1966 21952 2018 22004
rect 2018 21952 2020 22004
rect 2044 21952 2082 22004
rect 2082 21952 2094 22004
rect 2094 21952 2100 22004
rect 2124 21952 2146 22004
rect 2146 21952 2158 22004
rect 2158 21952 2180 22004
rect 2204 21952 2210 22004
rect 2210 21952 2222 22004
rect 2222 21952 2260 22004
rect 2284 21952 2286 22004
rect 2286 21952 2338 22004
rect 2338 21952 2340 22004
rect 1964 21950 2020 21952
rect 2044 21950 2100 21952
rect 2124 21950 2180 21952
rect 2204 21950 2260 21952
rect 2284 21950 2340 21952
rect 1964 20672 2020 20674
rect 2044 20672 2100 20674
rect 2124 20672 2180 20674
rect 2204 20672 2260 20674
rect 2284 20672 2340 20674
rect 1964 20620 1966 20672
rect 1966 20620 2018 20672
rect 2018 20620 2020 20672
rect 2044 20620 2082 20672
rect 2082 20620 2094 20672
rect 2094 20620 2100 20672
rect 2124 20620 2146 20672
rect 2146 20620 2158 20672
rect 2158 20620 2180 20672
rect 2204 20620 2210 20672
rect 2210 20620 2222 20672
rect 2222 20620 2260 20672
rect 2284 20620 2286 20672
rect 2286 20620 2338 20672
rect 2338 20620 2340 20672
rect 1964 20618 2020 20620
rect 2044 20618 2100 20620
rect 2124 20618 2180 20620
rect 2204 20618 2260 20620
rect 2284 20618 2340 20620
rect 1556 20174 1612 20230
rect 1964 19340 2020 19342
rect 2044 19340 2100 19342
rect 2124 19340 2180 19342
rect 2204 19340 2260 19342
rect 2284 19340 2340 19342
rect 1964 19288 1966 19340
rect 1966 19288 2018 19340
rect 2018 19288 2020 19340
rect 2044 19288 2082 19340
rect 2082 19288 2094 19340
rect 2094 19288 2100 19340
rect 2124 19288 2146 19340
rect 2146 19288 2158 19340
rect 2158 19288 2180 19340
rect 2204 19288 2210 19340
rect 2210 19288 2222 19340
rect 2222 19288 2260 19340
rect 2284 19288 2286 19340
rect 2286 19288 2338 19340
rect 2338 19288 2340 19340
rect 1964 19286 2020 19288
rect 2044 19286 2100 19288
rect 2124 19286 2180 19288
rect 2204 19286 2260 19288
rect 2284 19286 2340 19288
rect 1556 18694 1612 18750
rect 1964 18008 2020 18010
rect 2044 18008 2100 18010
rect 2124 18008 2180 18010
rect 2204 18008 2260 18010
rect 2284 18008 2340 18010
rect 1964 17956 1966 18008
rect 1966 17956 2018 18008
rect 2018 17956 2020 18008
rect 2044 17956 2082 18008
rect 2082 17956 2094 18008
rect 2094 17956 2100 18008
rect 2124 17956 2146 18008
rect 2146 17956 2158 18008
rect 2158 17956 2180 18008
rect 2204 17956 2210 18008
rect 2210 17956 2222 18008
rect 2222 17956 2260 18008
rect 2284 17956 2286 18008
rect 2286 17956 2338 18008
rect 2338 17956 2340 18008
rect 1964 17954 2020 17956
rect 2044 17954 2100 17956
rect 2124 17954 2180 17956
rect 2204 17954 2260 17956
rect 2284 17954 2340 17956
rect 1268 17231 1324 17270
rect 1268 17214 1270 17231
rect 1270 17214 1322 17231
rect 1322 17214 1324 17231
rect 1964 16676 2020 16678
rect 2044 16676 2100 16678
rect 2124 16676 2180 16678
rect 2204 16676 2260 16678
rect 2284 16676 2340 16678
rect 1964 16624 1966 16676
rect 1966 16624 2018 16676
rect 2018 16624 2020 16676
rect 2044 16624 2082 16676
rect 2082 16624 2094 16676
rect 2094 16624 2100 16676
rect 2124 16624 2146 16676
rect 2146 16624 2158 16676
rect 2158 16624 2180 16676
rect 2204 16624 2210 16676
rect 2210 16624 2222 16676
rect 2222 16624 2260 16676
rect 2284 16624 2286 16676
rect 2286 16624 2338 16676
rect 2338 16624 2340 16676
rect 1964 16622 2020 16624
rect 2044 16622 2100 16624
rect 2124 16622 2180 16624
rect 2204 16622 2260 16624
rect 2284 16622 2340 16624
rect 788 15751 844 15790
rect 788 15734 790 15751
rect 790 15734 842 15751
rect 842 15734 844 15751
rect 1964 15344 2020 15346
rect 2044 15344 2100 15346
rect 2124 15344 2180 15346
rect 2204 15344 2260 15346
rect 2284 15344 2340 15346
rect 1964 15292 1966 15344
rect 1966 15292 2018 15344
rect 2018 15292 2020 15344
rect 2044 15292 2082 15344
rect 2082 15292 2094 15344
rect 2094 15292 2100 15344
rect 2124 15292 2146 15344
rect 2146 15292 2158 15344
rect 2158 15292 2180 15344
rect 2204 15292 2210 15344
rect 2210 15292 2222 15344
rect 2222 15292 2260 15344
rect 2284 15292 2286 15344
rect 2286 15292 2338 15344
rect 2338 15292 2340 15344
rect 1964 15290 2020 15292
rect 2044 15290 2100 15292
rect 2124 15290 2180 15292
rect 2204 15290 2260 15292
rect 2284 15290 2340 15292
rect 788 14271 844 14310
rect 788 14254 790 14271
rect 790 14254 842 14271
rect 842 14254 844 14271
rect 1964 14012 2020 14014
rect 2044 14012 2100 14014
rect 2124 14012 2180 14014
rect 2204 14012 2260 14014
rect 2284 14012 2340 14014
rect 1964 13960 1966 14012
rect 1966 13960 2018 14012
rect 2018 13960 2020 14012
rect 2044 13960 2082 14012
rect 2082 13960 2094 14012
rect 2094 13960 2100 14012
rect 2124 13960 2146 14012
rect 2146 13960 2158 14012
rect 2158 13960 2180 14012
rect 2204 13960 2210 14012
rect 2210 13960 2222 14012
rect 2222 13960 2260 14012
rect 2284 13960 2286 14012
rect 2286 13960 2338 14012
rect 2338 13960 2340 14012
rect 1964 13958 2020 13960
rect 2044 13958 2100 13960
rect 2124 13958 2180 13960
rect 2204 13958 2260 13960
rect 2284 13958 2340 13960
rect 1556 12774 1612 12830
rect 1964 12680 2020 12682
rect 2044 12680 2100 12682
rect 2124 12680 2180 12682
rect 2204 12680 2260 12682
rect 2284 12680 2340 12682
rect 1964 12628 1966 12680
rect 1966 12628 2018 12680
rect 2018 12628 2020 12680
rect 2044 12628 2082 12680
rect 2082 12628 2094 12680
rect 2094 12628 2100 12680
rect 2124 12628 2146 12680
rect 2146 12628 2158 12680
rect 2158 12628 2180 12680
rect 2204 12628 2210 12680
rect 2210 12628 2222 12680
rect 2222 12628 2260 12680
rect 2284 12628 2286 12680
rect 2286 12628 2338 12680
rect 2338 12628 2340 12680
rect 1964 12626 2020 12628
rect 2044 12626 2100 12628
rect 2124 12626 2180 12628
rect 2204 12626 2260 12628
rect 2284 12626 2340 12628
rect 1556 11294 1612 11350
rect 1964 11348 2020 11350
rect 2044 11348 2100 11350
rect 2124 11348 2180 11350
rect 2204 11348 2260 11350
rect 2284 11348 2340 11350
rect 1964 11296 1966 11348
rect 1966 11296 2018 11348
rect 2018 11296 2020 11348
rect 2044 11296 2082 11348
rect 2082 11296 2094 11348
rect 2094 11296 2100 11348
rect 2124 11296 2146 11348
rect 2146 11296 2158 11348
rect 2158 11296 2180 11348
rect 2204 11296 2210 11348
rect 2210 11296 2222 11348
rect 2222 11296 2260 11348
rect 2284 11296 2286 11348
rect 2286 11296 2338 11348
rect 2338 11296 2340 11348
rect 1964 11294 2020 11296
rect 2044 11294 2100 11296
rect 2124 11294 2180 11296
rect 2204 11294 2260 11296
rect 2284 11294 2340 11296
rect 1556 9814 1612 9870
rect 4964 25334 5020 25336
rect 5044 25334 5100 25336
rect 5124 25334 5180 25336
rect 5204 25334 5260 25336
rect 5284 25334 5340 25336
rect 4964 25282 4966 25334
rect 4966 25282 5018 25334
rect 5018 25282 5020 25334
rect 5044 25282 5082 25334
rect 5082 25282 5094 25334
rect 5094 25282 5100 25334
rect 5124 25282 5146 25334
rect 5146 25282 5158 25334
rect 5158 25282 5180 25334
rect 5204 25282 5210 25334
rect 5210 25282 5222 25334
rect 5222 25282 5260 25334
rect 5284 25282 5286 25334
rect 5286 25282 5338 25334
rect 5338 25282 5340 25334
rect 4964 25280 5020 25282
rect 5044 25280 5100 25282
rect 5124 25280 5180 25282
rect 5204 25280 5260 25282
rect 5284 25280 5340 25282
rect 4964 24002 5020 24004
rect 5044 24002 5100 24004
rect 5124 24002 5180 24004
rect 5204 24002 5260 24004
rect 5284 24002 5340 24004
rect 4964 23950 4966 24002
rect 4966 23950 5018 24002
rect 5018 23950 5020 24002
rect 5044 23950 5082 24002
rect 5082 23950 5094 24002
rect 5094 23950 5100 24002
rect 5124 23950 5146 24002
rect 5146 23950 5158 24002
rect 5158 23950 5180 24002
rect 5204 23950 5210 24002
rect 5210 23950 5222 24002
rect 5222 23950 5260 24002
rect 5284 23950 5286 24002
rect 5286 23950 5338 24002
rect 5338 23950 5340 24002
rect 4964 23948 5020 23950
rect 5044 23948 5100 23950
rect 5124 23948 5180 23950
rect 5204 23948 5260 23950
rect 5284 23948 5340 23950
rect 4964 22670 5020 22672
rect 5044 22670 5100 22672
rect 5124 22670 5180 22672
rect 5204 22670 5260 22672
rect 5284 22670 5340 22672
rect 4964 22618 4966 22670
rect 4966 22618 5018 22670
rect 5018 22618 5020 22670
rect 5044 22618 5082 22670
rect 5082 22618 5094 22670
rect 5094 22618 5100 22670
rect 5124 22618 5146 22670
rect 5146 22618 5158 22670
rect 5158 22618 5180 22670
rect 5204 22618 5210 22670
rect 5210 22618 5222 22670
rect 5222 22618 5260 22670
rect 5284 22618 5286 22670
rect 5286 22618 5338 22670
rect 5338 22618 5340 22670
rect 4964 22616 5020 22618
rect 5044 22616 5100 22618
rect 5124 22616 5180 22618
rect 5204 22616 5260 22618
rect 5284 22616 5340 22618
rect 4964 21338 5020 21340
rect 5044 21338 5100 21340
rect 5124 21338 5180 21340
rect 5204 21338 5260 21340
rect 5284 21338 5340 21340
rect 4964 21286 4966 21338
rect 4966 21286 5018 21338
rect 5018 21286 5020 21338
rect 5044 21286 5082 21338
rect 5082 21286 5094 21338
rect 5094 21286 5100 21338
rect 5124 21286 5146 21338
rect 5146 21286 5158 21338
rect 5158 21286 5180 21338
rect 5204 21286 5210 21338
rect 5210 21286 5222 21338
rect 5222 21286 5260 21338
rect 5284 21286 5286 21338
rect 5286 21286 5338 21338
rect 5338 21286 5340 21338
rect 4964 21284 5020 21286
rect 5044 21284 5100 21286
rect 5124 21284 5180 21286
rect 5204 21284 5260 21286
rect 5284 21284 5340 21286
rect 4964 20006 5020 20008
rect 5044 20006 5100 20008
rect 5124 20006 5180 20008
rect 5204 20006 5260 20008
rect 5284 20006 5340 20008
rect 4964 19954 4966 20006
rect 4966 19954 5018 20006
rect 5018 19954 5020 20006
rect 5044 19954 5082 20006
rect 5082 19954 5094 20006
rect 5094 19954 5100 20006
rect 5124 19954 5146 20006
rect 5146 19954 5158 20006
rect 5158 19954 5180 20006
rect 5204 19954 5210 20006
rect 5210 19954 5222 20006
rect 5222 19954 5260 20006
rect 5284 19954 5286 20006
rect 5286 19954 5338 20006
rect 5338 19954 5340 20006
rect 4964 19952 5020 19954
rect 5044 19952 5100 19954
rect 5124 19952 5180 19954
rect 5204 19952 5260 19954
rect 5284 19952 5340 19954
rect 4964 18674 5020 18676
rect 5044 18674 5100 18676
rect 5124 18674 5180 18676
rect 5204 18674 5260 18676
rect 5284 18674 5340 18676
rect 4964 18622 4966 18674
rect 4966 18622 5018 18674
rect 5018 18622 5020 18674
rect 5044 18622 5082 18674
rect 5082 18622 5094 18674
rect 5094 18622 5100 18674
rect 5124 18622 5146 18674
rect 5146 18622 5158 18674
rect 5158 18622 5180 18674
rect 5204 18622 5210 18674
rect 5210 18622 5222 18674
rect 5222 18622 5260 18674
rect 5284 18622 5286 18674
rect 5286 18622 5338 18674
rect 5338 18622 5340 18674
rect 4964 18620 5020 18622
rect 5044 18620 5100 18622
rect 5124 18620 5180 18622
rect 5204 18620 5260 18622
rect 5284 18620 5340 18622
rect 4964 17342 5020 17344
rect 5044 17342 5100 17344
rect 5124 17342 5180 17344
rect 5204 17342 5260 17344
rect 5284 17342 5340 17344
rect 4964 17290 4966 17342
rect 4966 17290 5018 17342
rect 5018 17290 5020 17342
rect 5044 17290 5082 17342
rect 5082 17290 5094 17342
rect 5094 17290 5100 17342
rect 5124 17290 5146 17342
rect 5146 17290 5158 17342
rect 5158 17290 5180 17342
rect 5204 17290 5210 17342
rect 5210 17290 5222 17342
rect 5222 17290 5260 17342
rect 5284 17290 5286 17342
rect 5286 17290 5338 17342
rect 5338 17290 5340 17342
rect 4964 17288 5020 17290
rect 5044 17288 5100 17290
rect 5124 17288 5180 17290
rect 5204 17288 5260 17290
rect 5284 17288 5340 17290
rect 4964 16010 5020 16012
rect 5044 16010 5100 16012
rect 5124 16010 5180 16012
rect 5204 16010 5260 16012
rect 5284 16010 5340 16012
rect 4964 15958 4966 16010
rect 4966 15958 5018 16010
rect 5018 15958 5020 16010
rect 5044 15958 5082 16010
rect 5082 15958 5094 16010
rect 5094 15958 5100 16010
rect 5124 15958 5146 16010
rect 5146 15958 5158 16010
rect 5158 15958 5180 16010
rect 5204 15958 5210 16010
rect 5210 15958 5222 16010
rect 5222 15958 5260 16010
rect 5284 15958 5286 16010
rect 5286 15958 5338 16010
rect 5338 15958 5340 16010
rect 4964 15956 5020 15958
rect 5044 15956 5100 15958
rect 5124 15956 5180 15958
rect 5204 15956 5260 15958
rect 5284 15956 5340 15958
rect 4964 14678 5020 14680
rect 5044 14678 5100 14680
rect 5124 14678 5180 14680
rect 5204 14678 5260 14680
rect 5284 14678 5340 14680
rect 4964 14626 4966 14678
rect 4966 14626 5018 14678
rect 5018 14626 5020 14678
rect 5044 14626 5082 14678
rect 5082 14626 5094 14678
rect 5094 14626 5100 14678
rect 5124 14626 5146 14678
rect 5146 14626 5158 14678
rect 5158 14626 5180 14678
rect 5204 14626 5210 14678
rect 5210 14626 5222 14678
rect 5222 14626 5260 14678
rect 5284 14626 5286 14678
rect 5286 14626 5338 14678
rect 5338 14626 5340 14678
rect 4964 14624 5020 14626
rect 5044 14624 5100 14626
rect 5124 14624 5180 14626
rect 5204 14624 5260 14626
rect 5284 14624 5340 14626
rect 4964 13346 5020 13348
rect 5044 13346 5100 13348
rect 5124 13346 5180 13348
rect 5204 13346 5260 13348
rect 5284 13346 5340 13348
rect 4964 13294 4966 13346
rect 4966 13294 5018 13346
rect 5018 13294 5020 13346
rect 5044 13294 5082 13346
rect 5082 13294 5094 13346
rect 5094 13294 5100 13346
rect 5124 13294 5146 13346
rect 5146 13294 5158 13346
rect 5158 13294 5180 13346
rect 5204 13294 5210 13346
rect 5210 13294 5222 13346
rect 5222 13294 5260 13346
rect 5284 13294 5286 13346
rect 5286 13294 5338 13346
rect 5338 13294 5340 13346
rect 4964 13292 5020 13294
rect 5044 13292 5100 13294
rect 5124 13292 5180 13294
rect 5204 13292 5260 13294
rect 5284 13292 5340 13294
rect 1652 8334 1708 8390
rect 1964 10016 2020 10018
rect 2044 10016 2100 10018
rect 2124 10016 2180 10018
rect 2204 10016 2260 10018
rect 2284 10016 2340 10018
rect 1964 9964 1966 10016
rect 1966 9964 2018 10016
rect 2018 9964 2020 10016
rect 2044 9964 2082 10016
rect 2082 9964 2094 10016
rect 2094 9964 2100 10016
rect 2124 9964 2146 10016
rect 2146 9964 2158 10016
rect 2158 9964 2180 10016
rect 2204 9964 2210 10016
rect 2210 9964 2222 10016
rect 2222 9964 2260 10016
rect 2284 9964 2286 10016
rect 2286 9964 2338 10016
rect 2338 9964 2340 10016
rect 1964 9962 2020 9964
rect 2044 9962 2100 9964
rect 2124 9962 2180 9964
rect 2204 9962 2260 9964
rect 2284 9962 2340 9964
rect 1964 8684 2020 8686
rect 2044 8684 2100 8686
rect 2124 8684 2180 8686
rect 2204 8684 2260 8686
rect 2284 8684 2340 8686
rect 1964 8632 1966 8684
rect 1966 8632 2018 8684
rect 2018 8632 2020 8684
rect 2044 8632 2082 8684
rect 2082 8632 2094 8684
rect 2094 8632 2100 8684
rect 2124 8632 2146 8684
rect 2146 8632 2158 8684
rect 2158 8632 2180 8684
rect 2204 8632 2210 8684
rect 2210 8632 2222 8684
rect 2222 8632 2260 8684
rect 2284 8632 2286 8684
rect 2286 8632 2338 8684
rect 2338 8632 2340 8684
rect 1964 8630 2020 8632
rect 2044 8630 2100 8632
rect 2124 8630 2180 8632
rect 2204 8630 2260 8632
rect 2284 8630 2340 8632
rect 4964 12014 5020 12016
rect 5044 12014 5100 12016
rect 5124 12014 5180 12016
rect 5204 12014 5260 12016
rect 5284 12014 5340 12016
rect 4964 11962 4966 12014
rect 4966 11962 5018 12014
rect 5018 11962 5020 12014
rect 5044 11962 5082 12014
rect 5082 11962 5094 12014
rect 5094 11962 5100 12014
rect 5124 11962 5146 12014
rect 5146 11962 5158 12014
rect 5158 11962 5180 12014
rect 5204 11962 5210 12014
rect 5210 11962 5222 12014
rect 5222 11962 5260 12014
rect 5284 11962 5286 12014
rect 5286 11962 5338 12014
rect 5338 11962 5340 12014
rect 4964 11960 5020 11962
rect 5044 11960 5100 11962
rect 5124 11960 5180 11962
rect 5204 11960 5260 11962
rect 5284 11960 5340 11962
rect 1652 6854 1708 6910
rect 1964 7352 2020 7354
rect 2044 7352 2100 7354
rect 2124 7352 2180 7354
rect 2204 7352 2260 7354
rect 2284 7352 2340 7354
rect 1964 7300 1966 7352
rect 1966 7300 2018 7352
rect 2018 7300 2020 7352
rect 2044 7300 2082 7352
rect 2082 7300 2094 7352
rect 2094 7300 2100 7352
rect 2124 7300 2146 7352
rect 2146 7300 2158 7352
rect 2158 7300 2180 7352
rect 2204 7300 2210 7352
rect 2210 7300 2222 7352
rect 2222 7300 2260 7352
rect 2284 7300 2286 7352
rect 2286 7300 2338 7352
rect 2338 7300 2340 7352
rect 1964 7298 2020 7300
rect 2044 7298 2100 7300
rect 2124 7298 2180 7300
rect 2204 7298 2260 7300
rect 2284 7298 2340 7300
rect 1964 6020 2020 6022
rect 2044 6020 2100 6022
rect 2124 6020 2180 6022
rect 2204 6020 2260 6022
rect 2284 6020 2340 6022
rect 1964 5968 1966 6020
rect 1966 5968 2018 6020
rect 2018 5968 2020 6020
rect 2044 5968 2082 6020
rect 2082 5968 2094 6020
rect 2094 5968 2100 6020
rect 2124 5968 2146 6020
rect 2146 5968 2158 6020
rect 2158 5968 2180 6020
rect 2204 5968 2210 6020
rect 2210 5968 2222 6020
rect 2222 5968 2260 6020
rect 2284 5968 2286 6020
rect 2286 5968 2338 6020
rect 2338 5968 2340 6020
rect 1964 5966 2020 5968
rect 2044 5966 2100 5968
rect 2124 5966 2180 5968
rect 2204 5966 2260 5968
rect 2284 5966 2340 5968
rect 1964 4688 2020 4690
rect 2044 4688 2100 4690
rect 2124 4688 2180 4690
rect 2204 4688 2260 4690
rect 2284 4688 2340 4690
rect 1964 4636 1966 4688
rect 1966 4636 2018 4688
rect 2018 4636 2020 4688
rect 2044 4636 2082 4688
rect 2082 4636 2094 4688
rect 2094 4636 2100 4688
rect 2124 4636 2146 4688
rect 2146 4636 2158 4688
rect 2158 4636 2180 4688
rect 2204 4636 2210 4688
rect 2210 4636 2222 4688
rect 2222 4636 2260 4688
rect 2284 4636 2286 4688
rect 2286 4636 2338 4688
rect 2338 4636 2340 4688
rect 1964 4634 2020 4636
rect 2044 4634 2100 4636
rect 2124 4634 2180 4636
rect 2204 4634 2260 4636
rect 2284 4634 2340 4636
rect 884 3894 940 3950
rect 1964 3356 2020 3358
rect 2044 3356 2100 3358
rect 2124 3356 2180 3358
rect 2204 3356 2260 3358
rect 2284 3356 2340 3358
rect 1964 3304 1966 3356
rect 1966 3304 2018 3356
rect 2018 3304 2020 3356
rect 2044 3304 2082 3356
rect 2082 3304 2094 3356
rect 2094 3304 2100 3356
rect 2124 3304 2146 3356
rect 2146 3304 2158 3356
rect 2158 3304 2180 3356
rect 2204 3304 2210 3356
rect 2210 3304 2222 3356
rect 2222 3304 2260 3356
rect 2284 3304 2286 3356
rect 2286 3304 2338 3356
rect 2338 3304 2340 3356
rect 1964 3302 2020 3304
rect 2044 3302 2100 3304
rect 2124 3302 2180 3304
rect 2204 3302 2260 3304
rect 2284 3302 2340 3304
rect 4964 10682 5020 10684
rect 5044 10682 5100 10684
rect 5124 10682 5180 10684
rect 5204 10682 5260 10684
rect 5284 10682 5340 10684
rect 4964 10630 4966 10682
rect 4966 10630 5018 10682
rect 5018 10630 5020 10682
rect 5044 10630 5082 10682
rect 5082 10630 5094 10682
rect 5094 10630 5100 10682
rect 5124 10630 5146 10682
rect 5146 10630 5158 10682
rect 5158 10630 5180 10682
rect 5204 10630 5210 10682
rect 5210 10630 5222 10682
rect 5222 10630 5260 10682
rect 5284 10630 5286 10682
rect 5286 10630 5338 10682
rect 5338 10630 5340 10682
rect 4964 10628 5020 10630
rect 5044 10628 5100 10630
rect 5124 10628 5180 10630
rect 5204 10628 5260 10630
rect 5284 10628 5340 10630
rect 4964 9350 5020 9352
rect 5044 9350 5100 9352
rect 5124 9350 5180 9352
rect 5204 9350 5260 9352
rect 5284 9350 5340 9352
rect 4964 9298 4966 9350
rect 4966 9298 5018 9350
rect 5018 9298 5020 9350
rect 5044 9298 5082 9350
rect 5082 9298 5094 9350
rect 5094 9298 5100 9350
rect 5124 9298 5146 9350
rect 5146 9298 5158 9350
rect 5158 9298 5180 9350
rect 5204 9298 5210 9350
rect 5210 9298 5222 9350
rect 5222 9298 5260 9350
rect 5284 9298 5286 9350
rect 5286 9298 5338 9350
rect 5338 9298 5340 9350
rect 4964 9296 5020 9298
rect 5044 9296 5100 9298
rect 5124 9296 5180 9298
rect 5204 9296 5260 9298
rect 5284 9296 5340 9298
rect 4964 8018 5020 8020
rect 5044 8018 5100 8020
rect 5124 8018 5180 8020
rect 5204 8018 5260 8020
rect 5284 8018 5340 8020
rect 4964 7966 4966 8018
rect 4966 7966 5018 8018
rect 5018 7966 5020 8018
rect 5044 7966 5082 8018
rect 5082 7966 5094 8018
rect 5094 7966 5100 8018
rect 5124 7966 5146 8018
rect 5146 7966 5158 8018
rect 5158 7966 5180 8018
rect 5204 7966 5210 8018
rect 5210 7966 5222 8018
rect 5222 7966 5260 8018
rect 5284 7966 5286 8018
rect 5286 7966 5338 8018
rect 5338 7966 5340 8018
rect 4964 7964 5020 7966
rect 5044 7964 5100 7966
rect 5124 7964 5180 7966
rect 5204 7964 5260 7966
rect 5284 7964 5340 7966
rect 4964 6686 5020 6688
rect 5044 6686 5100 6688
rect 5124 6686 5180 6688
rect 5204 6686 5260 6688
rect 5284 6686 5340 6688
rect 4964 6634 4966 6686
rect 4966 6634 5018 6686
rect 5018 6634 5020 6686
rect 5044 6634 5082 6686
rect 5082 6634 5094 6686
rect 5094 6634 5100 6686
rect 5124 6634 5146 6686
rect 5146 6634 5158 6686
rect 5158 6634 5180 6686
rect 5204 6634 5210 6686
rect 5210 6634 5222 6686
rect 5222 6634 5260 6686
rect 5284 6634 5286 6686
rect 5286 6634 5338 6686
rect 5338 6634 5340 6686
rect 4964 6632 5020 6634
rect 5044 6632 5100 6634
rect 5124 6632 5180 6634
rect 5204 6632 5260 6634
rect 5284 6632 5340 6634
rect 4964 5354 5020 5356
rect 5044 5354 5100 5356
rect 5124 5354 5180 5356
rect 5204 5354 5260 5356
rect 5284 5354 5340 5356
rect 4964 5302 4966 5354
rect 4966 5302 5018 5354
rect 5018 5302 5020 5354
rect 5044 5302 5082 5354
rect 5082 5302 5094 5354
rect 5094 5302 5100 5354
rect 5124 5302 5146 5354
rect 5146 5302 5158 5354
rect 5158 5302 5180 5354
rect 5204 5302 5210 5354
rect 5210 5302 5222 5354
rect 5222 5302 5260 5354
rect 5284 5302 5286 5354
rect 5286 5302 5338 5354
rect 5338 5302 5340 5354
rect 4964 5300 5020 5302
rect 5044 5300 5100 5302
rect 5124 5300 5180 5302
rect 5204 5300 5260 5302
rect 5284 5300 5340 5302
rect 4964 4022 5020 4024
rect 5044 4022 5100 4024
rect 5124 4022 5180 4024
rect 5204 4022 5260 4024
rect 5284 4022 5340 4024
rect 4964 3970 4966 4022
rect 4966 3970 5018 4022
rect 5018 3970 5020 4022
rect 5044 3970 5082 4022
rect 5082 3970 5094 4022
rect 5094 3970 5100 4022
rect 5124 3970 5146 4022
rect 5146 3970 5158 4022
rect 5158 3970 5180 4022
rect 5204 3970 5210 4022
rect 5210 3970 5222 4022
rect 5222 3970 5260 4022
rect 5284 3970 5286 4022
rect 5286 3970 5338 4022
rect 5338 3970 5340 4022
rect 4964 3968 5020 3970
rect 5044 3968 5100 3970
rect 5124 3968 5180 3970
rect 5204 3968 5260 3970
rect 5284 3968 5340 3970
rect 7964 24668 8020 24670
rect 8044 24668 8100 24670
rect 8124 24668 8180 24670
rect 8204 24668 8260 24670
rect 8284 24668 8340 24670
rect 7964 24616 7966 24668
rect 7966 24616 8018 24668
rect 8018 24616 8020 24668
rect 8044 24616 8082 24668
rect 8082 24616 8094 24668
rect 8094 24616 8100 24668
rect 8124 24616 8146 24668
rect 8146 24616 8158 24668
rect 8158 24616 8180 24668
rect 8204 24616 8210 24668
rect 8210 24616 8222 24668
rect 8222 24616 8260 24668
rect 8284 24616 8286 24668
rect 8286 24616 8338 24668
rect 8338 24616 8340 24668
rect 7964 24614 8020 24616
rect 8044 24614 8100 24616
rect 8124 24614 8180 24616
rect 8204 24614 8260 24616
rect 8284 24614 8340 24616
rect 7964 23336 8020 23338
rect 8044 23336 8100 23338
rect 8124 23336 8180 23338
rect 8204 23336 8260 23338
rect 8284 23336 8340 23338
rect 7964 23284 7966 23336
rect 7966 23284 8018 23336
rect 8018 23284 8020 23336
rect 8044 23284 8082 23336
rect 8082 23284 8094 23336
rect 8094 23284 8100 23336
rect 8124 23284 8146 23336
rect 8146 23284 8158 23336
rect 8158 23284 8180 23336
rect 8204 23284 8210 23336
rect 8210 23284 8222 23336
rect 8222 23284 8260 23336
rect 8284 23284 8286 23336
rect 8286 23284 8338 23336
rect 8338 23284 8340 23336
rect 7964 23282 8020 23284
rect 8044 23282 8100 23284
rect 8124 23282 8180 23284
rect 8204 23282 8260 23284
rect 8284 23282 8340 23284
rect 10100 22542 10156 22598
rect 7964 22004 8020 22006
rect 8044 22004 8100 22006
rect 8124 22004 8180 22006
rect 8204 22004 8260 22006
rect 8284 22004 8340 22006
rect 7964 21952 7966 22004
rect 7966 21952 8018 22004
rect 8018 21952 8020 22004
rect 8044 21952 8082 22004
rect 8082 21952 8094 22004
rect 8094 21952 8100 22004
rect 8124 21952 8146 22004
rect 8146 21952 8158 22004
rect 8158 21952 8180 22004
rect 8204 21952 8210 22004
rect 8210 21952 8222 22004
rect 8222 21952 8260 22004
rect 8284 21952 8286 22004
rect 8286 21952 8338 22004
rect 8338 21952 8340 22004
rect 7964 21950 8020 21952
rect 8044 21950 8100 21952
rect 8124 21950 8180 21952
rect 8204 21950 8260 21952
rect 8284 21950 8340 21952
rect 7964 20672 8020 20674
rect 8044 20672 8100 20674
rect 8124 20672 8180 20674
rect 8204 20672 8260 20674
rect 8284 20672 8340 20674
rect 7964 20620 7966 20672
rect 7966 20620 8018 20672
rect 8018 20620 8020 20672
rect 8044 20620 8082 20672
rect 8082 20620 8094 20672
rect 8094 20620 8100 20672
rect 8124 20620 8146 20672
rect 8146 20620 8158 20672
rect 8158 20620 8180 20672
rect 8204 20620 8210 20672
rect 8210 20620 8222 20672
rect 8222 20620 8260 20672
rect 8284 20620 8286 20672
rect 8286 20620 8338 20672
rect 8338 20620 8340 20672
rect 7964 20618 8020 20620
rect 8044 20618 8100 20620
rect 8124 20618 8180 20620
rect 8204 20618 8260 20620
rect 8284 20618 8340 20620
rect 10100 20191 10156 20230
rect 10100 20174 10102 20191
rect 10102 20174 10154 20191
rect 10154 20174 10156 20191
rect 7964 19340 8020 19342
rect 8044 19340 8100 19342
rect 8124 19340 8180 19342
rect 8204 19340 8260 19342
rect 8284 19340 8340 19342
rect 7964 19288 7966 19340
rect 7966 19288 8018 19340
rect 8018 19288 8020 19340
rect 8044 19288 8082 19340
rect 8082 19288 8094 19340
rect 8094 19288 8100 19340
rect 8124 19288 8146 19340
rect 8146 19288 8158 19340
rect 8158 19288 8180 19340
rect 8204 19288 8210 19340
rect 8210 19288 8222 19340
rect 8222 19288 8260 19340
rect 8284 19288 8286 19340
rect 8286 19288 8338 19340
rect 8338 19288 8340 19340
rect 7964 19286 8020 19288
rect 8044 19286 8100 19288
rect 8124 19286 8180 19288
rect 8204 19286 8260 19288
rect 8284 19286 8340 19288
rect 7964 18008 8020 18010
rect 8044 18008 8100 18010
rect 8124 18008 8180 18010
rect 8204 18008 8260 18010
rect 8284 18008 8340 18010
rect 7964 17956 7966 18008
rect 7966 17956 8018 18008
rect 8018 17956 8020 18008
rect 8044 17956 8082 18008
rect 8082 17956 8094 18008
rect 8094 17956 8100 18008
rect 8124 17956 8146 18008
rect 8146 17956 8158 18008
rect 8158 17956 8180 18008
rect 8204 17956 8210 18008
rect 8210 17956 8222 18008
rect 8222 17956 8260 18008
rect 8284 17956 8286 18008
rect 8286 17956 8338 18008
rect 8338 17956 8340 18008
rect 7964 17954 8020 17956
rect 8044 17954 8100 17956
rect 8124 17954 8180 17956
rect 8204 17954 8260 17956
rect 8284 17954 8340 17956
rect 7964 16676 8020 16678
rect 8044 16676 8100 16678
rect 8124 16676 8180 16678
rect 8204 16676 8260 16678
rect 8284 16676 8340 16678
rect 7964 16624 7966 16676
rect 7966 16624 8018 16676
rect 8018 16624 8020 16676
rect 8044 16624 8082 16676
rect 8082 16624 8094 16676
rect 8094 16624 8100 16676
rect 8124 16624 8146 16676
rect 8146 16624 8158 16676
rect 8158 16624 8180 16676
rect 8204 16624 8210 16676
rect 8210 16624 8222 16676
rect 8222 16624 8260 16676
rect 8284 16624 8286 16676
rect 8286 16624 8338 16676
rect 8338 16624 8340 16676
rect 7964 16622 8020 16624
rect 8044 16622 8100 16624
rect 8124 16622 8180 16624
rect 8204 16622 8260 16624
rect 8284 16622 8340 16624
rect 7964 15344 8020 15346
rect 8044 15344 8100 15346
rect 8124 15344 8180 15346
rect 8204 15344 8260 15346
rect 8284 15344 8340 15346
rect 7964 15292 7966 15344
rect 7966 15292 8018 15344
rect 8018 15292 8020 15344
rect 8044 15292 8082 15344
rect 8082 15292 8094 15344
rect 8094 15292 8100 15344
rect 8124 15292 8146 15344
rect 8146 15292 8158 15344
rect 8158 15292 8180 15344
rect 8204 15292 8210 15344
rect 8210 15292 8222 15344
rect 8222 15292 8260 15344
rect 8284 15292 8286 15344
rect 8286 15292 8338 15344
rect 8338 15292 8340 15344
rect 7964 15290 8020 15292
rect 8044 15290 8100 15292
rect 8124 15290 8180 15292
rect 8204 15290 8260 15292
rect 8284 15290 8340 15292
rect 6356 5522 6412 5578
rect 7964 14012 8020 14014
rect 8044 14012 8100 14014
rect 8124 14012 8180 14014
rect 8204 14012 8260 14014
rect 8284 14012 8340 14014
rect 7964 13960 7966 14012
rect 7966 13960 8018 14012
rect 8018 13960 8020 14012
rect 8044 13960 8082 14012
rect 8082 13960 8094 14012
rect 8094 13960 8100 14012
rect 8124 13960 8146 14012
rect 8146 13960 8158 14012
rect 8158 13960 8180 14012
rect 8204 13960 8210 14012
rect 8210 13960 8222 14012
rect 8222 13960 8260 14012
rect 8284 13960 8286 14012
rect 8286 13960 8338 14012
rect 8338 13960 8340 14012
rect 7964 13958 8020 13960
rect 8044 13958 8100 13960
rect 8124 13958 8180 13960
rect 8204 13958 8260 13960
rect 8284 13958 8340 13960
rect 7964 12680 8020 12682
rect 8044 12680 8100 12682
rect 8124 12680 8180 12682
rect 8204 12680 8260 12682
rect 8284 12680 8340 12682
rect 7964 12628 7966 12680
rect 7966 12628 8018 12680
rect 8018 12628 8020 12680
rect 8044 12628 8082 12680
rect 8082 12628 8094 12680
rect 8094 12628 8100 12680
rect 8124 12628 8146 12680
rect 8146 12628 8158 12680
rect 8158 12628 8180 12680
rect 8204 12628 8210 12680
rect 8210 12628 8222 12680
rect 8222 12628 8260 12680
rect 8284 12628 8286 12680
rect 8286 12628 8338 12680
rect 8338 12628 8340 12680
rect 7964 12626 8020 12628
rect 8044 12626 8100 12628
rect 8124 12626 8180 12628
rect 8204 12626 8260 12628
rect 8284 12626 8340 12628
rect 7964 11348 8020 11350
rect 8044 11348 8100 11350
rect 8124 11348 8180 11350
rect 8204 11348 8260 11350
rect 8284 11348 8340 11350
rect 7964 11296 7966 11348
rect 7966 11296 8018 11348
rect 8018 11296 8020 11348
rect 8044 11296 8082 11348
rect 8082 11296 8094 11348
rect 8094 11296 8100 11348
rect 8124 11296 8146 11348
rect 8146 11296 8158 11348
rect 8158 11296 8180 11348
rect 8204 11296 8210 11348
rect 8210 11296 8222 11348
rect 8222 11296 8260 11348
rect 8284 11296 8286 11348
rect 8286 11296 8338 11348
rect 8338 11296 8340 11348
rect 7964 11294 8020 11296
rect 8044 11294 8100 11296
rect 8124 11294 8180 11296
rect 8204 11294 8260 11296
rect 8284 11294 8340 11296
rect 7964 10016 8020 10018
rect 8044 10016 8100 10018
rect 8124 10016 8180 10018
rect 8204 10016 8260 10018
rect 8284 10016 8340 10018
rect 7964 9964 7966 10016
rect 7966 9964 8018 10016
rect 8018 9964 8020 10016
rect 8044 9964 8082 10016
rect 8082 9964 8094 10016
rect 8094 9964 8100 10016
rect 8124 9964 8146 10016
rect 8146 9964 8158 10016
rect 8158 9964 8180 10016
rect 8204 9964 8210 10016
rect 8210 9964 8222 10016
rect 8222 9964 8260 10016
rect 8284 9964 8286 10016
rect 8286 9964 8338 10016
rect 8338 9964 8340 10016
rect 7964 9962 8020 9964
rect 8044 9962 8100 9964
rect 8124 9962 8180 9964
rect 8204 9962 8260 9964
rect 8284 9962 8340 9964
rect 7964 8684 8020 8686
rect 8044 8684 8100 8686
rect 8124 8684 8180 8686
rect 8204 8684 8260 8686
rect 8284 8684 8340 8686
rect 7964 8632 7966 8684
rect 7966 8632 8018 8684
rect 8018 8632 8020 8684
rect 8044 8632 8082 8684
rect 8082 8632 8094 8684
rect 8094 8632 8100 8684
rect 8124 8632 8146 8684
rect 8146 8632 8158 8684
rect 8158 8632 8180 8684
rect 8204 8632 8210 8684
rect 8210 8632 8222 8684
rect 8222 8632 8260 8684
rect 8284 8632 8286 8684
rect 8286 8632 8338 8684
rect 8338 8632 8340 8684
rect 7964 8630 8020 8632
rect 8044 8630 8100 8632
rect 8124 8630 8180 8632
rect 8204 8630 8260 8632
rect 8284 8630 8340 8632
rect 7964 7352 8020 7354
rect 8044 7352 8100 7354
rect 8124 7352 8180 7354
rect 8204 7352 8260 7354
rect 8284 7352 8340 7354
rect 7964 7300 7966 7352
rect 7966 7300 8018 7352
rect 8018 7300 8020 7352
rect 8044 7300 8082 7352
rect 8082 7300 8094 7352
rect 8094 7300 8100 7352
rect 8124 7300 8146 7352
rect 8146 7300 8158 7352
rect 8158 7300 8180 7352
rect 8204 7300 8210 7352
rect 8210 7300 8222 7352
rect 8222 7300 8260 7352
rect 8284 7300 8286 7352
rect 8286 7300 8338 7352
rect 8338 7300 8340 7352
rect 7964 7298 8020 7300
rect 8044 7298 8100 7300
rect 8124 7298 8180 7300
rect 8204 7298 8260 7300
rect 8284 7298 8340 7300
rect 2228 2414 2284 2470
rect 4964 2690 5020 2692
rect 5044 2690 5100 2692
rect 5124 2690 5180 2692
rect 5204 2690 5260 2692
rect 5284 2690 5340 2692
rect 4964 2638 4966 2690
rect 4966 2638 5018 2690
rect 5018 2638 5020 2690
rect 5044 2638 5082 2690
rect 5082 2638 5094 2690
rect 5094 2638 5100 2690
rect 5124 2638 5146 2690
rect 5146 2638 5158 2690
rect 5158 2638 5180 2690
rect 5204 2638 5210 2690
rect 5210 2638 5222 2690
rect 5222 2638 5260 2690
rect 5284 2638 5286 2690
rect 5286 2638 5338 2690
rect 5338 2638 5340 2690
rect 4964 2636 5020 2638
rect 5044 2636 5100 2638
rect 5124 2636 5180 2638
rect 5204 2636 5260 2638
rect 5284 2636 5340 2638
rect 7964 6020 8020 6022
rect 8044 6020 8100 6022
rect 8124 6020 8180 6022
rect 8204 6020 8260 6022
rect 8284 6020 8340 6022
rect 7964 5968 7966 6020
rect 7966 5968 8018 6020
rect 8018 5968 8020 6020
rect 8044 5968 8082 6020
rect 8082 5968 8094 6020
rect 8094 5968 8100 6020
rect 8124 5968 8146 6020
rect 8146 5968 8158 6020
rect 8158 5968 8180 6020
rect 8204 5968 8210 6020
rect 8210 5968 8222 6020
rect 8222 5968 8260 6020
rect 8284 5968 8286 6020
rect 8286 5968 8338 6020
rect 8338 5968 8340 6020
rect 7964 5966 8020 5968
rect 8044 5966 8100 5968
rect 8124 5966 8180 5968
rect 8204 5966 8260 5968
rect 8284 5966 8340 5968
rect 7964 4688 8020 4690
rect 8044 4688 8100 4690
rect 8124 4688 8180 4690
rect 8204 4688 8260 4690
rect 8284 4688 8340 4690
rect 7964 4636 7966 4688
rect 7966 4636 8018 4688
rect 8018 4636 8020 4688
rect 8044 4636 8082 4688
rect 8082 4636 8094 4688
rect 8094 4636 8100 4688
rect 8124 4636 8146 4688
rect 8146 4636 8158 4688
rect 8158 4636 8180 4688
rect 8204 4636 8210 4688
rect 8210 4636 8222 4688
rect 8222 4636 8260 4688
rect 8284 4636 8286 4688
rect 8286 4636 8338 4688
rect 8338 4636 8340 4688
rect 7964 4634 8020 4636
rect 8044 4634 8100 4636
rect 8124 4634 8180 4636
rect 8204 4634 8260 4636
rect 8284 4634 8340 4636
rect 10100 17823 10156 17862
rect 10100 17806 10102 17823
rect 10102 17806 10154 17823
rect 10154 17806 10156 17823
rect 10100 15455 10156 15494
rect 10100 15438 10102 15455
rect 10102 15438 10154 15455
rect 10154 15438 10156 15455
rect 10100 13070 10156 13126
rect 10100 10741 10102 10758
rect 10102 10741 10154 10758
rect 10154 10741 10156 10758
rect 10100 10702 10156 10741
rect 7964 3356 8020 3358
rect 8044 3356 8100 3358
rect 8124 3356 8180 3358
rect 8204 3356 8260 3358
rect 8284 3356 8340 3358
rect 7964 3304 7966 3356
rect 7966 3304 8018 3356
rect 8018 3304 8020 3356
rect 8044 3304 8082 3356
rect 8082 3304 8094 3356
rect 8094 3304 8100 3356
rect 8124 3304 8146 3356
rect 8146 3304 8158 3356
rect 8158 3304 8180 3356
rect 8204 3304 8210 3356
rect 8210 3304 8222 3356
rect 8222 3304 8260 3356
rect 8284 3304 8286 3356
rect 8286 3304 8338 3356
rect 8338 3304 8340 3356
rect 7964 3302 8020 3304
rect 8044 3302 8100 3304
rect 8124 3302 8180 3304
rect 8204 3302 8260 3304
rect 8284 3302 8340 3304
rect 10100 8351 10156 8390
rect 10100 8334 10102 8351
rect 10102 8334 10154 8351
rect 10154 8334 10156 8351
rect 10100 5966 10156 6022
rect 10100 3615 10156 3654
rect 10100 3598 10102 3615
rect 10102 3598 10154 3615
rect 10154 3598 10156 3615
rect 9716 1230 9772 1286
<< metal3 >>
rect 9711 27336 9777 27339
rect 10922 27336 11722 27366
rect 9711 27334 11722 27336
rect 9711 27278 9716 27334
rect 9772 27278 11722 27334
rect 9711 27276 11722 27278
rect 9711 27273 9777 27276
rect 10922 27246 11722 27276
rect 0 26152 800 26182
rect 1647 26152 1713 26155
rect 0 26150 1713 26152
rect 0 26094 1652 26150
rect 1708 26094 1713 26150
rect 0 26092 1713 26094
rect 0 26062 800 26092
rect 1647 26089 1713 26092
rect 1954 26006 2350 26007
rect 1954 25942 1960 26006
rect 2024 25942 2040 26006
rect 2104 25942 2120 26006
rect 2184 25942 2200 26006
rect 2264 25942 2280 26006
rect 2344 25942 2350 26006
rect 1954 25941 2350 25942
rect 7954 26006 8350 26007
rect 7954 25942 7960 26006
rect 8024 25942 8040 26006
rect 8104 25942 8120 26006
rect 8184 25942 8200 26006
rect 8264 25942 8280 26006
rect 8344 25942 8350 26006
rect 7954 25941 8350 25942
rect 4954 25340 5350 25341
rect 4954 25276 4960 25340
rect 5024 25276 5040 25340
rect 5104 25276 5120 25340
rect 5184 25276 5200 25340
rect 5264 25276 5280 25340
rect 5344 25276 5350 25340
rect 4954 25275 5350 25276
rect 0 24672 800 24702
rect 879 24672 945 24675
rect 0 24670 945 24672
rect 0 24614 884 24670
rect 940 24614 945 24670
rect 0 24612 945 24614
rect 0 24582 800 24612
rect 879 24609 945 24612
rect 1954 24674 2350 24675
rect 1954 24610 1960 24674
rect 2024 24610 2040 24674
rect 2104 24610 2120 24674
rect 2184 24610 2200 24674
rect 2264 24610 2280 24674
rect 2344 24610 2350 24674
rect 1954 24609 2350 24610
rect 7954 24674 8350 24675
rect 7954 24610 7960 24674
rect 8024 24610 8040 24674
rect 8104 24610 8120 24674
rect 8184 24610 8200 24674
rect 8264 24610 8280 24674
rect 8344 24610 8350 24674
rect 7954 24609 8350 24610
rect 4954 24008 5350 24009
rect 4954 23944 4960 24008
rect 5024 23944 5040 24008
rect 5104 23944 5120 24008
rect 5184 23944 5200 24008
rect 5264 23944 5280 24008
rect 5344 23944 5350 24008
rect 4954 23943 5350 23944
rect 1954 23342 2350 23343
rect 1954 23278 1960 23342
rect 2024 23278 2040 23342
rect 2104 23278 2120 23342
rect 2184 23278 2200 23342
rect 2264 23278 2280 23342
rect 2344 23278 2350 23342
rect 1954 23277 2350 23278
rect 7954 23342 8350 23343
rect 7954 23278 7960 23342
rect 8024 23278 8040 23342
rect 8104 23278 8120 23342
rect 8184 23278 8200 23342
rect 8264 23278 8280 23342
rect 8344 23278 8350 23342
rect 7954 23277 8350 23278
rect 0 23195 800 23222
rect 0 23190 849 23195
rect 0 23134 788 23190
rect 844 23134 849 23190
rect 0 23129 849 23134
rect 0 23102 800 23129
rect 4954 22676 5350 22677
rect 4954 22612 4960 22676
rect 5024 22612 5040 22676
rect 5104 22612 5120 22676
rect 5184 22612 5200 22676
rect 5264 22612 5280 22676
rect 5344 22612 5350 22676
rect 4954 22611 5350 22612
rect 10095 22600 10161 22603
rect 10922 22600 11722 22630
rect 10095 22598 11722 22600
rect 10095 22542 10100 22598
rect 10156 22542 11722 22598
rect 10095 22540 11722 22542
rect 10095 22537 10161 22540
rect 10922 22510 11722 22540
rect 1954 22010 2350 22011
rect 1954 21946 1960 22010
rect 2024 21946 2040 22010
rect 2104 21946 2120 22010
rect 2184 21946 2200 22010
rect 2264 21946 2280 22010
rect 2344 21946 2350 22010
rect 1954 21945 2350 21946
rect 7954 22010 8350 22011
rect 7954 21946 7960 22010
rect 8024 21946 8040 22010
rect 8104 21946 8120 22010
rect 8184 21946 8200 22010
rect 8264 21946 8280 22010
rect 8344 21946 8350 22010
rect 7954 21945 8350 21946
rect 0 21712 800 21742
rect 879 21712 945 21715
rect 0 21710 945 21712
rect 0 21654 884 21710
rect 940 21654 945 21710
rect 0 21652 945 21654
rect 0 21622 800 21652
rect 879 21649 945 21652
rect 4954 21344 5350 21345
rect 4954 21280 4960 21344
rect 5024 21280 5040 21344
rect 5104 21280 5120 21344
rect 5184 21280 5200 21344
rect 5264 21280 5280 21344
rect 5344 21280 5350 21344
rect 4954 21279 5350 21280
rect 1954 20678 2350 20679
rect 1954 20614 1960 20678
rect 2024 20614 2040 20678
rect 2104 20614 2120 20678
rect 2184 20614 2200 20678
rect 2264 20614 2280 20678
rect 2344 20614 2350 20678
rect 1954 20613 2350 20614
rect 7954 20678 8350 20679
rect 7954 20614 7960 20678
rect 8024 20614 8040 20678
rect 8104 20614 8120 20678
rect 8184 20614 8200 20678
rect 8264 20614 8280 20678
rect 8344 20614 8350 20678
rect 7954 20613 8350 20614
rect 0 20232 800 20262
rect 1551 20232 1617 20235
rect 0 20230 1617 20232
rect 0 20174 1556 20230
rect 1612 20174 1617 20230
rect 0 20172 1617 20174
rect 0 20142 800 20172
rect 1551 20169 1617 20172
rect 10095 20232 10161 20235
rect 10922 20232 11722 20262
rect 10095 20230 11722 20232
rect 10095 20174 10100 20230
rect 10156 20174 11722 20230
rect 10095 20172 11722 20174
rect 10095 20169 10161 20172
rect 10922 20142 11722 20172
rect 4954 20012 5350 20013
rect 4954 19948 4960 20012
rect 5024 19948 5040 20012
rect 5104 19948 5120 20012
rect 5184 19948 5200 20012
rect 5264 19948 5280 20012
rect 5344 19948 5350 20012
rect 4954 19947 5350 19948
rect 1954 19346 2350 19347
rect 1954 19282 1960 19346
rect 2024 19282 2040 19346
rect 2104 19282 2120 19346
rect 2184 19282 2200 19346
rect 2264 19282 2280 19346
rect 2344 19282 2350 19346
rect 1954 19281 2350 19282
rect 7954 19346 8350 19347
rect 7954 19282 7960 19346
rect 8024 19282 8040 19346
rect 8104 19282 8120 19346
rect 8184 19282 8200 19346
rect 8264 19282 8280 19346
rect 8344 19282 8350 19346
rect 7954 19281 8350 19282
rect 0 18752 800 18782
rect 1551 18752 1617 18755
rect 0 18750 1617 18752
rect 0 18694 1556 18750
rect 1612 18694 1617 18750
rect 0 18692 1617 18694
rect 0 18662 800 18692
rect 1551 18689 1617 18692
rect 4954 18680 5350 18681
rect 4954 18616 4960 18680
rect 5024 18616 5040 18680
rect 5104 18616 5120 18680
rect 5184 18616 5200 18680
rect 5264 18616 5280 18680
rect 5344 18616 5350 18680
rect 4954 18615 5350 18616
rect 1954 18014 2350 18015
rect 1954 17950 1960 18014
rect 2024 17950 2040 18014
rect 2104 17950 2120 18014
rect 2184 17950 2200 18014
rect 2264 17950 2280 18014
rect 2344 17950 2350 18014
rect 1954 17949 2350 17950
rect 7954 18014 8350 18015
rect 7954 17950 7960 18014
rect 8024 17950 8040 18014
rect 8104 17950 8120 18014
rect 8184 17950 8200 18014
rect 8264 17950 8280 18014
rect 8344 17950 8350 18014
rect 7954 17949 8350 17950
rect 10095 17864 10161 17867
rect 10922 17864 11722 17894
rect 10095 17862 11722 17864
rect 10095 17806 10100 17862
rect 10156 17806 11722 17862
rect 10095 17804 11722 17806
rect 10095 17801 10161 17804
rect 10922 17774 11722 17804
rect 4954 17348 5350 17349
rect 0 17272 800 17302
rect 4954 17284 4960 17348
rect 5024 17284 5040 17348
rect 5104 17284 5120 17348
rect 5184 17284 5200 17348
rect 5264 17284 5280 17348
rect 5344 17284 5350 17348
rect 4954 17283 5350 17284
rect 1263 17272 1329 17275
rect 0 17270 1329 17272
rect 0 17214 1268 17270
rect 1324 17214 1329 17270
rect 0 17212 1329 17214
rect 0 17182 800 17212
rect 1263 17209 1329 17212
rect 1954 16682 2350 16683
rect 1954 16618 1960 16682
rect 2024 16618 2040 16682
rect 2104 16618 2120 16682
rect 2184 16618 2200 16682
rect 2264 16618 2280 16682
rect 2344 16618 2350 16682
rect 1954 16617 2350 16618
rect 7954 16682 8350 16683
rect 7954 16618 7960 16682
rect 8024 16618 8040 16682
rect 8104 16618 8120 16682
rect 8184 16618 8200 16682
rect 8264 16618 8280 16682
rect 8344 16618 8350 16682
rect 7954 16617 8350 16618
rect 4954 16016 5350 16017
rect 4954 15952 4960 16016
rect 5024 15952 5040 16016
rect 5104 15952 5120 16016
rect 5184 15952 5200 16016
rect 5264 15952 5280 16016
rect 5344 15952 5350 16016
rect 4954 15951 5350 15952
rect 0 15795 800 15822
rect 0 15790 849 15795
rect 0 15734 788 15790
rect 844 15734 849 15790
rect 0 15729 849 15734
rect 0 15702 800 15729
rect 10095 15496 10161 15499
rect 10922 15496 11722 15526
rect 10095 15494 11722 15496
rect 10095 15438 10100 15494
rect 10156 15438 11722 15494
rect 10095 15436 11722 15438
rect 10095 15433 10161 15436
rect 10922 15406 11722 15436
rect 1954 15350 2350 15351
rect 1954 15286 1960 15350
rect 2024 15286 2040 15350
rect 2104 15286 2120 15350
rect 2184 15286 2200 15350
rect 2264 15286 2280 15350
rect 2344 15286 2350 15350
rect 1954 15285 2350 15286
rect 7954 15350 8350 15351
rect 7954 15286 7960 15350
rect 8024 15286 8040 15350
rect 8104 15286 8120 15350
rect 8184 15286 8200 15350
rect 8264 15286 8280 15350
rect 8344 15286 8350 15350
rect 7954 15285 8350 15286
rect 4954 14684 5350 14685
rect 4954 14620 4960 14684
rect 5024 14620 5040 14684
rect 5104 14620 5120 14684
rect 5184 14620 5200 14684
rect 5264 14620 5280 14684
rect 5344 14620 5350 14684
rect 4954 14619 5350 14620
rect 0 14315 800 14342
rect 0 14310 849 14315
rect 0 14254 788 14310
rect 844 14254 849 14310
rect 0 14249 849 14254
rect 0 14222 800 14249
rect 1954 14018 2350 14019
rect 1954 13954 1960 14018
rect 2024 13954 2040 14018
rect 2104 13954 2120 14018
rect 2184 13954 2200 14018
rect 2264 13954 2280 14018
rect 2344 13954 2350 14018
rect 1954 13953 2350 13954
rect 7954 14018 8350 14019
rect 7954 13954 7960 14018
rect 8024 13954 8040 14018
rect 8104 13954 8120 14018
rect 8184 13954 8200 14018
rect 8264 13954 8280 14018
rect 8344 13954 8350 14018
rect 7954 13953 8350 13954
rect 4954 13352 5350 13353
rect 4954 13288 4960 13352
rect 5024 13288 5040 13352
rect 5104 13288 5120 13352
rect 5184 13288 5200 13352
rect 5264 13288 5280 13352
rect 5344 13288 5350 13352
rect 4954 13287 5350 13288
rect 10095 13128 10161 13131
rect 10922 13128 11722 13158
rect 10095 13126 11722 13128
rect 10095 13070 10100 13126
rect 10156 13070 11722 13126
rect 10095 13068 11722 13070
rect 10095 13065 10161 13068
rect 10922 13038 11722 13068
rect 0 12832 800 12862
rect 1551 12832 1617 12835
rect 0 12830 1617 12832
rect 0 12774 1556 12830
rect 1612 12774 1617 12830
rect 0 12772 1617 12774
rect 0 12742 800 12772
rect 1551 12769 1617 12772
rect 1954 12686 2350 12687
rect 1954 12622 1960 12686
rect 2024 12622 2040 12686
rect 2104 12622 2120 12686
rect 2184 12622 2200 12686
rect 2264 12622 2280 12686
rect 2344 12622 2350 12686
rect 1954 12621 2350 12622
rect 7954 12686 8350 12687
rect 7954 12622 7960 12686
rect 8024 12622 8040 12686
rect 8104 12622 8120 12686
rect 8184 12622 8200 12686
rect 8264 12622 8280 12686
rect 8344 12622 8350 12686
rect 7954 12621 8350 12622
rect 4954 12020 5350 12021
rect 4954 11956 4960 12020
rect 5024 11956 5040 12020
rect 5104 11956 5120 12020
rect 5184 11956 5200 12020
rect 5264 11956 5280 12020
rect 5344 11956 5350 12020
rect 4954 11955 5350 11956
rect 0 11352 800 11382
rect 1551 11352 1617 11355
rect 0 11350 1617 11352
rect 0 11294 1556 11350
rect 1612 11294 1617 11350
rect 0 11292 1617 11294
rect 0 11262 800 11292
rect 1551 11289 1617 11292
rect 1954 11354 2350 11355
rect 1954 11290 1960 11354
rect 2024 11290 2040 11354
rect 2104 11290 2120 11354
rect 2184 11290 2200 11354
rect 2264 11290 2280 11354
rect 2344 11290 2350 11354
rect 1954 11289 2350 11290
rect 7954 11354 8350 11355
rect 7954 11290 7960 11354
rect 8024 11290 8040 11354
rect 8104 11290 8120 11354
rect 8184 11290 8200 11354
rect 8264 11290 8280 11354
rect 8344 11290 8350 11354
rect 7954 11289 8350 11290
rect 10095 10760 10161 10763
rect 10922 10760 11722 10790
rect 10095 10758 11722 10760
rect 10095 10702 10100 10758
rect 10156 10702 11722 10758
rect 10095 10700 11722 10702
rect 10095 10697 10161 10700
rect 4954 10688 5350 10689
rect 4954 10624 4960 10688
rect 5024 10624 5040 10688
rect 5104 10624 5120 10688
rect 5184 10624 5200 10688
rect 5264 10624 5280 10688
rect 5344 10624 5350 10688
rect 10922 10670 11722 10700
rect 4954 10623 5350 10624
rect 1954 10022 2350 10023
rect 1954 9958 1960 10022
rect 2024 9958 2040 10022
rect 2104 9958 2120 10022
rect 2184 9958 2200 10022
rect 2264 9958 2280 10022
rect 2344 9958 2350 10022
rect 1954 9957 2350 9958
rect 7954 10022 8350 10023
rect 7954 9958 7960 10022
rect 8024 9958 8040 10022
rect 8104 9958 8120 10022
rect 8184 9958 8200 10022
rect 8264 9958 8280 10022
rect 8344 9958 8350 10022
rect 7954 9957 8350 9958
rect 0 9872 800 9902
rect 1551 9872 1617 9875
rect 0 9870 1617 9872
rect 0 9814 1556 9870
rect 1612 9814 1617 9870
rect 0 9812 1617 9814
rect 0 9782 800 9812
rect 1551 9809 1617 9812
rect 4954 9356 5350 9357
rect 4954 9292 4960 9356
rect 5024 9292 5040 9356
rect 5104 9292 5120 9356
rect 5184 9292 5200 9356
rect 5264 9292 5280 9356
rect 5344 9292 5350 9356
rect 4954 9291 5350 9292
rect 1954 8690 2350 8691
rect 1954 8626 1960 8690
rect 2024 8626 2040 8690
rect 2104 8626 2120 8690
rect 2184 8626 2200 8690
rect 2264 8626 2280 8690
rect 2344 8626 2350 8690
rect 1954 8625 2350 8626
rect 7954 8690 8350 8691
rect 7954 8626 7960 8690
rect 8024 8626 8040 8690
rect 8104 8626 8120 8690
rect 8184 8626 8200 8690
rect 8264 8626 8280 8690
rect 8344 8626 8350 8690
rect 7954 8625 8350 8626
rect 0 8392 800 8422
rect 1647 8392 1713 8395
rect 0 8390 1713 8392
rect 0 8334 1652 8390
rect 1708 8334 1713 8390
rect 0 8332 1713 8334
rect 0 8302 800 8332
rect 1647 8329 1713 8332
rect 10095 8392 10161 8395
rect 10922 8392 11722 8422
rect 10095 8390 11722 8392
rect 10095 8334 10100 8390
rect 10156 8334 11722 8390
rect 10095 8332 11722 8334
rect 10095 8329 10161 8332
rect 10922 8302 11722 8332
rect 4954 8024 5350 8025
rect 4954 7960 4960 8024
rect 5024 7960 5040 8024
rect 5104 7960 5120 8024
rect 5184 7960 5200 8024
rect 5264 7960 5280 8024
rect 5344 7960 5350 8024
rect 4954 7959 5350 7960
rect 1954 7358 2350 7359
rect 1954 7294 1960 7358
rect 2024 7294 2040 7358
rect 2104 7294 2120 7358
rect 2184 7294 2200 7358
rect 2264 7294 2280 7358
rect 2344 7294 2350 7358
rect 1954 7293 2350 7294
rect 7954 7358 8350 7359
rect 7954 7294 7960 7358
rect 8024 7294 8040 7358
rect 8104 7294 8120 7358
rect 8184 7294 8200 7358
rect 8264 7294 8280 7358
rect 8344 7294 8350 7358
rect 7954 7293 8350 7294
rect 0 6912 800 6942
rect 1647 6912 1713 6915
rect 0 6910 1713 6912
rect 0 6854 1652 6910
rect 1708 6854 1713 6910
rect 0 6852 1713 6854
rect 0 6822 800 6852
rect 1647 6849 1713 6852
rect 4954 6692 5350 6693
rect 4954 6628 4960 6692
rect 5024 6628 5040 6692
rect 5104 6628 5120 6692
rect 5184 6628 5200 6692
rect 5264 6628 5280 6692
rect 5344 6628 5350 6692
rect 4954 6627 5350 6628
rect 1954 6026 2350 6027
rect 1954 5962 1960 6026
rect 2024 5962 2040 6026
rect 2104 5962 2120 6026
rect 2184 5962 2200 6026
rect 2264 5962 2280 6026
rect 2344 5962 2350 6026
rect 1954 5961 2350 5962
rect 7954 6026 8350 6027
rect 7954 5962 7960 6026
rect 8024 5962 8040 6026
rect 8104 5962 8120 6026
rect 8184 5962 8200 6026
rect 8264 5962 8280 6026
rect 8344 5962 8350 6026
rect 7954 5961 8350 5962
rect 10095 6024 10161 6027
rect 10922 6024 11722 6054
rect 10095 6022 11722 6024
rect 10095 5966 10100 6022
rect 10156 5966 11722 6022
rect 10095 5964 11722 5966
rect 10095 5961 10161 5964
rect 10922 5934 11722 5964
rect 6351 5580 6417 5583
rect 3138 5578 6417 5580
rect 3138 5522 6356 5578
rect 6412 5522 6417 5578
rect 3138 5520 6417 5522
rect 0 5432 800 5462
rect 3138 5432 3198 5520
rect 6351 5517 6417 5520
rect 0 5372 3198 5432
rect 0 5342 800 5372
rect 4954 5360 5350 5361
rect 4954 5296 4960 5360
rect 5024 5296 5040 5360
rect 5104 5296 5120 5360
rect 5184 5296 5200 5360
rect 5264 5296 5280 5360
rect 5344 5296 5350 5360
rect 4954 5295 5350 5296
rect 1954 4694 2350 4695
rect 1954 4630 1960 4694
rect 2024 4630 2040 4694
rect 2104 4630 2120 4694
rect 2184 4630 2200 4694
rect 2264 4630 2280 4694
rect 2344 4630 2350 4694
rect 1954 4629 2350 4630
rect 7954 4694 8350 4695
rect 7954 4630 7960 4694
rect 8024 4630 8040 4694
rect 8104 4630 8120 4694
rect 8184 4630 8200 4694
rect 8264 4630 8280 4694
rect 8344 4630 8350 4694
rect 7954 4629 8350 4630
rect 4954 4028 5350 4029
rect 0 3952 800 3982
rect 4954 3964 4960 4028
rect 5024 3964 5040 4028
rect 5104 3964 5120 4028
rect 5184 3964 5200 4028
rect 5264 3964 5280 4028
rect 5344 3964 5350 4028
rect 4954 3963 5350 3964
rect 879 3952 945 3955
rect 0 3950 945 3952
rect 0 3894 884 3950
rect 940 3894 945 3950
rect 0 3892 945 3894
rect 0 3862 800 3892
rect 879 3889 945 3892
rect 10095 3656 10161 3659
rect 10922 3656 11722 3686
rect 10095 3654 11722 3656
rect 10095 3598 10100 3654
rect 10156 3598 11722 3654
rect 10095 3596 11722 3598
rect 10095 3593 10161 3596
rect 10922 3566 11722 3596
rect 1954 3362 2350 3363
rect 1954 3298 1960 3362
rect 2024 3298 2040 3362
rect 2104 3298 2120 3362
rect 2184 3298 2200 3362
rect 2264 3298 2280 3362
rect 2344 3298 2350 3362
rect 1954 3297 2350 3298
rect 7954 3362 8350 3363
rect 7954 3298 7960 3362
rect 8024 3298 8040 3362
rect 8104 3298 8120 3362
rect 8184 3298 8200 3362
rect 8264 3298 8280 3362
rect 8344 3298 8350 3362
rect 7954 3297 8350 3298
rect 4954 2696 5350 2697
rect 4954 2632 4960 2696
rect 5024 2632 5040 2696
rect 5104 2632 5120 2696
rect 5184 2632 5200 2696
rect 5264 2632 5280 2696
rect 5344 2632 5350 2696
rect 4954 2631 5350 2632
rect 0 2472 800 2502
rect 2223 2472 2289 2475
rect 0 2470 2289 2472
rect 0 2414 2228 2470
rect 2284 2414 2289 2470
rect 0 2412 2289 2414
rect 0 2382 800 2412
rect 2223 2409 2289 2412
rect 9711 1288 9777 1291
rect 10922 1288 11722 1318
rect 9711 1286 11722 1288
rect 9711 1230 9716 1286
rect 9772 1230 11722 1286
rect 9711 1228 11722 1230
rect 9711 1225 9777 1228
rect 10922 1198 11722 1228
<< via3 >>
rect 1960 26002 2024 26006
rect 1960 25946 1964 26002
rect 1964 25946 2020 26002
rect 2020 25946 2024 26002
rect 1960 25942 2024 25946
rect 2040 26002 2104 26006
rect 2040 25946 2044 26002
rect 2044 25946 2100 26002
rect 2100 25946 2104 26002
rect 2040 25942 2104 25946
rect 2120 26002 2184 26006
rect 2120 25946 2124 26002
rect 2124 25946 2180 26002
rect 2180 25946 2184 26002
rect 2120 25942 2184 25946
rect 2200 26002 2264 26006
rect 2200 25946 2204 26002
rect 2204 25946 2260 26002
rect 2260 25946 2264 26002
rect 2200 25942 2264 25946
rect 2280 26002 2344 26006
rect 2280 25946 2284 26002
rect 2284 25946 2340 26002
rect 2340 25946 2344 26002
rect 2280 25942 2344 25946
rect 7960 26002 8024 26006
rect 7960 25946 7964 26002
rect 7964 25946 8020 26002
rect 8020 25946 8024 26002
rect 7960 25942 8024 25946
rect 8040 26002 8104 26006
rect 8040 25946 8044 26002
rect 8044 25946 8100 26002
rect 8100 25946 8104 26002
rect 8040 25942 8104 25946
rect 8120 26002 8184 26006
rect 8120 25946 8124 26002
rect 8124 25946 8180 26002
rect 8180 25946 8184 26002
rect 8120 25942 8184 25946
rect 8200 26002 8264 26006
rect 8200 25946 8204 26002
rect 8204 25946 8260 26002
rect 8260 25946 8264 26002
rect 8200 25942 8264 25946
rect 8280 26002 8344 26006
rect 8280 25946 8284 26002
rect 8284 25946 8340 26002
rect 8340 25946 8344 26002
rect 8280 25942 8344 25946
rect 4960 25336 5024 25340
rect 4960 25280 4964 25336
rect 4964 25280 5020 25336
rect 5020 25280 5024 25336
rect 4960 25276 5024 25280
rect 5040 25336 5104 25340
rect 5040 25280 5044 25336
rect 5044 25280 5100 25336
rect 5100 25280 5104 25336
rect 5040 25276 5104 25280
rect 5120 25336 5184 25340
rect 5120 25280 5124 25336
rect 5124 25280 5180 25336
rect 5180 25280 5184 25336
rect 5120 25276 5184 25280
rect 5200 25336 5264 25340
rect 5200 25280 5204 25336
rect 5204 25280 5260 25336
rect 5260 25280 5264 25336
rect 5200 25276 5264 25280
rect 5280 25336 5344 25340
rect 5280 25280 5284 25336
rect 5284 25280 5340 25336
rect 5340 25280 5344 25336
rect 5280 25276 5344 25280
rect 1960 24670 2024 24674
rect 1960 24614 1964 24670
rect 1964 24614 2020 24670
rect 2020 24614 2024 24670
rect 1960 24610 2024 24614
rect 2040 24670 2104 24674
rect 2040 24614 2044 24670
rect 2044 24614 2100 24670
rect 2100 24614 2104 24670
rect 2040 24610 2104 24614
rect 2120 24670 2184 24674
rect 2120 24614 2124 24670
rect 2124 24614 2180 24670
rect 2180 24614 2184 24670
rect 2120 24610 2184 24614
rect 2200 24670 2264 24674
rect 2200 24614 2204 24670
rect 2204 24614 2260 24670
rect 2260 24614 2264 24670
rect 2200 24610 2264 24614
rect 2280 24670 2344 24674
rect 2280 24614 2284 24670
rect 2284 24614 2340 24670
rect 2340 24614 2344 24670
rect 2280 24610 2344 24614
rect 7960 24670 8024 24674
rect 7960 24614 7964 24670
rect 7964 24614 8020 24670
rect 8020 24614 8024 24670
rect 7960 24610 8024 24614
rect 8040 24670 8104 24674
rect 8040 24614 8044 24670
rect 8044 24614 8100 24670
rect 8100 24614 8104 24670
rect 8040 24610 8104 24614
rect 8120 24670 8184 24674
rect 8120 24614 8124 24670
rect 8124 24614 8180 24670
rect 8180 24614 8184 24670
rect 8120 24610 8184 24614
rect 8200 24670 8264 24674
rect 8200 24614 8204 24670
rect 8204 24614 8260 24670
rect 8260 24614 8264 24670
rect 8200 24610 8264 24614
rect 8280 24670 8344 24674
rect 8280 24614 8284 24670
rect 8284 24614 8340 24670
rect 8340 24614 8344 24670
rect 8280 24610 8344 24614
rect 4960 24004 5024 24008
rect 4960 23948 4964 24004
rect 4964 23948 5020 24004
rect 5020 23948 5024 24004
rect 4960 23944 5024 23948
rect 5040 24004 5104 24008
rect 5040 23948 5044 24004
rect 5044 23948 5100 24004
rect 5100 23948 5104 24004
rect 5040 23944 5104 23948
rect 5120 24004 5184 24008
rect 5120 23948 5124 24004
rect 5124 23948 5180 24004
rect 5180 23948 5184 24004
rect 5120 23944 5184 23948
rect 5200 24004 5264 24008
rect 5200 23948 5204 24004
rect 5204 23948 5260 24004
rect 5260 23948 5264 24004
rect 5200 23944 5264 23948
rect 5280 24004 5344 24008
rect 5280 23948 5284 24004
rect 5284 23948 5340 24004
rect 5340 23948 5344 24004
rect 5280 23944 5344 23948
rect 1960 23338 2024 23342
rect 1960 23282 1964 23338
rect 1964 23282 2020 23338
rect 2020 23282 2024 23338
rect 1960 23278 2024 23282
rect 2040 23338 2104 23342
rect 2040 23282 2044 23338
rect 2044 23282 2100 23338
rect 2100 23282 2104 23338
rect 2040 23278 2104 23282
rect 2120 23338 2184 23342
rect 2120 23282 2124 23338
rect 2124 23282 2180 23338
rect 2180 23282 2184 23338
rect 2120 23278 2184 23282
rect 2200 23338 2264 23342
rect 2200 23282 2204 23338
rect 2204 23282 2260 23338
rect 2260 23282 2264 23338
rect 2200 23278 2264 23282
rect 2280 23338 2344 23342
rect 2280 23282 2284 23338
rect 2284 23282 2340 23338
rect 2340 23282 2344 23338
rect 2280 23278 2344 23282
rect 7960 23338 8024 23342
rect 7960 23282 7964 23338
rect 7964 23282 8020 23338
rect 8020 23282 8024 23338
rect 7960 23278 8024 23282
rect 8040 23338 8104 23342
rect 8040 23282 8044 23338
rect 8044 23282 8100 23338
rect 8100 23282 8104 23338
rect 8040 23278 8104 23282
rect 8120 23338 8184 23342
rect 8120 23282 8124 23338
rect 8124 23282 8180 23338
rect 8180 23282 8184 23338
rect 8120 23278 8184 23282
rect 8200 23338 8264 23342
rect 8200 23282 8204 23338
rect 8204 23282 8260 23338
rect 8260 23282 8264 23338
rect 8200 23278 8264 23282
rect 8280 23338 8344 23342
rect 8280 23282 8284 23338
rect 8284 23282 8340 23338
rect 8340 23282 8344 23338
rect 8280 23278 8344 23282
rect 4960 22672 5024 22676
rect 4960 22616 4964 22672
rect 4964 22616 5020 22672
rect 5020 22616 5024 22672
rect 4960 22612 5024 22616
rect 5040 22672 5104 22676
rect 5040 22616 5044 22672
rect 5044 22616 5100 22672
rect 5100 22616 5104 22672
rect 5040 22612 5104 22616
rect 5120 22672 5184 22676
rect 5120 22616 5124 22672
rect 5124 22616 5180 22672
rect 5180 22616 5184 22672
rect 5120 22612 5184 22616
rect 5200 22672 5264 22676
rect 5200 22616 5204 22672
rect 5204 22616 5260 22672
rect 5260 22616 5264 22672
rect 5200 22612 5264 22616
rect 5280 22672 5344 22676
rect 5280 22616 5284 22672
rect 5284 22616 5340 22672
rect 5340 22616 5344 22672
rect 5280 22612 5344 22616
rect 1960 22006 2024 22010
rect 1960 21950 1964 22006
rect 1964 21950 2020 22006
rect 2020 21950 2024 22006
rect 1960 21946 2024 21950
rect 2040 22006 2104 22010
rect 2040 21950 2044 22006
rect 2044 21950 2100 22006
rect 2100 21950 2104 22006
rect 2040 21946 2104 21950
rect 2120 22006 2184 22010
rect 2120 21950 2124 22006
rect 2124 21950 2180 22006
rect 2180 21950 2184 22006
rect 2120 21946 2184 21950
rect 2200 22006 2264 22010
rect 2200 21950 2204 22006
rect 2204 21950 2260 22006
rect 2260 21950 2264 22006
rect 2200 21946 2264 21950
rect 2280 22006 2344 22010
rect 2280 21950 2284 22006
rect 2284 21950 2340 22006
rect 2340 21950 2344 22006
rect 2280 21946 2344 21950
rect 7960 22006 8024 22010
rect 7960 21950 7964 22006
rect 7964 21950 8020 22006
rect 8020 21950 8024 22006
rect 7960 21946 8024 21950
rect 8040 22006 8104 22010
rect 8040 21950 8044 22006
rect 8044 21950 8100 22006
rect 8100 21950 8104 22006
rect 8040 21946 8104 21950
rect 8120 22006 8184 22010
rect 8120 21950 8124 22006
rect 8124 21950 8180 22006
rect 8180 21950 8184 22006
rect 8120 21946 8184 21950
rect 8200 22006 8264 22010
rect 8200 21950 8204 22006
rect 8204 21950 8260 22006
rect 8260 21950 8264 22006
rect 8200 21946 8264 21950
rect 8280 22006 8344 22010
rect 8280 21950 8284 22006
rect 8284 21950 8340 22006
rect 8340 21950 8344 22006
rect 8280 21946 8344 21950
rect 4960 21340 5024 21344
rect 4960 21284 4964 21340
rect 4964 21284 5020 21340
rect 5020 21284 5024 21340
rect 4960 21280 5024 21284
rect 5040 21340 5104 21344
rect 5040 21284 5044 21340
rect 5044 21284 5100 21340
rect 5100 21284 5104 21340
rect 5040 21280 5104 21284
rect 5120 21340 5184 21344
rect 5120 21284 5124 21340
rect 5124 21284 5180 21340
rect 5180 21284 5184 21340
rect 5120 21280 5184 21284
rect 5200 21340 5264 21344
rect 5200 21284 5204 21340
rect 5204 21284 5260 21340
rect 5260 21284 5264 21340
rect 5200 21280 5264 21284
rect 5280 21340 5344 21344
rect 5280 21284 5284 21340
rect 5284 21284 5340 21340
rect 5340 21284 5344 21340
rect 5280 21280 5344 21284
rect 1960 20674 2024 20678
rect 1960 20618 1964 20674
rect 1964 20618 2020 20674
rect 2020 20618 2024 20674
rect 1960 20614 2024 20618
rect 2040 20674 2104 20678
rect 2040 20618 2044 20674
rect 2044 20618 2100 20674
rect 2100 20618 2104 20674
rect 2040 20614 2104 20618
rect 2120 20674 2184 20678
rect 2120 20618 2124 20674
rect 2124 20618 2180 20674
rect 2180 20618 2184 20674
rect 2120 20614 2184 20618
rect 2200 20674 2264 20678
rect 2200 20618 2204 20674
rect 2204 20618 2260 20674
rect 2260 20618 2264 20674
rect 2200 20614 2264 20618
rect 2280 20674 2344 20678
rect 2280 20618 2284 20674
rect 2284 20618 2340 20674
rect 2340 20618 2344 20674
rect 2280 20614 2344 20618
rect 7960 20674 8024 20678
rect 7960 20618 7964 20674
rect 7964 20618 8020 20674
rect 8020 20618 8024 20674
rect 7960 20614 8024 20618
rect 8040 20674 8104 20678
rect 8040 20618 8044 20674
rect 8044 20618 8100 20674
rect 8100 20618 8104 20674
rect 8040 20614 8104 20618
rect 8120 20674 8184 20678
rect 8120 20618 8124 20674
rect 8124 20618 8180 20674
rect 8180 20618 8184 20674
rect 8120 20614 8184 20618
rect 8200 20674 8264 20678
rect 8200 20618 8204 20674
rect 8204 20618 8260 20674
rect 8260 20618 8264 20674
rect 8200 20614 8264 20618
rect 8280 20674 8344 20678
rect 8280 20618 8284 20674
rect 8284 20618 8340 20674
rect 8340 20618 8344 20674
rect 8280 20614 8344 20618
rect 4960 20008 5024 20012
rect 4960 19952 4964 20008
rect 4964 19952 5020 20008
rect 5020 19952 5024 20008
rect 4960 19948 5024 19952
rect 5040 20008 5104 20012
rect 5040 19952 5044 20008
rect 5044 19952 5100 20008
rect 5100 19952 5104 20008
rect 5040 19948 5104 19952
rect 5120 20008 5184 20012
rect 5120 19952 5124 20008
rect 5124 19952 5180 20008
rect 5180 19952 5184 20008
rect 5120 19948 5184 19952
rect 5200 20008 5264 20012
rect 5200 19952 5204 20008
rect 5204 19952 5260 20008
rect 5260 19952 5264 20008
rect 5200 19948 5264 19952
rect 5280 20008 5344 20012
rect 5280 19952 5284 20008
rect 5284 19952 5340 20008
rect 5340 19952 5344 20008
rect 5280 19948 5344 19952
rect 1960 19342 2024 19346
rect 1960 19286 1964 19342
rect 1964 19286 2020 19342
rect 2020 19286 2024 19342
rect 1960 19282 2024 19286
rect 2040 19342 2104 19346
rect 2040 19286 2044 19342
rect 2044 19286 2100 19342
rect 2100 19286 2104 19342
rect 2040 19282 2104 19286
rect 2120 19342 2184 19346
rect 2120 19286 2124 19342
rect 2124 19286 2180 19342
rect 2180 19286 2184 19342
rect 2120 19282 2184 19286
rect 2200 19342 2264 19346
rect 2200 19286 2204 19342
rect 2204 19286 2260 19342
rect 2260 19286 2264 19342
rect 2200 19282 2264 19286
rect 2280 19342 2344 19346
rect 2280 19286 2284 19342
rect 2284 19286 2340 19342
rect 2340 19286 2344 19342
rect 2280 19282 2344 19286
rect 7960 19342 8024 19346
rect 7960 19286 7964 19342
rect 7964 19286 8020 19342
rect 8020 19286 8024 19342
rect 7960 19282 8024 19286
rect 8040 19342 8104 19346
rect 8040 19286 8044 19342
rect 8044 19286 8100 19342
rect 8100 19286 8104 19342
rect 8040 19282 8104 19286
rect 8120 19342 8184 19346
rect 8120 19286 8124 19342
rect 8124 19286 8180 19342
rect 8180 19286 8184 19342
rect 8120 19282 8184 19286
rect 8200 19342 8264 19346
rect 8200 19286 8204 19342
rect 8204 19286 8260 19342
rect 8260 19286 8264 19342
rect 8200 19282 8264 19286
rect 8280 19342 8344 19346
rect 8280 19286 8284 19342
rect 8284 19286 8340 19342
rect 8340 19286 8344 19342
rect 8280 19282 8344 19286
rect 4960 18676 5024 18680
rect 4960 18620 4964 18676
rect 4964 18620 5020 18676
rect 5020 18620 5024 18676
rect 4960 18616 5024 18620
rect 5040 18676 5104 18680
rect 5040 18620 5044 18676
rect 5044 18620 5100 18676
rect 5100 18620 5104 18676
rect 5040 18616 5104 18620
rect 5120 18676 5184 18680
rect 5120 18620 5124 18676
rect 5124 18620 5180 18676
rect 5180 18620 5184 18676
rect 5120 18616 5184 18620
rect 5200 18676 5264 18680
rect 5200 18620 5204 18676
rect 5204 18620 5260 18676
rect 5260 18620 5264 18676
rect 5200 18616 5264 18620
rect 5280 18676 5344 18680
rect 5280 18620 5284 18676
rect 5284 18620 5340 18676
rect 5340 18620 5344 18676
rect 5280 18616 5344 18620
rect 1960 18010 2024 18014
rect 1960 17954 1964 18010
rect 1964 17954 2020 18010
rect 2020 17954 2024 18010
rect 1960 17950 2024 17954
rect 2040 18010 2104 18014
rect 2040 17954 2044 18010
rect 2044 17954 2100 18010
rect 2100 17954 2104 18010
rect 2040 17950 2104 17954
rect 2120 18010 2184 18014
rect 2120 17954 2124 18010
rect 2124 17954 2180 18010
rect 2180 17954 2184 18010
rect 2120 17950 2184 17954
rect 2200 18010 2264 18014
rect 2200 17954 2204 18010
rect 2204 17954 2260 18010
rect 2260 17954 2264 18010
rect 2200 17950 2264 17954
rect 2280 18010 2344 18014
rect 2280 17954 2284 18010
rect 2284 17954 2340 18010
rect 2340 17954 2344 18010
rect 2280 17950 2344 17954
rect 7960 18010 8024 18014
rect 7960 17954 7964 18010
rect 7964 17954 8020 18010
rect 8020 17954 8024 18010
rect 7960 17950 8024 17954
rect 8040 18010 8104 18014
rect 8040 17954 8044 18010
rect 8044 17954 8100 18010
rect 8100 17954 8104 18010
rect 8040 17950 8104 17954
rect 8120 18010 8184 18014
rect 8120 17954 8124 18010
rect 8124 17954 8180 18010
rect 8180 17954 8184 18010
rect 8120 17950 8184 17954
rect 8200 18010 8264 18014
rect 8200 17954 8204 18010
rect 8204 17954 8260 18010
rect 8260 17954 8264 18010
rect 8200 17950 8264 17954
rect 8280 18010 8344 18014
rect 8280 17954 8284 18010
rect 8284 17954 8340 18010
rect 8340 17954 8344 18010
rect 8280 17950 8344 17954
rect 4960 17344 5024 17348
rect 4960 17288 4964 17344
rect 4964 17288 5020 17344
rect 5020 17288 5024 17344
rect 4960 17284 5024 17288
rect 5040 17344 5104 17348
rect 5040 17288 5044 17344
rect 5044 17288 5100 17344
rect 5100 17288 5104 17344
rect 5040 17284 5104 17288
rect 5120 17344 5184 17348
rect 5120 17288 5124 17344
rect 5124 17288 5180 17344
rect 5180 17288 5184 17344
rect 5120 17284 5184 17288
rect 5200 17344 5264 17348
rect 5200 17288 5204 17344
rect 5204 17288 5260 17344
rect 5260 17288 5264 17344
rect 5200 17284 5264 17288
rect 5280 17344 5344 17348
rect 5280 17288 5284 17344
rect 5284 17288 5340 17344
rect 5340 17288 5344 17344
rect 5280 17284 5344 17288
rect 1960 16678 2024 16682
rect 1960 16622 1964 16678
rect 1964 16622 2020 16678
rect 2020 16622 2024 16678
rect 1960 16618 2024 16622
rect 2040 16678 2104 16682
rect 2040 16622 2044 16678
rect 2044 16622 2100 16678
rect 2100 16622 2104 16678
rect 2040 16618 2104 16622
rect 2120 16678 2184 16682
rect 2120 16622 2124 16678
rect 2124 16622 2180 16678
rect 2180 16622 2184 16678
rect 2120 16618 2184 16622
rect 2200 16678 2264 16682
rect 2200 16622 2204 16678
rect 2204 16622 2260 16678
rect 2260 16622 2264 16678
rect 2200 16618 2264 16622
rect 2280 16678 2344 16682
rect 2280 16622 2284 16678
rect 2284 16622 2340 16678
rect 2340 16622 2344 16678
rect 2280 16618 2344 16622
rect 7960 16678 8024 16682
rect 7960 16622 7964 16678
rect 7964 16622 8020 16678
rect 8020 16622 8024 16678
rect 7960 16618 8024 16622
rect 8040 16678 8104 16682
rect 8040 16622 8044 16678
rect 8044 16622 8100 16678
rect 8100 16622 8104 16678
rect 8040 16618 8104 16622
rect 8120 16678 8184 16682
rect 8120 16622 8124 16678
rect 8124 16622 8180 16678
rect 8180 16622 8184 16678
rect 8120 16618 8184 16622
rect 8200 16678 8264 16682
rect 8200 16622 8204 16678
rect 8204 16622 8260 16678
rect 8260 16622 8264 16678
rect 8200 16618 8264 16622
rect 8280 16678 8344 16682
rect 8280 16622 8284 16678
rect 8284 16622 8340 16678
rect 8340 16622 8344 16678
rect 8280 16618 8344 16622
rect 4960 16012 5024 16016
rect 4960 15956 4964 16012
rect 4964 15956 5020 16012
rect 5020 15956 5024 16012
rect 4960 15952 5024 15956
rect 5040 16012 5104 16016
rect 5040 15956 5044 16012
rect 5044 15956 5100 16012
rect 5100 15956 5104 16012
rect 5040 15952 5104 15956
rect 5120 16012 5184 16016
rect 5120 15956 5124 16012
rect 5124 15956 5180 16012
rect 5180 15956 5184 16012
rect 5120 15952 5184 15956
rect 5200 16012 5264 16016
rect 5200 15956 5204 16012
rect 5204 15956 5260 16012
rect 5260 15956 5264 16012
rect 5200 15952 5264 15956
rect 5280 16012 5344 16016
rect 5280 15956 5284 16012
rect 5284 15956 5340 16012
rect 5340 15956 5344 16012
rect 5280 15952 5344 15956
rect 1960 15346 2024 15350
rect 1960 15290 1964 15346
rect 1964 15290 2020 15346
rect 2020 15290 2024 15346
rect 1960 15286 2024 15290
rect 2040 15346 2104 15350
rect 2040 15290 2044 15346
rect 2044 15290 2100 15346
rect 2100 15290 2104 15346
rect 2040 15286 2104 15290
rect 2120 15346 2184 15350
rect 2120 15290 2124 15346
rect 2124 15290 2180 15346
rect 2180 15290 2184 15346
rect 2120 15286 2184 15290
rect 2200 15346 2264 15350
rect 2200 15290 2204 15346
rect 2204 15290 2260 15346
rect 2260 15290 2264 15346
rect 2200 15286 2264 15290
rect 2280 15346 2344 15350
rect 2280 15290 2284 15346
rect 2284 15290 2340 15346
rect 2340 15290 2344 15346
rect 2280 15286 2344 15290
rect 7960 15346 8024 15350
rect 7960 15290 7964 15346
rect 7964 15290 8020 15346
rect 8020 15290 8024 15346
rect 7960 15286 8024 15290
rect 8040 15346 8104 15350
rect 8040 15290 8044 15346
rect 8044 15290 8100 15346
rect 8100 15290 8104 15346
rect 8040 15286 8104 15290
rect 8120 15346 8184 15350
rect 8120 15290 8124 15346
rect 8124 15290 8180 15346
rect 8180 15290 8184 15346
rect 8120 15286 8184 15290
rect 8200 15346 8264 15350
rect 8200 15290 8204 15346
rect 8204 15290 8260 15346
rect 8260 15290 8264 15346
rect 8200 15286 8264 15290
rect 8280 15346 8344 15350
rect 8280 15290 8284 15346
rect 8284 15290 8340 15346
rect 8340 15290 8344 15346
rect 8280 15286 8344 15290
rect 4960 14680 5024 14684
rect 4960 14624 4964 14680
rect 4964 14624 5020 14680
rect 5020 14624 5024 14680
rect 4960 14620 5024 14624
rect 5040 14680 5104 14684
rect 5040 14624 5044 14680
rect 5044 14624 5100 14680
rect 5100 14624 5104 14680
rect 5040 14620 5104 14624
rect 5120 14680 5184 14684
rect 5120 14624 5124 14680
rect 5124 14624 5180 14680
rect 5180 14624 5184 14680
rect 5120 14620 5184 14624
rect 5200 14680 5264 14684
rect 5200 14624 5204 14680
rect 5204 14624 5260 14680
rect 5260 14624 5264 14680
rect 5200 14620 5264 14624
rect 5280 14680 5344 14684
rect 5280 14624 5284 14680
rect 5284 14624 5340 14680
rect 5340 14624 5344 14680
rect 5280 14620 5344 14624
rect 1960 14014 2024 14018
rect 1960 13958 1964 14014
rect 1964 13958 2020 14014
rect 2020 13958 2024 14014
rect 1960 13954 2024 13958
rect 2040 14014 2104 14018
rect 2040 13958 2044 14014
rect 2044 13958 2100 14014
rect 2100 13958 2104 14014
rect 2040 13954 2104 13958
rect 2120 14014 2184 14018
rect 2120 13958 2124 14014
rect 2124 13958 2180 14014
rect 2180 13958 2184 14014
rect 2120 13954 2184 13958
rect 2200 14014 2264 14018
rect 2200 13958 2204 14014
rect 2204 13958 2260 14014
rect 2260 13958 2264 14014
rect 2200 13954 2264 13958
rect 2280 14014 2344 14018
rect 2280 13958 2284 14014
rect 2284 13958 2340 14014
rect 2340 13958 2344 14014
rect 2280 13954 2344 13958
rect 7960 14014 8024 14018
rect 7960 13958 7964 14014
rect 7964 13958 8020 14014
rect 8020 13958 8024 14014
rect 7960 13954 8024 13958
rect 8040 14014 8104 14018
rect 8040 13958 8044 14014
rect 8044 13958 8100 14014
rect 8100 13958 8104 14014
rect 8040 13954 8104 13958
rect 8120 14014 8184 14018
rect 8120 13958 8124 14014
rect 8124 13958 8180 14014
rect 8180 13958 8184 14014
rect 8120 13954 8184 13958
rect 8200 14014 8264 14018
rect 8200 13958 8204 14014
rect 8204 13958 8260 14014
rect 8260 13958 8264 14014
rect 8200 13954 8264 13958
rect 8280 14014 8344 14018
rect 8280 13958 8284 14014
rect 8284 13958 8340 14014
rect 8340 13958 8344 14014
rect 8280 13954 8344 13958
rect 4960 13348 5024 13352
rect 4960 13292 4964 13348
rect 4964 13292 5020 13348
rect 5020 13292 5024 13348
rect 4960 13288 5024 13292
rect 5040 13348 5104 13352
rect 5040 13292 5044 13348
rect 5044 13292 5100 13348
rect 5100 13292 5104 13348
rect 5040 13288 5104 13292
rect 5120 13348 5184 13352
rect 5120 13292 5124 13348
rect 5124 13292 5180 13348
rect 5180 13292 5184 13348
rect 5120 13288 5184 13292
rect 5200 13348 5264 13352
rect 5200 13292 5204 13348
rect 5204 13292 5260 13348
rect 5260 13292 5264 13348
rect 5200 13288 5264 13292
rect 5280 13348 5344 13352
rect 5280 13292 5284 13348
rect 5284 13292 5340 13348
rect 5340 13292 5344 13348
rect 5280 13288 5344 13292
rect 1960 12682 2024 12686
rect 1960 12626 1964 12682
rect 1964 12626 2020 12682
rect 2020 12626 2024 12682
rect 1960 12622 2024 12626
rect 2040 12682 2104 12686
rect 2040 12626 2044 12682
rect 2044 12626 2100 12682
rect 2100 12626 2104 12682
rect 2040 12622 2104 12626
rect 2120 12682 2184 12686
rect 2120 12626 2124 12682
rect 2124 12626 2180 12682
rect 2180 12626 2184 12682
rect 2120 12622 2184 12626
rect 2200 12682 2264 12686
rect 2200 12626 2204 12682
rect 2204 12626 2260 12682
rect 2260 12626 2264 12682
rect 2200 12622 2264 12626
rect 2280 12682 2344 12686
rect 2280 12626 2284 12682
rect 2284 12626 2340 12682
rect 2340 12626 2344 12682
rect 2280 12622 2344 12626
rect 7960 12682 8024 12686
rect 7960 12626 7964 12682
rect 7964 12626 8020 12682
rect 8020 12626 8024 12682
rect 7960 12622 8024 12626
rect 8040 12682 8104 12686
rect 8040 12626 8044 12682
rect 8044 12626 8100 12682
rect 8100 12626 8104 12682
rect 8040 12622 8104 12626
rect 8120 12682 8184 12686
rect 8120 12626 8124 12682
rect 8124 12626 8180 12682
rect 8180 12626 8184 12682
rect 8120 12622 8184 12626
rect 8200 12682 8264 12686
rect 8200 12626 8204 12682
rect 8204 12626 8260 12682
rect 8260 12626 8264 12682
rect 8200 12622 8264 12626
rect 8280 12682 8344 12686
rect 8280 12626 8284 12682
rect 8284 12626 8340 12682
rect 8340 12626 8344 12682
rect 8280 12622 8344 12626
rect 4960 12016 5024 12020
rect 4960 11960 4964 12016
rect 4964 11960 5020 12016
rect 5020 11960 5024 12016
rect 4960 11956 5024 11960
rect 5040 12016 5104 12020
rect 5040 11960 5044 12016
rect 5044 11960 5100 12016
rect 5100 11960 5104 12016
rect 5040 11956 5104 11960
rect 5120 12016 5184 12020
rect 5120 11960 5124 12016
rect 5124 11960 5180 12016
rect 5180 11960 5184 12016
rect 5120 11956 5184 11960
rect 5200 12016 5264 12020
rect 5200 11960 5204 12016
rect 5204 11960 5260 12016
rect 5260 11960 5264 12016
rect 5200 11956 5264 11960
rect 5280 12016 5344 12020
rect 5280 11960 5284 12016
rect 5284 11960 5340 12016
rect 5340 11960 5344 12016
rect 5280 11956 5344 11960
rect 1960 11350 2024 11354
rect 1960 11294 1964 11350
rect 1964 11294 2020 11350
rect 2020 11294 2024 11350
rect 1960 11290 2024 11294
rect 2040 11350 2104 11354
rect 2040 11294 2044 11350
rect 2044 11294 2100 11350
rect 2100 11294 2104 11350
rect 2040 11290 2104 11294
rect 2120 11350 2184 11354
rect 2120 11294 2124 11350
rect 2124 11294 2180 11350
rect 2180 11294 2184 11350
rect 2120 11290 2184 11294
rect 2200 11350 2264 11354
rect 2200 11294 2204 11350
rect 2204 11294 2260 11350
rect 2260 11294 2264 11350
rect 2200 11290 2264 11294
rect 2280 11350 2344 11354
rect 2280 11294 2284 11350
rect 2284 11294 2340 11350
rect 2340 11294 2344 11350
rect 2280 11290 2344 11294
rect 7960 11350 8024 11354
rect 7960 11294 7964 11350
rect 7964 11294 8020 11350
rect 8020 11294 8024 11350
rect 7960 11290 8024 11294
rect 8040 11350 8104 11354
rect 8040 11294 8044 11350
rect 8044 11294 8100 11350
rect 8100 11294 8104 11350
rect 8040 11290 8104 11294
rect 8120 11350 8184 11354
rect 8120 11294 8124 11350
rect 8124 11294 8180 11350
rect 8180 11294 8184 11350
rect 8120 11290 8184 11294
rect 8200 11350 8264 11354
rect 8200 11294 8204 11350
rect 8204 11294 8260 11350
rect 8260 11294 8264 11350
rect 8200 11290 8264 11294
rect 8280 11350 8344 11354
rect 8280 11294 8284 11350
rect 8284 11294 8340 11350
rect 8340 11294 8344 11350
rect 8280 11290 8344 11294
rect 4960 10684 5024 10688
rect 4960 10628 4964 10684
rect 4964 10628 5020 10684
rect 5020 10628 5024 10684
rect 4960 10624 5024 10628
rect 5040 10684 5104 10688
rect 5040 10628 5044 10684
rect 5044 10628 5100 10684
rect 5100 10628 5104 10684
rect 5040 10624 5104 10628
rect 5120 10684 5184 10688
rect 5120 10628 5124 10684
rect 5124 10628 5180 10684
rect 5180 10628 5184 10684
rect 5120 10624 5184 10628
rect 5200 10684 5264 10688
rect 5200 10628 5204 10684
rect 5204 10628 5260 10684
rect 5260 10628 5264 10684
rect 5200 10624 5264 10628
rect 5280 10684 5344 10688
rect 5280 10628 5284 10684
rect 5284 10628 5340 10684
rect 5340 10628 5344 10684
rect 5280 10624 5344 10628
rect 1960 10018 2024 10022
rect 1960 9962 1964 10018
rect 1964 9962 2020 10018
rect 2020 9962 2024 10018
rect 1960 9958 2024 9962
rect 2040 10018 2104 10022
rect 2040 9962 2044 10018
rect 2044 9962 2100 10018
rect 2100 9962 2104 10018
rect 2040 9958 2104 9962
rect 2120 10018 2184 10022
rect 2120 9962 2124 10018
rect 2124 9962 2180 10018
rect 2180 9962 2184 10018
rect 2120 9958 2184 9962
rect 2200 10018 2264 10022
rect 2200 9962 2204 10018
rect 2204 9962 2260 10018
rect 2260 9962 2264 10018
rect 2200 9958 2264 9962
rect 2280 10018 2344 10022
rect 2280 9962 2284 10018
rect 2284 9962 2340 10018
rect 2340 9962 2344 10018
rect 2280 9958 2344 9962
rect 7960 10018 8024 10022
rect 7960 9962 7964 10018
rect 7964 9962 8020 10018
rect 8020 9962 8024 10018
rect 7960 9958 8024 9962
rect 8040 10018 8104 10022
rect 8040 9962 8044 10018
rect 8044 9962 8100 10018
rect 8100 9962 8104 10018
rect 8040 9958 8104 9962
rect 8120 10018 8184 10022
rect 8120 9962 8124 10018
rect 8124 9962 8180 10018
rect 8180 9962 8184 10018
rect 8120 9958 8184 9962
rect 8200 10018 8264 10022
rect 8200 9962 8204 10018
rect 8204 9962 8260 10018
rect 8260 9962 8264 10018
rect 8200 9958 8264 9962
rect 8280 10018 8344 10022
rect 8280 9962 8284 10018
rect 8284 9962 8340 10018
rect 8340 9962 8344 10018
rect 8280 9958 8344 9962
rect 4960 9352 5024 9356
rect 4960 9296 4964 9352
rect 4964 9296 5020 9352
rect 5020 9296 5024 9352
rect 4960 9292 5024 9296
rect 5040 9352 5104 9356
rect 5040 9296 5044 9352
rect 5044 9296 5100 9352
rect 5100 9296 5104 9352
rect 5040 9292 5104 9296
rect 5120 9352 5184 9356
rect 5120 9296 5124 9352
rect 5124 9296 5180 9352
rect 5180 9296 5184 9352
rect 5120 9292 5184 9296
rect 5200 9352 5264 9356
rect 5200 9296 5204 9352
rect 5204 9296 5260 9352
rect 5260 9296 5264 9352
rect 5200 9292 5264 9296
rect 5280 9352 5344 9356
rect 5280 9296 5284 9352
rect 5284 9296 5340 9352
rect 5340 9296 5344 9352
rect 5280 9292 5344 9296
rect 1960 8686 2024 8690
rect 1960 8630 1964 8686
rect 1964 8630 2020 8686
rect 2020 8630 2024 8686
rect 1960 8626 2024 8630
rect 2040 8686 2104 8690
rect 2040 8630 2044 8686
rect 2044 8630 2100 8686
rect 2100 8630 2104 8686
rect 2040 8626 2104 8630
rect 2120 8686 2184 8690
rect 2120 8630 2124 8686
rect 2124 8630 2180 8686
rect 2180 8630 2184 8686
rect 2120 8626 2184 8630
rect 2200 8686 2264 8690
rect 2200 8630 2204 8686
rect 2204 8630 2260 8686
rect 2260 8630 2264 8686
rect 2200 8626 2264 8630
rect 2280 8686 2344 8690
rect 2280 8630 2284 8686
rect 2284 8630 2340 8686
rect 2340 8630 2344 8686
rect 2280 8626 2344 8630
rect 7960 8686 8024 8690
rect 7960 8630 7964 8686
rect 7964 8630 8020 8686
rect 8020 8630 8024 8686
rect 7960 8626 8024 8630
rect 8040 8686 8104 8690
rect 8040 8630 8044 8686
rect 8044 8630 8100 8686
rect 8100 8630 8104 8686
rect 8040 8626 8104 8630
rect 8120 8686 8184 8690
rect 8120 8630 8124 8686
rect 8124 8630 8180 8686
rect 8180 8630 8184 8686
rect 8120 8626 8184 8630
rect 8200 8686 8264 8690
rect 8200 8630 8204 8686
rect 8204 8630 8260 8686
rect 8260 8630 8264 8686
rect 8200 8626 8264 8630
rect 8280 8686 8344 8690
rect 8280 8630 8284 8686
rect 8284 8630 8340 8686
rect 8340 8630 8344 8686
rect 8280 8626 8344 8630
rect 4960 8020 5024 8024
rect 4960 7964 4964 8020
rect 4964 7964 5020 8020
rect 5020 7964 5024 8020
rect 4960 7960 5024 7964
rect 5040 8020 5104 8024
rect 5040 7964 5044 8020
rect 5044 7964 5100 8020
rect 5100 7964 5104 8020
rect 5040 7960 5104 7964
rect 5120 8020 5184 8024
rect 5120 7964 5124 8020
rect 5124 7964 5180 8020
rect 5180 7964 5184 8020
rect 5120 7960 5184 7964
rect 5200 8020 5264 8024
rect 5200 7964 5204 8020
rect 5204 7964 5260 8020
rect 5260 7964 5264 8020
rect 5200 7960 5264 7964
rect 5280 8020 5344 8024
rect 5280 7964 5284 8020
rect 5284 7964 5340 8020
rect 5340 7964 5344 8020
rect 5280 7960 5344 7964
rect 1960 7354 2024 7358
rect 1960 7298 1964 7354
rect 1964 7298 2020 7354
rect 2020 7298 2024 7354
rect 1960 7294 2024 7298
rect 2040 7354 2104 7358
rect 2040 7298 2044 7354
rect 2044 7298 2100 7354
rect 2100 7298 2104 7354
rect 2040 7294 2104 7298
rect 2120 7354 2184 7358
rect 2120 7298 2124 7354
rect 2124 7298 2180 7354
rect 2180 7298 2184 7354
rect 2120 7294 2184 7298
rect 2200 7354 2264 7358
rect 2200 7298 2204 7354
rect 2204 7298 2260 7354
rect 2260 7298 2264 7354
rect 2200 7294 2264 7298
rect 2280 7354 2344 7358
rect 2280 7298 2284 7354
rect 2284 7298 2340 7354
rect 2340 7298 2344 7354
rect 2280 7294 2344 7298
rect 7960 7354 8024 7358
rect 7960 7298 7964 7354
rect 7964 7298 8020 7354
rect 8020 7298 8024 7354
rect 7960 7294 8024 7298
rect 8040 7354 8104 7358
rect 8040 7298 8044 7354
rect 8044 7298 8100 7354
rect 8100 7298 8104 7354
rect 8040 7294 8104 7298
rect 8120 7354 8184 7358
rect 8120 7298 8124 7354
rect 8124 7298 8180 7354
rect 8180 7298 8184 7354
rect 8120 7294 8184 7298
rect 8200 7354 8264 7358
rect 8200 7298 8204 7354
rect 8204 7298 8260 7354
rect 8260 7298 8264 7354
rect 8200 7294 8264 7298
rect 8280 7354 8344 7358
rect 8280 7298 8284 7354
rect 8284 7298 8340 7354
rect 8340 7298 8344 7354
rect 8280 7294 8344 7298
rect 4960 6688 5024 6692
rect 4960 6632 4964 6688
rect 4964 6632 5020 6688
rect 5020 6632 5024 6688
rect 4960 6628 5024 6632
rect 5040 6688 5104 6692
rect 5040 6632 5044 6688
rect 5044 6632 5100 6688
rect 5100 6632 5104 6688
rect 5040 6628 5104 6632
rect 5120 6688 5184 6692
rect 5120 6632 5124 6688
rect 5124 6632 5180 6688
rect 5180 6632 5184 6688
rect 5120 6628 5184 6632
rect 5200 6688 5264 6692
rect 5200 6632 5204 6688
rect 5204 6632 5260 6688
rect 5260 6632 5264 6688
rect 5200 6628 5264 6632
rect 5280 6688 5344 6692
rect 5280 6632 5284 6688
rect 5284 6632 5340 6688
rect 5340 6632 5344 6688
rect 5280 6628 5344 6632
rect 1960 6022 2024 6026
rect 1960 5966 1964 6022
rect 1964 5966 2020 6022
rect 2020 5966 2024 6022
rect 1960 5962 2024 5966
rect 2040 6022 2104 6026
rect 2040 5966 2044 6022
rect 2044 5966 2100 6022
rect 2100 5966 2104 6022
rect 2040 5962 2104 5966
rect 2120 6022 2184 6026
rect 2120 5966 2124 6022
rect 2124 5966 2180 6022
rect 2180 5966 2184 6022
rect 2120 5962 2184 5966
rect 2200 6022 2264 6026
rect 2200 5966 2204 6022
rect 2204 5966 2260 6022
rect 2260 5966 2264 6022
rect 2200 5962 2264 5966
rect 2280 6022 2344 6026
rect 2280 5966 2284 6022
rect 2284 5966 2340 6022
rect 2340 5966 2344 6022
rect 2280 5962 2344 5966
rect 7960 6022 8024 6026
rect 7960 5966 7964 6022
rect 7964 5966 8020 6022
rect 8020 5966 8024 6022
rect 7960 5962 8024 5966
rect 8040 6022 8104 6026
rect 8040 5966 8044 6022
rect 8044 5966 8100 6022
rect 8100 5966 8104 6022
rect 8040 5962 8104 5966
rect 8120 6022 8184 6026
rect 8120 5966 8124 6022
rect 8124 5966 8180 6022
rect 8180 5966 8184 6022
rect 8120 5962 8184 5966
rect 8200 6022 8264 6026
rect 8200 5966 8204 6022
rect 8204 5966 8260 6022
rect 8260 5966 8264 6022
rect 8200 5962 8264 5966
rect 8280 6022 8344 6026
rect 8280 5966 8284 6022
rect 8284 5966 8340 6022
rect 8340 5966 8344 6022
rect 8280 5962 8344 5966
rect 4960 5356 5024 5360
rect 4960 5300 4964 5356
rect 4964 5300 5020 5356
rect 5020 5300 5024 5356
rect 4960 5296 5024 5300
rect 5040 5356 5104 5360
rect 5040 5300 5044 5356
rect 5044 5300 5100 5356
rect 5100 5300 5104 5356
rect 5040 5296 5104 5300
rect 5120 5356 5184 5360
rect 5120 5300 5124 5356
rect 5124 5300 5180 5356
rect 5180 5300 5184 5356
rect 5120 5296 5184 5300
rect 5200 5356 5264 5360
rect 5200 5300 5204 5356
rect 5204 5300 5260 5356
rect 5260 5300 5264 5356
rect 5200 5296 5264 5300
rect 5280 5356 5344 5360
rect 5280 5300 5284 5356
rect 5284 5300 5340 5356
rect 5340 5300 5344 5356
rect 5280 5296 5344 5300
rect 1960 4690 2024 4694
rect 1960 4634 1964 4690
rect 1964 4634 2020 4690
rect 2020 4634 2024 4690
rect 1960 4630 2024 4634
rect 2040 4690 2104 4694
rect 2040 4634 2044 4690
rect 2044 4634 2100 4690
rect 2100 4634 2104 4690
rect 2040 4630 2104 4634
rect 2120 4690 2184 4694
rect 2120 4634 2124 4690
rect 2124 4634 2180 4690
rect 2180 4634 2184 4690
rect 2120 4630 2184 4634
rect 2200 4690 2264 4694
rect 2200 4634 2204 4690
rect 2204 4634 2260 4690
rect 2260 4634 2264 4690
rect 2200 4630 2264 4634
rect 2280 4690 2344 4694
rect 2280 4634 2284 4690
rect 2284 4634 2340 4690
rect 2340 4634 2344 4690
rect 2280 4630 2344 4634
rect 7960 4690 8024 4694
rect 7960 4634 7964 4690
rect 7964 4634 8020 4690
rect 8020 4634 8024 4690
rect 7960 4630 8024 4634
rect 8040 4690 8104 4694
rect 8040 4634 8044 4690
rect 8044 4634 8100 4690
rect 8100 4634 8104 4690
rect 8040 4630 8104 4634
rect 8120 4690 8184 4694
rect 8120 4634 8124 4690
rect 8124 4634 8180 4690
rect 8180 4634 8184 4690
rect 8120 4630 8184 4634
rect 8200 4690 8264 4694
rect 8200 4634 8204 4690
rect 8204 4634 8260 4690
rect 8260 4634 8264 4690
rect 8200 4630 8264 4634
rect 8280 4690 8344 4694
rect 8280 4634 8284 4690
rect 8284 4634 8340 4690
rect 8340 4634 8344 4690
rect 8280 4630 8344 4634
rect 4960 4024 5024 4028
rect 4960 3968 4964 4024
rect 4964 3968 5020 4024
rect 5020 3968 5024 4024
rect 4960 3964 5024 3968
rect 5040 4024 5104 4028
rect 5040 3968 5044 4024
rect 5044 3968 5100 4024
rect 5100 3968 5104 4024
rect 5040 3964 5104 3968
rect 5120 4024 5184 4028
rect 5120 3968 5124 4024
rect 5124 3968 5180 4024
rect 5180 3968 5184 4024
rect 5120 3964 5184 3968
rect 5200 4024 5264 4028
rect 5200 3968 5204 4024
rect 5204 3968 5260 4024
rect 5260 3968 5264 4024
rect 5200 3964 5264 3968
rect 5280 4024 5344 4028
rect 5280 3968 5284 4024
rect 5284 3968 5340 4024
rect 5340 3968 5344 4024
rect 5280 3964 5344 3968
rect 1960 3358 2024 3362
rect 1960 3302 1964 3358
rect 1964 3302 2020 3358
rect 2020 3302 2024 3358
rect 1960 3298 2024 3302
rect 2040 3358 2104 3362
rect 2040 3302 2044 3358
rect 2044 3302 2100 3358
rect 2100 3302 2104 3358
rect 2040 3298 2104 3302
rect 2120 3358 2184 3362
rect 2120 3302 2124 3358
rect 2124 3302 2180 3358
rect 2180 3302 2184 3358
rect 2120 3298 2184 3302
rect 2200 3358 2264 3362
rect 2200 3302 2204 3358
rect 2204 3302 2260 3358
rect 2260 3302 2264 3358
rect 2200 3298 2264 3302
rect 2280 3358 2344 3362
rect 2280 3302 2284 3358
rect 2284 3302 2340 3358
rect 2340 3302 2344 3358
rect 2280 3298 2344 3302
rect 7960 3358 8024 3362
rect 7960 3302 7964 3358
rect 7964 3302 8020 3358
rect 8020 3302 8024 3358
rect 7960 3298 8024 3302
rect 8040 3358 8104 3362
rect 8040 3302 8044 3358
rect 8044 3302 8100 3358
rect 8100 3302 8104 3358
rect 8040 3298 8104 3302
rect 8120 3358 8184 3362
rect 8120 3302 8124 3358
rect 8124 3302 8180 3358
rect 8180 3302 8184 3358
rect 8120 3298 8184 3302
rect 8200 3358 8264 3362
rect 8200 3302 8204 3358
rect 8204 3302 8260 3358
rect 8260 3302 8264 3358
rect 8200 3298 8264 3302
rect 8280 3358 8344 3362
rect 8280 3302 8284 3358
rect 8284 3302 8340 3358
rect 8340 3302 8344 3358
rect 8280 3298 8344 3302
rect 4960 2692 5024 2696
rect 4960 2636 4964 2692
rect 4964 2636 5020 2692
rect 5020 2636 5024 2692
rect 4960 2632 5024 2636
rect 5040 2692 5104 2696
rect 5040 2636 5044 2692
rect 5044 2636 5100 2692
rect 5100 2636 5104 2692
rect 5040 2632 5104 2636
rect 5120 2692 5184 2696
rect 5120 2636 5124 2692
rect 5124 2636 5180 2692
rect 5180 2636 5184 2692
rect 5120 2632 5184 2636
rect 5200 2692 5264 2696
rect 5200 2636 5204 2692
rect 5204 2636 5260 2692
rect 5260 2636 5264 2692
rect 5200 2632 5264 2636
rect 5280 2692 5344 2696
rect 5280 2636 5284 2692
rect 5284 2636 5340 2692
rect 5340 2636 5344 2692
rect 5280 2632 5344 2636
<< metal4 >>
rect 1952 26006 2352 26022
rect 1952 25942 1960 26006
rect 2024 25942 2040 26006
rect 2104 25942 2120 26006
rect 2184 25942 2200 26006
rect 2264 25942 2280 26006
rect 2344 25942 2352 26006
rect 1952 24674 2352 25942
rect 1952 24610 1960 24674
rect 2024 24610 2040 24674
rect 2104 24610 2120 24674
rect 2184 24610 2200 24674
rect 2264 24610 2280 24674
rect 2344 24610 2352 24674
rect 1952 23342 2352 24610
rect 1952 23278 1960 23342
rect 2024 23278 2040 23342
rect 2104 23278 2120 23342
rect 2184 23278 2200 23342
rect 2264 23278 2280 23342
rect 2344 23278 2352 23342
rect 1952 22010 2352 23278
rect 1952 21946 1960 22010
rect 2024 21946 2040 22010
rect 2104 21946 2120 22010
rect 2184 21946 2200 22010
rect 2264 21946 2280 22010
rect 2344 21946 2352 22010
rect 1952 20678 2352 21946
rect 1952 20614 1960 20678
rect 2024 20614 2040 20678
rect 2104 20614 2120 20678
rect 2184 20614 2200 20678
rect 2264 20614 2280 20678
rect 2344 20614 2352 20678
rect 1952 19346 2352 20614
rect 1952 19282 1960 19346
rect 2024 19282 2040 19346
rect 2104 19282 2120 19346
rect 2184 19282 2200 19346
rect 2264 19282 2280 19346
rect 2344 19282 2352 19346
rect 1952 18014 2352 19282
rect 1952 17950 1960 18014
rect 2024 17950 2040 18014
rect 2104 17950 2120 18014
rect 2184 17950 2200 18014
rect 2264 17950 2280 18014
rect 2344 17950 2352 18014
rect 1952 16682 2352 17950
rect 1952 16618 1960 16682
rect 2024 16618 2040 16682
rect 2104 16618 2120 16682
rect 2184 16618 2200 16682
rect 2264 16618 2280 16682
rect 2344 16618 2352 16682
rect 1952 15350 2352 16618
rect 1952 15286 1960 15350
rect 2024 15286 2040 15350
rect 2104 15286 2120 15350
rect 2184 15286 2200 15350
rect 2264 15286 2280 15350
rect 2344 15286 2352 15350
rect 1952 14018 2352 15286
rect 1952 13954 1960 14018
rect 2024 13954 2040 14018
rect 2104 13954 2120 14018
rect 2184 13954 2200 14018
rect 2264 13954 2280 14018
rect 2344 13954 2352 14018
rect 1952 12686 2352 13954
rect 1952 12622 1960 12686
rect 2024 12622 2040 12686
rect 2104 12622 2120 12686
rect 2184 12622 2200 12686
rect 2264 12622 2280 12686
rect 2344 12622 2352 12686
rect 1952 11354 2352 12622
rect 1952 11290 1960 11354
rect 2024 11290 2040 11354
rect 2104 11290 2120 11354
rect 2184 11290 2200 11354
rect 2264 11290 2280 11354
rect 2344 11290 2352 11354
rect 1952 10022 2352 11290
rect 1952 9958 1960 10022
rect 2024 9958 2040 10022
rect 2104 9958 2120 10022
rect 2184 9958 2200 10022
rect 2264 9958 2280 10022
rect 2344 9958 2352 10022
rect 1952 8690 2352 9958
rect 1952 8626 1960 8690
rect 2024 8626 2040 8690
rect 2104 8626 2120 8690
rect 2184 8626 2200 8690
rect 2264 8626 2280 8690
rect 2344 8626 2352 8690
rect 1952 7358 2352 8626
rect 1952 7294 1960 7358
rect 2024 7294 2040 7358
rect 2104 7294 2120 7358
rect 2184 7294 2200 7358
rect 2264 7294 2280 7358
rect 2344 7294 2352 7358
rect 1952 6026 2352 7294
rect 1952 5962 1960 6026
rect 2024 5962 2040 6026
rect 2104 5962 2120 6026
rect 2184 5962 2200 6026
rect 2264 5962 2280 6026
rect 2344 5962 2352 6026
rect 1952 4694 2352 5962
rect 1952 4630 1960 4694
rect 2024 4630 2040 4694
rect 2104 4630 2120 4694
rect 2184 4630 2200 4694
rect 2264 4630 2280 4694
rect 2344 4630 2352 4694
rect 1952 3362 2352 4630
rect 1952 3298 1960 3362
rect 2024 3298 2040 3362
rect 2104 3298 2120 3362
rect 2184 3298 2200 3362
rect 2264 3298 2280 3362
rect 2344 3298 2352 3362
rect 1952 2616 2352 3298
rect 4952 25340 5352 26022
rect 4952 25276 4960 25340
rect 5024 25276 5040 25340
rect 5104 25276 5120 25340
rect 5184 25276 5200 25340
rect 5264 25276 5280 25340
rect 5344 25276 5352 25340
rect 4952 24008 5352 25276
rect 4952 23944 4960 24008
rect 5024 23944 5040 24008
rect 5104 23944 5120 24008
rect 5184 23944 5200 24008
rect 5264 23944 5280 24008
rect 5344 23944 5352 24008
rect 4952 22676 5352 23944
rect 4952 22612 4960 22676
rect 5024 22612 5040 22676
rect 5104 22612 5120 22676
rect 5184 22612 5200 22676
rect 5264 22612 5280 22676
rect 5344 22612 5352 22676
rect 4952 21344 5352 22612
rect 4952 21280 4960 21344
rect 5024 21280 5040 21344
rect 5104 21280 5120 21344
rect 5184 21280 5200 21344
rect 5264 21280 5280 21344
rect 5344 21280 5352 21344
rect 4952 20012 5352 21280
rect 4952 19948 4960 20012
rect 5024 19948 5040 20012
rect 5104 19948 5120 20012
rect 5184 19948 5200 20012
rect 5264 19948 5280 20012
rect 5344 19948 5352 20012
rect 4952 18680 5352 19948
rect 4952 18616 4960 18680
rect 5024 18616 5040 18680
rect 5104 18616 5120 18680
rect 5184 18616 5200 18680
rect 5264 18616 5280 18680
rect 5344 18616 5352 18680
rect 4952 17348 5352 18616
rect 4952 17284 4960 17348
rect 5024 17284 5040 17348
rect 5104 17284 5120 17348
rect 5184 17284 5200 17348
rect 5264 17284 5280 17348
rect 5344 17284 5352 17348
rect 4952 16016 5352 17284
rect 4952 15952 4960 16016
rect 5024 15952 5040 16016
rect 5104 15952 5120 16016
rect 5184 15952 5200 16016
rect 5264 15952 5280 16016
rect 5344 15952 5352 16016
rect 4952 14684 5352 15952
rect 4952 14620 4960 14684
rect 5024 14620 5040 14684
rect 5104 14620 5120 14684
rect 5184 14620 5200 14684
rect 5264 14620 5280 14684
rect 5344 14620 5352 14684
rect 4952 13352 5352 14620
rect 4952 13288 4960 13352
rect 5024 13288 5040 13352
rect 5104 13288 5120 13352
rect 5184 13288 5200 13352
rect 5264 13288 5280 13352
rect 5344 13288 5352 13352
rect 4952 12020 5352 13288
rect 4952 11956 4960 12020
rect 5024 11956 5040 12020
rect 5104 11956 5120 12020
rect 5184 11956 5200 12020
rect 5264 11956 5280 12020
rect 5344 11956 5352 12020
rect 4952 10688 5352 11956
rect 4952 10624 4960 10688
rect 5024 10624 5040 10688
rect 5104 10624 5120 10688
rect 5184 10624 5200 10688
rect 5264 10624 5280 10688
rect 5344 10624 5352 10688
rect 4952 9356 5352 10624
rect 4952 9292 4960 9356
rect 5024 9292 5040 9356
rect 5104 9292 5120 9356
rect 5184 9292 5200 9356
rect 5264 9292 5280 9356
rect 5344 9292 5352 9356
rect 4952 8024 5352 9292
rect 4952 7960 4960 8024
rect 5024 7960 5040 8024
rect 5104 7960 5120 8024
rect 5184 7960 5200 8024
rect 5264 7960 5280 8024
rect 5344 7960 5352 8024
rect 4952 6692 5352 7960
rect 4952 6628 4960 6692
rect 5024 6628 5040 6692
rect 5104 6628 5120 6692
rect 5184 6628 5200 6692
rect 5264 6628 5280 6692
rect 5344 6628 5352 6692
rect 4952 5360 5352 6628
rect 4952 5296 4960 5360
rect 5024 5296 5040 5360
rect 5104 5296 5120 5360
rect 5184 5296 5200 5360
rect 5264 5296 5280 5360
rect 5344 5296 5352 5360
rect 4952 4028 5352 5296
rect 4952 3964 4960 4028
rect 5024 3964 5040 4028
rect 5104 3964 5120 4028
rect 5184 3964 5200 4028
rect 5264 3964 5280 4028
rect 5344 3964 5352 4028
rect 4952 2696 5352 3964
rect 4952 2632 4960 2696
rect 5024 2632 5040 2696
rect 5104 2632 5120 2696
rect 5184 2632 5200 2696
rect 5264 2632 5280 2696
rect 5344 2632 5352 2696
rect 4952 2616 5352 2632
rect 7952 26006 8352 26022
rect 7952 25942 7960 26006
rect 8024 25942 8040 26006
rect 8104 25942 8120 26006
rect 8184 25942 8200 26006
rect 8264 25942 8280 26006
rect 8344 25942 8352 26006
rect 7952 24674 8352 25942
rect 7952 24610 7960 24674
rect 8024 24610 8040 24674
rect 8104 24610 8120 24674
rect 8184 24610 8200 24674
rect 8264 24610 8280 24674
rect 8344 24610 8352 24674
rect 7952 23342 8352 24610
rect 7952 23278 7960 23342
rect 8024 23278 8040 23342
rect 8104 23278 8120 23342
rect 8184 23278 8200 23342
rect 8264 23278 8280 23342
rect 8344 23278 8352 23342
rect 7952 22010 8352 23278
rect 7952 21946 7960 22010
rect 8024 21946 8040 22010
rect 8104 21946 8120 22010
rect 8184 21946 8200 22010
rect 8264 21946 8280 22010
rect 8344 21946 8352 22010
rect 7952 20678 8352 21946
rect 7952 20614 7960 20678
rect 8024 20614 8040 20678
rect 8104 20614 8120 20678
rect 8184 20614 8200 20678
rect 8264 20614 8280 20678
rect 8344 20614 8352 20678
rect 7952 19346 8352 20614
rect 7952 19282 7960 19346
rect 8024 19282 8040 19346
rect 8104 19282 8120 19346
rect 8184 19282 8200 19346
rect 8264 19282 8280 19346
rect 8344 19282 8352 19346
rect 7952 18014 8352 19282
rect 7952 17950 7960 18014
rect 8024 17950 8040 18014
rect 8104 17950 8120 18014
rect 8184 17950 8200 18014
rect 8264 17950 8280 18014
rect 8344 17950 8352 18014
rect 7952 16682 8352 17950
rect 7952 16618 7960 16682
rect 8024 16618 8040 16682
rect 8104 16618 8120 16682
rect 8184 16618 8200 16682
rect 8264 16618 8280 16682
rect 8344 16618 8352 16682
rect 7952 15350 8352 16618
rect 7952 15286 7960 15350
rect 8024 15286 8040 15350
rect 8104 15286 8120 15350
rect 8184 15286 8200 15350
rect 8264 15286 8280 15350
rect 8344 15286 8352 15350
rect 7952 14018 8352 15286
rect 7952 13954 7960 14018
rect 8024 13954 8040 14018
rect 8104 13954 8120 14018
rect 8184 13954 8200 14018
rect 8264 13954 8280 14018
rect 8344 13954 8352 14018
rect 7952 12686 8352 13954
rect 7952 12622 7960 12686
rect 8024 12622 8040 12686
rect 8104 12622 8120 12686
rect 8184 12622 8200 12686
rect 8264 12622 8280 12686
rect 8344 12622 8352 12686
rect 7952 11354 8352 12622
rect 7952 11290 7960 11354
rect 8024 11290 8040 11354
rect 8104 11290 8120 11354
rect 8184 11290 8200 11354
rect 8264 11290 8280 11354
rect 8344 11290 8352 11354
rect 7952 10022 8352 11290
rect 7952 9958 7960 10022
rect 8024 9958 8040 10022
rect 8104 9958 8120 10022
rect 8184 9958 8200 10022
rect 8264 9958 8280 10022
rect 8344 9958 8352 10022
rect 7952 8690 8352 9958
rect 7952 8626 7960 8690
rect 8024 8626 8040 8690
rect 8104 8626 8120 8690
rect 8184 8626 8200 8690
rect 8264 8626 8280 8690
rect 8344 8626 8352 8690
rect 7952 7358 8352 8626
rect 7952 7294 7960 7358
rect 8024 7294 8040 7358
rect 8104 7294 8120 7358
rect 8184 7294 8200 7358
rect 8264 7294 8280 7358
rect 8344 7294 8352 7358
rect 7952 6026 8352 7294
rect 7952 5962 7960 6026
rect 8024 5962 8040 6026
rect 8104 5962 8120 6026
rect 8184 5962 8200 6026
rect 8264 5962 8280 6026
rect 8344 5962 8352 6026
rect 7952 4694 8352 5962
rect 7952 4630 7960 4694
rect 8024 4630 8040 4694
rect 8104 4630 8120 4694
rect 8184 4630 8200 4694
rect 8264 4630 8280 4694
rect 8344 4630 8352 4694
rect 7952 3362 8352 4630
rect 7952 3298 7960 3362
rect 8024 3298 8040 3362
rect 8104 3298 8120 3362
rect 8184 3298 8200 3362
rect 8264 3298 8280 3362
rect 8344 3298 8352 3362
rect 7952 2616 8352 3298
use sky130_fd_sc_hs__and2_1  _18_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749223325
transform 1 0 7872 0 1 22644
box -38 -49 518 715
use sky130_fd_sc_hs__clkbuf_1  _19_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 8736 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__or4bb_1  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 9120 0 -1 6660
box -38 -49 998 715
use sky130_fd_sc_hs__nand2_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749010377
transform -1 0 5088 0 1 5328
box -38 -49 326 715
use sky130_fd_sc_hs__or3b_1  _22_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 5088 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__o21a_1  _23_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 6240 0 1 3996
box -38 -49 614 715
use sky130_fd_sc_hs__and2_1  _24_
timestamp 1749223325
transform -1 0 6336 0 -1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__a21bo_1  _25_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 6336 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__clkbuf_1  _26_
timestamp 1704896540
transform 1 0 5184 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__nor2_1  _27_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 6528 0 1 3996
box -38 -49 326 715
use sky130_fd_sc_hs__xor2_1  _28_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 9120 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__and2_1  _29_
timestamp 1749223325
transform 1 0 8256 0 1 3996
box -38 -49 518 715
use sky130_fd_sc_hs__clkbuf_1  _30_
timestamp 1704896540
transform -1 0 9504 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__and3_1  _31_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 9024 0 1 5328
box -38 -49 614 715
use sky130_fd_sc_hs__a21oi_1  _32_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 9120 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__nor3_1  _33_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 9984 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__xor2_1  _34_
timestamp 1704896540
transform -1 0 8928 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__and2_1  _35_
timestamp 1749223325
transform -1 0 8352 0 -1 7992
box -38 -49 518 715
use sky130_fd_sc_hs__clkbuf_1  _36_
timestamp 1704896540
transform -1 0 7200 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__dfxtp_1  _37_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 6240 0 -1 5328
box -38 -49 1670 715
use sky130_fd_sc_hs__dfxtp_4  _38_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 6432 0 -1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__dfrtp_1  _39_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 3744 0 1 6660
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _40_
timestamp 1704896540
transform 1 0 1632 0 -1 7992
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _41_
timestamp 1704896540
transform -1 0 3840 0 -1 6660
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _42_
timestamp 1704896540
transform 1 0 1536 0 1 11988
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _43_
timestamp 1704896540
transform -1 0 3744 0 1 14652
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _44_
timestamp 1704896540
transform -1 0 3744 0 1 15984
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _45_
timestamp 1704896540
transform -1 0 3744 0 1 17316
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _46_
timestamp 1704896540
transform -1 0 3744 0 1 18648
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _47_
timestamp 1704896540
transform -1 0 3744 0 1 19980
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _48_
timestamp 1704896540
transform 1 0 1536 0 1 21312
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_2  _49_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 3840 0 1 21312
box -38 -49 2342 715
use sky130_fd_sc_hs__dfxtp_1  _50_
timestamp 1704896540
transform 1 0 6528 0 -1 3996
box -38 -49 1670 715
use sky130_fd_sc_hs__dfxtp_1  _51_
timestamp 1704896540
transform 1 0 6624 0 1 3996
box -38 -49 1670 715
use sky130_fd_sc_hs__dfxtp_1  _52_
timestamp 1704896540
transform 1 0 6528 0 -1 6660
box -38 -49 1670 715
use sky130_fd_sc_hs__dfxtp_1  _53_
timestamp 1704896540
transform 1 0 6240 0 1 6660
box -38 -49 1670 715
use sky130_fd_sc_hs__dfrtp_1  _54_
timestamp 1704896540
transform 1 0 6432 0 -1 23976
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _55_
timestamp 1704896540
transform 1 0 5568 0 1 22644
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _56_
timestamp 1704896540
transform 1 0 5376 0 1 19980
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _57_
timestamp 1704896540
transform 1 0 4992 0 1 18648
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _58_
timestamp 1704896540
transform 1 0 4416 0 1 17316
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _59_
timestamp 1704896540
transform 1 0 3552 0 -1 17316
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _60_
timestamp 1704896540
transform 1 0 2880 0 -1 15984
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _61_
timestamp 1704896540
transform 1 0 2400 0 -1 11988
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _62_
timestamp 1704896540
transform 1 0 2304 0 -1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _63_
timestamp 1704896540
transform 1 0 1536 0 1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _64_
timestamp 1704896540
transform 1 0 6240 0 1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _65_
timestamp 1704896540
transform 1 0 6144 0 1 11988
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _66_
timestamp 1704896540
transform 1 0 6432 0 -1 11988
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _67_
timestamp 1704896540
transform 1 0 5088 0 1 13320
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _68_
timestamp 1704896540
transform 1 0 4128 0 -1 14652
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _69_
timestamp 1704896540
transform 1 0 2976 0 -1 13320
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _70_
timestamp 1704896540
transform 1 0 3840 0 1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _71_
timestamp 1704896540
transform 1 0 1632 0 -1 5328
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _72_
timestamp 1704896540
transform -1 0 3744 0 1 3996
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _73_
timestamp 1704896540
transform 1 0 1536 0 1 5328
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _74_
timestamp 1704896540
transform 1 0 7776 0 -1 22644
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _75_
timestamp 1704896540
transform 1 0 7776 0 -1 21312
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _76_
timestamp 1704896540
transform 1 0 7776 0 -1 19980
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _77_
timestamp 1704896540
transform 1 0 7776 0 -1 17316
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _78_
timestamp 1704896540
transform 1 0 7776 0 -1 18648
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _79_
timestamp 1704896540
transform 1 0 7488 0 -1 15984
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _80_
timestamp 1704896540
transform 1 0 7488 0 -1 14652
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _81_
timestamp 1704896540
transform 1 0 7680 0 -1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _82_
timestamp 1704896540
transform 1 0 7776 0 -1 13320
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _83_
timestamp 1704896540
transform 1 0 7776 0 -1 9324
box -38 -49 2246 715
use sky130_fd_sc_hs__clkbuf_16  clkbuf_0_CLK $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 6336 0 1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__clkbuf_16  clkbuf_1_0__f_CLK
timestamp 1704896540
transform 1 0 6912 0 1 2664
box -38 -49 1958 715
use sky130_fd_sc_hs__clkbuf_16  clkbuf_1_1__f_CLK
timestamp 1704896540
transform -1 0 8064 0 1 7992
box -38 -49 1958 715
use sky130_fd_sc_hs__fill_2  FILLER_0_0_4 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 1536 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 1728 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_0_23 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 3360 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_0_28
timestamp 1704896540
transform 1 0 3840 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_0_30
timestamp 1704896540
transform 1 0 4032 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_0_35 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 4512 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_0_47
timestamp 1704896540
transform 1 0 5664 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_0_51
timestamp 1704896540
transform 1 0 6048 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_0_53
timestamp 1704896540
transform 1 0 6240 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_0_59
timestamp 1704896540
transform 1 0 6816 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_0_80
timestamp 1704896540
transform 1 0 8832 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_1_16
timestamp 1704896540
transform 1 0 2688 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_1_24
timestamp 1704896540
transform 1 0 3456 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_1_32
timestamp 1704896540
transform 1 0 4224 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_1_40
timestamp 1704896540
transform 1 0 4992 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_1_48
timestamp 1704896540
transform 1 0 5760 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 6432 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_1_77
timestamp 1704896540
transform 1 0 8544 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_1_85
timestamp 1704896540
transform 1 0 9312 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_2_28
timestamp 1704896540
transform 1 0 3840 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_2_36
timestamp 1704896540
transform 1 0 4608 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_2_44
timestamp 1704896540
transform 1 0 5376 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_2_46
timestamp 1704896540
transform 1 0 5568 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_2_56
timestamp 1704896540
transform 1 0 6528 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_2_79
timestamp 1704896540
transform 1 0 8736 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_2_82
timestamp 1704896540
transform 1 0 9024 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_2_90
timestamp 1704896540
transform 1 0 9792 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_3_4
timestamp 1704896540
transform 1 0 1536 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_3_28
timestamp 1704896540
transform 1 0 3840 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_3_53
timestamp 1704896540
transform 1 0 6240 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_3_87
timestamp 1704896540
transform 1 0 9504 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_3_91
timestamp 1704896540
transform 1 0 9888 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_3_93
timestamp 1704896540
transform 1 0 10080 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_4_28
timestamp 1704896540
transform 1 0 3840 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_4_36
timestamp 1704896540
transform 1 0 4608 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_4_49
timestamp 1704896540
transform 1 0 5856 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_4_53
timestamp 1704896540
transform 1 0 6240 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_4_74
timestamp 1704896540
transform 1 0 8256 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_4_78
timestamp 1704896540
transform 1 0 8640 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_4_80
timestamp 1704896540
transform 1 0 8832 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_4_92
timestamp 1704896540
transform 1 0 9984 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_5_4
timestamp 1704896540
transform 1 0 1536 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_5_28
timestamp 1704896540
transform 1 0 3840 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_5_36
timestamp 1704896540
transform 1 0 4608 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_5_40
timestamp 1704896540
transform 1 0 4992 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 6432 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_5_87
timestamp 1704896540
transform 1 0 9504 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_5_89
timestamp 1704896540
transform 1 0 9696 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_6_28
timestamp 1704896540
transform 1 0 3840 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_6_36
timestamp 1704896540
transform 1 0 4608 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_6_44
timestamp 1704896540
transform 1 0 5376 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_6_52
timestamp 1704896540
transform 1 0 6144 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_6_70
timestamp 1704896540
transform 1 0 7872 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_6_72
timestamp 1704896540
transform 1 0 8064 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_6_82
timestamp 1704896540
transform 1 0 9024 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_6_90
timestamp 1704896540
transform 1 0 9792 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_7_4
timestamp 1704896540
transform 1 0 1536 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_7_28
timestamp 1704896540
transform 1 0 3840 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_7_36
timestamp 1704896540
transform 1 0 4608 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_7_44
timestamp 1704896540
transform 1 0 5376 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_7_52
timestamp 1704896540
transform 1 0 6144 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6432 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  FILLER_0_7_63
timestamp 1704896540
transform 1 0 7200 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_7_67
timestamp 1704896540
transform 1 0 7584 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_7_69
timestamp 1704896540
transform 1 0 7776 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_7_75
timestamp 1704896540
transform 1 0 8352 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_7_83
timestamp 1704896540
transform 1 0 9120 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_7_91
timestamp 1704896540
transform 1 0 9888 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_7_93
timestamp 1704896540
transform 1 0 10080 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_8_10
timestamp 1704896540
transform 1 0 2112 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_8_18
timestamp 1704896540
transform 1 0 2880 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_8_26
timestamp 1704896540
transform 1 0 3648 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_8_28
timestamp 1704896540
transform 1 0 3840 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_8_36
timestamp 1704896540
transform 1 0 4608 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_8_44
timestamp 1704896540
transform 1 0 5376 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_8_72
timestamp 1704896540
transform 1 0 8064 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_8_80
timestamp 1704896540
transform 1 0 8832 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_8_82
timestamp 1704896540
transform 1 0 9024 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_9_8
timestamp 1704896540
transform 1 0 1920 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_9_16
timestamp 1704896540
transform 1 0 2688 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_9_24
timestamp 1704896540
transform 1 0 3456 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_9_32
timestamp 1704896540
transform 1 0 4224 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_9_40
timestamp 1704896540
transform 1 0 4992 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_9_48
timestamp 1704896540
transform 1 0 5760 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_9_52
timestamp 1704896540
transform 1 0 6144 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_9_55
timestamp 1704896540
transform 1 0 6432 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_9_63
timestamp 1704896540
transform 1 0 7200 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_9_67
timestamp 1704896540
transform 1 0 7584 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_9_92
timestamp 1704896540
transform 1 0 9984 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_4
timestamp 1704896540
transform 1 0 1536 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_12
timestamp 1704896540
transform 1 0 2304 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_10_20
timestamp 1704896540
transform 1 0 3072 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_10_24
timestamp 1704896540
transform 1 0 3456 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_10_26
timestamp 1704896540
transform 1 0 3648 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_28
timestamp 1704896540
transform 1 0 3840 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_36
timestamp 1704896540
transform 1 0 4608 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_44
timestamp 1704896540
transform 1 0 5376 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_52
timestamp 1704896540
transform 1 0 6144 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_60
timestamp 1704896540
transform 1 0 6912 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_68
timestamp 1704896540
transform 1 0 7680 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_10_76
timestamp 1704896540
transform 1 0 8448 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_10_80
timestamp 1704896540
transform 1 0 8832 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_82
timestamp 1704896540
transform 1 0 9024 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_10_90
timestamp 1704896540
transform 1 0 9792 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  FILLER_0_11_8
timestamp 1704896540
transform 1 0 1920 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_11_35
timestamp 1704896540
transform 1 0 4512 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_11_43
timestamp 1704896540
transform 1 0 5280 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_11_51
timestamp 1704896540
transform 1 0 6048 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_11_53
timestamp 1704896540
transform 1 0 6240 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_11_55
timestamp 1704896540
transform 1 0 6432 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_11_63
timestamp 1704896540
transform 1 0 7200 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_11_67
timestamp 1704896540
transform 1 0 7584 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_11_91
timestamp 1704896540
transform 1 0 9888 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_11_93
timestamp 1704896540
transform 1 0 10080 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_12_51
timestamp 1704896540
transform 1 0 6048 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_12_76
timestamp 1704896540
transform 1 0 8448 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_12_80
timestamp 1704896540
transform 1 0 8832 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_12_82
timestamp 1704896540
transform 1 0 9024 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_13_8
timestamp 1704896540
transform 1 0 1920 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_13_12
timestamp 1704896540
transform 1 0 2304 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_36
timestamp 1704896540
transform 1 0 4608 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_44
timestamp 1704896540
transform 1 0 5376 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_13_52
timestamp 1704896540
transform 1 0 6144 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_78
timestamp 1704896540
transform 1 0 8640 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_86
timestamp 1704896540
transform 1 0 9408 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_14_28
timestamp 1704896540
transform 1 0 3840 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_14_36
timestamp 1704896540
transform 1 0 4608 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_14_44
timestamp 1704896540
transform 1 0 5376 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_14_75
timestamp 1704896540
transform 1 0 8352 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_14_79
timestamp 1704896540
transform 1 0 8736 0 1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_14_82
timestamp 1704896540
transform 1 0 9024 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_14_90
timestamp 1704896540
transform 1 0 9792 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_15_8
timestamp 1704896540
transform 1 0 1920 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_15_16
timestamp 1704896540
transform 1 0 2688 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_15_18
timestamp 1704896540
transform 1 0 2880 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_15_42
timestamp 1704896540
transform 1 0 5184 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_15_50
timestamp 1704896540
transform 1 0 5952 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_15_55
timestamp 1704896540
transform 1 0 6432 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_15_63
timestamp 1704896540
transform 1 0 7200 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_15_67
timestamp 1704896540
transform 1 0 7584 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_15_92
timestamp 1704896540
transform 1 0 9984 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_4
timestamp 1704896540
transform 1 0 1536 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_12
timestamp 1704896540
transform 1 0 2304 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_16_20
timestamp 1704896540
transform 1 0 3072 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_16_24
timestamp 1704896540
transform 1 0 3456 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_16_26
timestamp 1704896540
transform 1 0 3648 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_28
timestamp 1704896540
transform 1 0 3840 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_16_36
timestamp 1704896540
transform 1 0 4608 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_16_40
timestamp 1704896540
transform 1 0 4992 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_64
timestamp 1704896540
transform 1 0 7296 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_72
timestamp 1704896540
transform 1 0 8064 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_16_80
timestamp 1704896540
transform 1 0 8832 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_82
timestamp 1704896540
transform 1 0 9024 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_17_8
timestamp 1704896540
transform 1 0 1920 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_17_16
timestamp 1704896540
transform 1 0 2688 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_17_24
timestamp 1704896540
transform 1 0 3456 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_17_28
timestamp 1704896540
transform 1 0 3840 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_17_30
timestamp 1704896540
transform 1 0 4032 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_17_55
timestamp 1704896540
transform 1 0 6432 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_17_63
timestamp 1704896540
transform 1 0 7200 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_17_65
timestamp 1704896540
transform 1 0 7392 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_17_89
timestamp 1704896540
transform 1 0 9696 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_17_93
timestamp 1704896540
transform 1 0 10080 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_18_28
timestamp 1704896540
transform 1 0 3840 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_18_36
timestamp 1704896540
transform 1 0 4608 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_18_44
timestamp 1704896540
transform 1 0 5376 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_18_52
timestamp 1704896540
transform 1 0 6144 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_18_60
timestamp 1704896540
transform 1 0 6912 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_18_68
timestamp 1704896540
transform 1 0 7680 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_18_76
timestamp 1704896540
transform 1 0 8448 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_18_80
timestamp 1704896540
transform 1 0 8832 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_18_82
timestamp 1704896540
transform 1 0 9024 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_18_90
timestamp 1704896540
transform 1 0 9792 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_19_8
timestamp 1704896540
transform 1 0 1920 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_19_16
timestamp 1704896540
transform 1 0 2688 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_19_41
timestamp 1704896540
transform 1 0 5088 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_19_49
timestamp 1704896540
transform 1 0 5856 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_19_53
timestamp 1704896540
transform 1 0 6240 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_19_55
timestamp 1704896540
transform 1 0 6432 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_19_63
timestamp 1704896540
transform 1 0 7200 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_19_65
timestamp 1704896540
transform 1 0 7392 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_19_89
timestamp 1704896540
transform 1 0 9696 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_20_28
timestamp 1704896540
transform 1 0 3840 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_20_36
timestamp 1704896540
transform 1 0 4608 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_20_44
timestamp 1704896540
transform 1 0 5376 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_20_52
timestamp 1704896540
transform 1 0 6144 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_20_60
timestamp 1704896540
transform 1 0 6912 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_20_68
timestamp 1704896540
transform 1 0 7680 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_20_76
timestamp 1704896540
transform 1 0 8448 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_20_80
timestamp 1704896540
transform 1 0 8832 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_20_82
timestamp 1704896540
transform 1 0 9024 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_20_90
timestamp 1704896540
transform 1 0 9792 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_21_8
timestamp 1704896540
transform 1 0 1920 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_21_16
timestamp 1704896540
transform 1 0 2688 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_21_24
timestamp 1704896540
transform 1 0 3456 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_21_48
timestamp 1704896540
transform 1 0 5760 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_21_52
timestamp 1704896540
transform 1 0 6144 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_21_55
timestamp 1704896540
transform 1 0 6432 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_21_63
timestamp 1704896540
transform 1 0 7200 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_21_67
timestamp 1704896540
transform 1 0 7584 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_21_92
timestamp 1704896540
transform 1 0 9984 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_22_28
timestamp 1704896540
transform 1 0 3840 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_22_32
timestamp 1704896540
transform 1 0 4224 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_22_57
timestamp 1704896540
transform 1 0 6624 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_22_65
timestamp 1704896540
transform 1 0 7392 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_22_73
timestamp 1704896540
transform 1 0 8160 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_22_82
timestamp 1704896540
transform 1 0 9024 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_23_8
timestamp 1704896540
transform 1 0 1920 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_23_16
timestamp 1704896540
transform 1 0 2688 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_23_24
timestamp 1704896540
transform 1 0 3456 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_23_32
timestamp 1704896540
transform 1 0 4224 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_23_40
timestamp 1704896540
transform 1 0 4992 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_23_48
timestamp 1704896540
transform 1 0 5760 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_23_52
timestamp 1704896540
transform 1 0 6144 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_23_55
timestamp 1704896540
transform 1 0 6432 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_23_63
timestamp 1704896540
transform 1 0 7200 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_23_67
timestamp 1704896540
transform 1 0 7584 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_23_92
timestamp 1704896540
transform 1 0 9984 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_24_28
timestamp 1704896540
transform 1 0 3840 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_24_36
timestamp 1704896540
transform 1 0 4608 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_24_63
timestamp 1704896540
transform 1 0 7200 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_24_71
timestamp 1704896540
transform 1 0 7968 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_24_79
timestamp 1704896540
transform 1 0 8736 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_24_82
timestamp 1704896540
transform 1 0 9024 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_24_90
timestamp 1704896540
transform 1 0 9792 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_25_8
timestamp 1704896540
transform 1 0 1920 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_25_16
timestamp 1704896540
transform 1 0 2688 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_25_24
timestamp 1704896540
transform 1 0 3456 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_25_32
timestamp 1704896540
transform 1 0 4224 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_25_40
timestamp 1704896540
transform 1 0 4992 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_25_48
timestamp 1704896540
transform 1 0 5760 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_25_52
timestamp 1704896540
transform 1 0 6144 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_25_55
timestamp 1704896540
transform 1 0 6432 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_25_63
timestamp 1704896540
transform 1 0 7200 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_25_67
timestamp 1704896540
transform 1 0 7584 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_25_92
timestamp 1704896540
transform 1 0 9984 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_26_28
timestamp 1704896540
transform 1 0 3840 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_26_36
timestamp 1704896540
transform 1 0 4608 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_26_67
timestamp 1704896540
transform 1 0 7584 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_26_75
timestamp 1704896540
transform 1 0 8352 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_26_79
timestamp 1704896540
transform 1 0 8736 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_26_82
timestamp 1704896540
transform 1 0 9024 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_27_4
timestamp 1704896540
transform 1 0 1536 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_27_12
timestamp 1704896540
transform 1 0 2304 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_27_20
timestamp 1704896540
transform 1 0 3072 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_27_28
timestamp 1704896540
transform 1 0 3840 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_27_36
timestamp 1704896540
transform 1 0 4608 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_27_44
timestamp 1704896540
transform 1 0 5376 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_27_52
timestamp 1704896540
transform 1 0 6144 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_27_55
timestamp 1704896540
transform 1 0 6432 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_27_63
timestamp 1704896540
transform 1 0 7200 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_27_67
timestamp 1704896540
transform 1 0 7584 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_27_92
timestamp 1704896540
transform 1 0 9984 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_28_52
timestamp 1704896540
transform 1 0 6144 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_28_60
timestamp 1704896540
transform 1 0 6912 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_28_68
timestamp 1704896540
transform 1 0 7680 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_28_76
timestamp 1704896540
transform 1 0 8448 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_28_80
timestamp 1704896540
transform 1 0 8832 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_28_82
timestamp 1704896540
transform 1 0 9024 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_28_90
timestamp 1704896540
transform 1 0 9792 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_29_8
timestamp 1704896540
transform 1 0 1920 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_29_16
timestamp 1704896540
transform 1 0 2688 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_29_24
timestamp 1704896540
transform 1 0 3456 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_29_32
timestamp 1704896540
transform 1 0 4224 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_29_40
timestamp 1704896540
transform 1 0 4992 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_29_48
timestamp 1704896540
transform 1 0 5760 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_29_52
timestamp 1704896540
transform 1 0 6144 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_29_55
timestamp 1704896540
transform 1 0 6432 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_29_63
timestamp 1704896540
transform 1 0 7200 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_29_67
timestamp 1704896540
transform 1 0 7584 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_29_92
timestamp 1704896540
transform 1 0 9984 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_30_4
timestamp 1704896540
transform 1 0 1536 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_30_12
timestamp 1704896540
transform 1 0 2304 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_30_20
timestamp 1704896540
transform 1 0 3072 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_30_24
timestamp 1704896540
transform 1 0 3456 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_30_26
timestamp 1704896540
transform 1 0 3648 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_30_28
timestamp 1704896540
transform 1 0 3840 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_30_36
timestamp 1704896540
transform 1 0 4608 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_30_44
timestamp 1704896540
transform 1 0 5376 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_30_69
timestamp 1704896540
transform 1 0 7776 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_30_75
timestamp 1704896540
transform 1 0 8352 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_30_79
timestamp 1704896540
transform 1 0 8736 0 1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_30_82
timestamp 1704896540
transform 1 0 9024 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_31_8
timestamp 1704896540
transform 1 0 1920 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_31_16
timestamp 1704896540
transform 1 0 2688 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_31_24
timestamp 1704896540
transform 1 0 3456 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_31_32
timestamp 1704896540
transform 1 0 4224 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_31_40
timestamp 1704896540
transform 1 0 4992 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_31_48
timestamp 1704896540
transform 1 0 5760 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_31_52
timestamp 1704896540
transform 1 0 6144 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_31_78
timestamp 1704896540
transform 1 0 8640 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_31_83
timestamp 1704896540
transform 1 0 9120 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_31_91
timestamp 1704896540
transform 1 0 9888 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_31_93
timestamp 1704896540
transform 1 0 10080 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_4
timestamp 1704896540
transform 1 0 1536 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_12
timestamp 1704896540
transform 1 0 2304 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_32_20
timestamp 1704896540
transform 1 0 3072 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_32_24
timestamp 1704896540
transform 1 0 3456 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_32_26
timestamp 1704896540
transform 1 0 3648 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_28
timestamp 1704896540
transform 1 0 3840 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_36
timestamp 1704896540
transform 1 0 4608 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_44
timestamp 1704896540
transform 1 0 5376 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_52
timestamp 1704896540
transform 1 0 6144 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_60
timestamp 1704896540
transform 1 0 6912 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_68
timestamp 1704896540
transform 1 0 7680 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_32_76
timestamp 1704896540
transform 1 0 8448 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_32_80
timestamp 1704896540
transform 1 0 8832 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_82
timestamp 1704896540
transform 1 0 9024 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_32_90
timestamp 1704896540
transform 1 0 9792 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_12
timestamp 1704896540
transform 1 0 2304 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_20
timestamp 1704896540
transform 1 0 3072 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_28
timestamp 1704896540
transform 1 0 3840 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_36
timestamp 1704896540
transform 1 0 4608 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_44
timestamp 1704896540
transform 1 0 5376 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_33_52
timestamp 1704896540
transform 1 0 6144 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_55
timestamp 1704896540
transform 1 0 6432 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_63
timestamp 1704896540
transform 1 0 7200 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_71
timestamp 1704896540
transform 1 0 7968 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_79
timestamp 1704896540
transform 1 0 8736 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_33_87
timestamp 1704896540
transform 1 0 9504 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_33_89
timestamp 1704896540
transform 1 0 9696 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_4
timestamp 1704896540
transform 1 0 1536 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_34_6
timestamp 1704896540
transform 1 0 1728 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_34_15
timestamp 1704896540
transform 1 0 2592 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  FILLER_0_34_23
timestamp 1704896540
transform 1 0 3360 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_28
timestamp 1704896540
transform 1 0 3840 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_34_30
timestamp 1704896540
transform 1 0 4032 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_34_35
timestamp 1704896540
transform 1 0 4512 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_34_47
timestamp 1704896540
transform 1 0 5664 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_51
timestamp 1704896540
transform 1 0 6048 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_34_53
timestamp 1704896540
transform 1 0 6240 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_34_59
timestamp 1704896540
transform 1 0 6816 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_34_71
timestamp 1704896540
transform 1 0 7968 0 1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_79
timestamp 1704896540
transform 1 0 8736 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__clkbuf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 1920 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  input2
timestamp 1704896540
transform -1 0 1920 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__buf_8  input3 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 1536 0 -1 3996
box -38 -49 1190 715
use sky130_fd_sc_hs__clkbuf_4  input4 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 2112 0 1 7992
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_1  output5
timestamp 1704896540
transform -1 0 1920 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output6
timestamp 1704896540
transform -1 0 1920 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output7
timestamp 1704896540
transform -1 0 1920 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output8
timestamp 1704896540
transform -1 0 1920 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output9
timestamp 1704896540
transform -1 0 1920 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output10
timestamp 1704896540
transform -1 0 1920 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output11
timestamp 1704896540
transform -1 0 1920 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output12
timestamp 1704896540
transform -1 0 1920 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output13
timestamp 1704896540
transform -1 0 1920 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output14
timestamp 1704896540
transform -1 0 1920 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output15
timestamp 1704896540
transform 1 0 9408 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output16
timestamp 1704896540
transform -1 0 2592 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output17
timestamp 1704896540
transform -1 0 2592 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output18
timestamp 1704896540
transform 1 0 9408 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output19
timestamp 1704896540
transform 1 0 9792 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output20
timestamp 1704896540
transform 1 0 9792 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output21
timestamp 1704896540
transform 1 0 9792 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output22
timestamp 1704896540
transform 1 0 9792 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output23
timestamp 1704896540
transform 1 0 9792 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output24
timestamp 1704896540
transform 1 0 9792 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output25
timestamp 1704896540
transform 1 0 9792 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output26
timestamp 1704896540
transform 1 0 9792 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output27
timestamp 1704896540
transform 1 0 9792 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output28
timestamp 1704896540
transform -1 0 2976 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output29
timestamp 1704896540
transform -1 0 2208 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output30
timestamp 1704896540
transform -1 0 3360 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output31
timestamp 1704896540
transform -1 0 4512 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output32
timestamp 1704896540
transform -1 0 5664 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output33
timestamp 1704896540
transform -1 0 6816 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output34
timestamp 1704896540
transform -1 0 8544 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output35
timestamp 1704896540
transform -1 0 9408 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output36
timestamp 1704896540
transform -1 0 10176 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output37
timestamp 1704896540
transform 1 0 9408 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output38
timestamp 1704896540
transform -1 0 2304 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output39
timestamp 1704896540
transform -1 0 2208 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output40
timestamp 1704896540
transform -1 0 3360 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output41
timestamp 1704896540
transform -1 0 4512 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output42
timestamp 1704896540
transform -1 0 5664 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output43
timestamp 1704896540
transform -1 0 6816 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output44
timestamp 1704896540
transform -1 0 7968 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output45
timestamp 1704896540
transform -1 0 9408 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output46
timestamp 1704896540
transform -1 0 10176 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output47
timestamp 1704896540
transform 1 0 9792 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_0_Left_35
timestamp 1704896540
transform 1 0 1152 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 10560 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_1_Left_36
timestamp 1704896540
transform 1 0 1152 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 10560 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_2_Left_37
timestamp 1704896540
transform 1 0 1152 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 10560 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_3_Left_38
timestamp 1704896540
transform 1 0 1152 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 10560 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_4_Left_39
timestamp 1704896540
transform 1 0 1152 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 10560 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_5_Left_40
timestamp 1704896540
transform 1 0 1152 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 10560 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_6_Left_41
timestamp 1704896540
transform 1 0 1152 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 10560 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_7_Left_42
timestamp 1704896540
transform 1 0 1152 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 10560 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_8_Left_43
timestamp 1704896540
transform 1 0 1152 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 10560 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_9_Left_44
timestamp 1704896540
transform 1 0 1152 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 10560 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_10_Left_45
timestamp 1704896540
transform 1 0 1152 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 10560 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_11_Left_46
timestamp 1704896540
transform 1 0 1152 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 10560 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_12_Left_47
timestamp 1704896540
transform 1 0 1152 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 10560 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_13_Left_48
timestamp 1704896540
transform 1 0 1152 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 10560 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_14_Left_49
timestamp 1704896540
transform 1 0 1152 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 10560 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_15_Left_50
timestamp 1704896540
transform 1 0 1152 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 10560 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_16_Left_51
timestamp 1704896540
transform 1 0 1152 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 10560 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_17_Left_52
timestamp 1704896540
transform 1 0 1152 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 10560 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_18_Left_53
timestamp 1704896540
transform 1 0 1152 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 10560 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_19_Left_54
timestamp 1704896540
transform 1 0 1152 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 10560 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_20_Left_55
timestamp 1704896540
transform 1 0 1152 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 10560 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_21_Left_56
timestamp 1704896540
transform 1 0 1152 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 10560 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_22_Left_57
timestamp 1704896540
transform 1 0 1152 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 10560 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_23_Left_58
timestamp 1704896540
transform 1 0 1152 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 10560 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_24_Left_59
timestamp 1704896540
transform 1 0 1152 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 10560 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_25_Left_60
timestamp 1704896540
transform 1 0 1152 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 10560 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_26_Left_61
timestamp 1704896540
transform 1 0 1152 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 10560 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_27_Left_62
timestamp 1704896540
transform 1 0 1152 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 10560 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_28_Left_63
timestamp 1704896540
transform 1 0 1152 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 10560 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_29_Left_64
timestamp 1704896540
transform 1 0 1152 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_29_Right_29
timestamp 1704896540
transform -1 0 10560 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_30_Left_65
timestamp 1704896540
transform 1 0 1152 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_30_Right_30
timestamp 1704896540
transform -1 0 10560 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_31_Left_66
timestamp 1704896540
transform 1 0 1152 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_31_Right_31
timestamp 1704896540
transform -1 0 10560 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_32_Left_67
timestamp 1704896540
transform 1 0 1152 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_32_Right_32
timestamp 1704896540
transform -1 0 10560 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_33_Left_68
timestamp 1704896540
transform 1 0 1152 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_33_Right_33
timestamp 1704896540
transform -1 0 10560 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_34_Left_69
timestamp 1704896540
transform 1 0 1152 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_34_Right_34
timestamp 1704896540
transform -1 0 10560 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749010377
transform 1 0 3744 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1749010377
transform 1 0 6336 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1749010377
transform 1 0 8928 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_73
timestamp 1749010377
transform 1 0 6336 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_74
timestamp 1749010377
transform 1 0 3744 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_75
timestamp 1749010377
transform 1 0 8928 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_76
timestamp 1749010377
transform 1 0 6336 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_77
timestamp 1749010377
transform 1 0 3744 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_78
timestamp 1749010377
transform 1 0 8928 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_79
timestamp 1749010377
transform 1 0 6336 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_80
timestamp 1749010377
transform 1 0 3744 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_81
timestamp 1749010377
transform 1 0 8928 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp 1749010377
transform 1 0 6336 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp 1749010377
transform 1 0 3744 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_84
timestamp 1749010377
transform 1 0 8928 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_85
timestamp 1749010377
transform 1 0 6336 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_86
timestamp 1749010377
transform 1 0 3744 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_87
timestamp 1749010377
transform 1 0 8928 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_88
timestamp 1749010377
transform 1 0 6336 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_89
timestamp 1749010377
transform 1 0 3744 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_90
timestamp 1749010377
transform 1 0 8928 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_91
timestamp 1749010377
transform 1 0 6336 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_92
timestamp 1749010377
transform 1 0 3744 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_93
timestamp 1749010377
transform 1 0 8928 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_94
timestamp 1749010377
transform 1 0 6336 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_95
timestamp 1749010377
transform 1 0 3744 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_96
timestamp 1749010377
transform 1 0 8928 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_97
timestamp 1749010377
transform 1 0 6336 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_98
timestamp 1749010377
transform 1 0 3744 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_99
timestamp 1749010377
transform 1 0 8928 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_100
timestamp 1749010377
transform 1 0 6336 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_101
timestamp 1749010377
transform 1 0 3744 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_102
timestamp 1749010377
transform 1 0 8928 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_103
timestamp 1749010377
transform 1 0 6336 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_104
timestamp 1749010377
transform 1 0 3744 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_105
timestamp 1749010377
transform 1 0 8928 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_106
timestamp 1749010377
transform 1 0 6336 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_107
timestamp 1749010377
transform 1 0 3744 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_108
timestamp 1749010377
transform 1 0 8928 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_109
timestamp 1749010377
transform 1 0 6336 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_110
timestamp 1749010377
transform 1 0 3744 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_111
timestamp 1749010377
transform 1 0 8928 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_112
timestamp 1749010377
transform 1 0 6336 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_113
timestamp 1749010377
transform 1 0 3744 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_114
timestamp 1749010377
transform 1 0 8928 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_115
timestamp 1749010377
transform 1 0 6336 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_116
timestamp 1749010377
transform 1 0 3744 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_117
timestamp 1749010377
transform 1 0 8928 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_118
timestamp 1749010377
transform 1 0 6336 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_119
timestamp 1749010377
transform 1 0 3744 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_120
timestamp 1749010377
transform 1 0 8928 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_121
timestamp 1749010377
transform 1 0 6336 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_122
timestamp 1749010377
transform 1 0 3744 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_123
timestamp 1749010377
transform 1 0 6336 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_124
timestamp 1749010377
transform 1 0 8928 0 1 25308
box -38 -49 134 715
<< labels >>
flabel metal3 s 0 9782 800 9902 0 FreeSans 480 0 0 0 CF[0]
port 0 nsew signal output
flabel metal3 s 0 11262 800 11382 0 FreeSans 480 0 0 0 CF[1]
port 1 nsew signal output
flabel metal3 s 0 12742 800 12862 0 FreeSans 480 0 0 0 CF[2]
port 2 nsew signal output
flabel metal3 s 0 14222 800 14342 0 FreeSans 480 0 0 0 CF[3]
port 3 nsew signal output
flabel metal3 s 0 15702 800 15822 0 FreeSans 480 0 0 0 CF[4]
port 4 nsew signal output
flabel metal3 s 0 17182 800 17302 0 FreeSans 480 0 0 0 CF[5]
port 5 nsew signal output
flabel metal3 s 0 18662 800 18782 0 FreeSans 480 0 0 0 CF[6]
port 6 nsew signal output
flabel metal3 s 0 20142 800 20262 0 FreeSans 480 0 0 0 CF[7]
port 7 nsew signal output
flabel metal3 s 0 21622 800 21742 0 FreeSans 480 0 0 0 CF[8]
port 8 nsew signal output
flabel metal3 s 0 23102 800 23222 0 FreeSans 480 0 0 0 CF[9]
port 9 nsew signal output
flabel metal3 s 10922 27246 11722 27366 0 FreeSans 480 0 0 0 CKO
port 10 nsew signal output
flabel metal3 s 0 26062 800 26182 0 FreeSans 480 0 0 0 CKS
port 11 nsew signal output
flabel metal3 s 0 2382 800 2502 0 FreeSans 480 0 0 0 CKSB
port 12 nsew signal output
flabel metal3 s 0 5342 800 5462 0 FreeSans 480 0 0 0 CLK
port 13 nsew signal input
flabel metal3 s 0 8302 800 8422 0 FreeSans 480 0 0 0 CMP_N
port 14 nsew signal input
flabel metal3 s 0 24582 800 24702 0 FreeSans 480 0 0 0 CMP_P
port 15 nsew signal input
flabel metal3 s 10922 1198 11722 1318 0 FreeSans 480 0 0 0 DATA[0]
port 16 nsew signal output
flabel metal3 s 10922 3566 11722 3686 0 FreeSans 480 0 0 0 DATA[1]
port 17 nsew signal output
flabel metal3 s 10922 5934 11722 6054 0 FreeSans 480 0 0 0 DATA[2]
port 18 nsew signal output
flabel metal3 s 10922 8302 11722 8422 0 FreeSans 480 0 0 0 DATA[3]
port 19 nsew signal output
flabel metal3 s 10922 10670 11722 10790 0 FreeSans 480 0 0 0 DATA[4]
port 20 nsew signal output
flabel metal3 s 10922 13038 11722 13158 0 FreeSans 480 0 0 0 DATA[5]
port 21 nsew signal output
flabel metal3 s 10922 15406 11722 15526 0 FreeSans 480 0 0 0 DATA[6]
port 22 nsew signal output
flabel metal3 s 10922 17774 11722 17894 0 FreeSans 480 0 0 0 DATA[7]
port 23 nsew signal output
flabel metal3 s 10922 20142 11722 20262 0 FreeSans 480 0 0 0 DATA[8]
port 24 nsew signal output
flabel metal3 s 10922 22510 11722 22630 0 FreeSans 480 0 0 0 DATA[9]
port 25 nsew signal output
flabel metal3 s 0 3862 800 3982 0 FreeSans 480 0 0 0 EN
port 26 nsew signal input
flabel metal3 s 0 6822 800 6942 0 FreeSans 480 0 0 0 RDY
port 27 nsew signal input
flabel metal2 s 596 0 652 800 0 FreeSans 224 90 0 0 SWN[0]
port 28 nsew signal output
flabel metal2 s 1748 0 1804 800 0 FreeSans 224 90 0 0 SWN[1]
port 29 nsew signal output
flabel metal2 s 2900 0 2956 800 0 FreeSans 224 90 0 0 SWN[2]
port 30 nsew signal output
flabel metal2 s 4052 0 4108 800 0 FreeSans 224 90 0 0 SWN[3]
port 31 nsew signal output
flabel metal2 s 5204 0 5260 800 0 FreeSans 224 90 0 0 SWN[4]
port 32 nsew signal output
flabel metal2 s 6356 0 6412 800 0 FreeSans 224 90 0 0 SWN[5]
port 33 nsew signal output
flabel metal2 s 7508 0 7564 800 0 FreeSans 224 90 0 0 SWN[6]
port 34 nsew signal output
flabel metal2 s 8660 0 8716 800 0 FreeSans 224 90 0 0 SWN[7]
port 35 nsew signal output
flabel metal2 s 9812 0 9868 800 0 FreeSans 224 90 0 0 SWN[8]
port 36 nsew signal output
flabel metal2 s 10964 0 11020 800 0 FreeSans 224 90 0 0 SWN[9]
port 37 nsew signal output
flabel metal2 s 596 28074 652 28874 0 FreeSans 224 90 0 0 SWP[0]
port 38 nsew signal output
flabel metal2 s 1748 28074 1804 28874 0 FreeSans 224 90 0 0 SWP[1]
port 39 nsew signal output
flabel metal2 s 2900 28074 2956 28874 0 FreeSans 224 90 0 0 SWP[2]
port 40 nsew signal output
flabel metal2 s 4052 28074 4108 28874 0 FreeSans 224 90 0 0 SWP[3]
port 41 nsew signal output
flabel metal2 s 5204 28074 5260 28874 0 FreeSans 224 90 0 0 SWP[4]
port 42 nsew signal output
flabel metal2 s 6356 28074 6412 28874 0 FreeSans 224 90 0 0 SWP[5]
port 43 nsew signal output
flabel metal2 s 7508 28074 7564 28874 0 FreeSans 224 90 0 0 SWP[6]
port 44 nsew signal output
flabel metal2 s 8660 28074 8716 28874 0 FreeSans 224 90 0 0 SWP[7]
port 45 nsew signal output
flabel metal2 s 9812 28074 9868 28874 0 FreeSans 224 90 0 0 SWP[8]
port 46 nsew signal output
flabel metal2 s 10964 28074 11020 28874 0 FreeSans 224 90 0 0 SWP[9]
port 47 nsew signal output
flabel metal4 s 4952 2616 5352 26022 0 FreeSans 1920 90 0 0 VGND
port 48 nsew ground bidirectional
flabel metal4 s 1952 2616 2352 26022 0 FreeSans 1920 90 0 0 VPWR
port 49 nsew power bidirectional
flabel metal4 s 7952 2616 8352 26022 0 FreeSans 1920 90 0 0 VPWR
port 49 nsew power bidirectional
rlabel metal1 5856 25308 5856 25308 0 VGND
rlabel metal1 5856 25974 5856 25974 0 VPWR
rlabel metal3 1143 9842 1143 9842 0 CF[0]
rlabel metal3 1143 11322 1143 11322 0 CF[1]
rlabel metal3 1143 12802 1143 12802 0 CF[2]
rlabel metal3 759 14282 759 14282 0 CF[3]
rlabel metal3 759 15762 759 15762 0 CF[4]
rlabel metal1 1440 17205 1440 17205 0 CF[5]
rlabel metal2 1584 18629 1584 18629 0 CF[6]
rlabel metal2 1584 20035 1584 20035 0 CF[7]
rlabel metal3 807 21682 807 21682 0 CF[8]
rlabel metal3 759 23162 759 23162 0 CF[9]
rlabel metal2 9744 26584 9744 26584 0 CKO
rlabel metal1 1968 25789 1968 25789 0 CKS
rlabel metal3 1479 2442 1479 2442 0 CKSB
rlabel metal3 1935 5402 1935 5402 0 CLK
rlabel metal3 1191 8362 1191 8362 0 CMP_N
rlabel metal3 807 24642 807 24642 0 CMP_P
rlabel metal2 9744 2090 9744 2090 0 DATA[0]
rlabel via2 10128 3607 10128 3607 0 DATA[1]
rlabel metal2 10128 6049 10128 6049 0 DATA[2]
rlabel via2 10128 8343 10128 8343 0 DATA[3]
rlabel via2 10128 10748 10128 10748 0 DATA[4]
rlabel metal2 10128 13264 10128 13264 0 DATA[5]
rlabel via2 10128 15447 10128 15447 0 DATA[6]
rlabel via2 10128 17815 10128 17815 0 DATA[7]
rlabel via2 10128 20183 10128 20183 0 DATA[8]
rlabel metal2 10128 22662 10128 22662 0 DATA[9]
rlabel metal3 807 3922 807 3922 0 EN
rlabel metal3 1191 6882 1191 6882 0 RDY
rlabel metal2 624 1875 624 1875 0 SWN[0]
rlabel metal2 1831 666 1831 666 0 SWN[1]
rlabel metal2 2983 666 2983 666 0 SWN[2]
rlabel metal2 4135 666 4135 666 0 SWN[3]
rlabel metal2 5335 666 5335 666 0 SWN[4]
rlabel metal2 6439 666 6439 666 0 SWN[5]
rlabel metal2 7536 2097 7536 2097 0 SWN[6]
rlabel metal2 8791 666 8791 666 0 SWN[7]
rlabel metal2 9840 1801 9840 1801 0 SWN[8]
rlabel metal2 10992 2060 10992 2060 0 SWN[9]
rlabel metal1 1296 25197 1296 25197 0 SWP[0]
rlabel metal1 1824 25863 1824 25863 0 SWP[1]
rlabel metal2 2983 28194 2983 28194 0 SWP[2]
rlabel metal2 4135 28194 4135 28194 0 SWP[3]
rlabel metal2 5287 28194 5287 28194 0 SWP[4]
rlabel metal2 6439 28194 6439 28194 0 SWP[5]
rlabel metal2 7591 28194 7591 28194 0 SWP[6]
rlabel metal1 8880 25863 8880 25863 0 SWP[7]
rlabel metal2 9840 27021 9840 27021 0 SWP[8]
rlabel metal1 10560 25197 10560 25197 0 SWP[9]
rlabel metal1 6000 4551 6000 4551 0 _00_
rlabel metal2 6864 5587 6864 5587 0 _01_
rlabel metal1 6672 3737 6672 3737 0 _02_
rlabel metal2 8592 5254 8592 5254 0 _03_
rlabel metal1 7080 6253 7080 6253 0 _04_
rlabel metal1 6768 7067 6768 7067 0 _05_
rlabel metal1 8544 22829 8544 22829 0 _06_
rlabel metal1 5856 5661 5856 5661 0 _07_
rlabel metal1 5808 4366 5808 4366 0 _08_
rlabel metal1 5904 5439 5904 5439 0 _09_
rlabel metal1 6096 6549 6096 6549 0 _10_
rlabel metal1 5328 6290 5328 6290 0 _11_
rlabel metal2 8496 4514 8496 4514 0 _12_
rlabel metal1 9024 4181 9024 4181 0 _13_
rlabel metal2 9552 6364 9552 6364 0 _14_
rlabel metal1 9504 5217 9504 5217 0 _15_
rlabel metal1 8304 7215 8304 7215 0 _16_
rlabel metal1 7152 7622 7152 7622 0 _17_
rlabel metal1 6480 4255 6480 4255 0 clk_div_0.COUNT\[0\]
rlabel metal1 8736 5069 8736 5069 0 clk_div_0.COUNT\[1\]
rlabel metal1 9024 6327 9024 6327 0 clk_div_0.COUNT\[2\]
rlabel metal1 8307 6919 8307 6919 0 clk_div_0.COUNT\[3\]
rlabel metal2 7152 3663 7152 3663 0 clknet_0_CLK
rlabel metal2 6576 3367 6576 3367 0 clknet_1_0__leaf_CLK
rlabel metal1 6528 6327 6528 6327 0 clknet_1_1__leaf_CLK
rlabel metal1 8064 18315 8064 18315 0 cyclic_flag_0.FINAL
rlabel metal1 2256 5587 2256 5587 0 net1
rlabel via1 4272 17649 4272 17649 0 net10
rlabel metal1 4560 18981 4560 18981 0 net11
rlabel metal1 5856 20313 5856 20313 0 net12
rlabel metal1 6000 22940 6000 22940 0 net13
rlabel metal1 6816 23643 6816 23643 0 net14
rlabel metal1 9264 23865 9264 23865 0 net15
rlabel metal1 5616 5587 5616 5587 0 net16
rlabel metal2 4656 3922 4656 3922 0 net17
rlabel metal1 9792 2997 9792 2997 0 net18
rlabel metal1 9792 3663 9792 3663 0 net19
rlabel metal2 5616 23939 5616 23939 0 net2
rlabel metal1 9792 10101 9792 10101 0 net20
rlabel metal1 9696 8325 9696 8325 0 net21
rlabel metal2 9840 13209 9840 13209 0 net22
rlabel metal1 9792 13653 9792 13653 0 net23
rlabel metal2 9840 16206 9840 16206 0 net24
rlabel metal2 9840 18537 9840 18537 0 net25
rlabel metal2 9840 20535 9840 20535 0 net26
rlabel metal2 9840 22755 9840 22755 0 net27
rlabel metal2 2928 4218 2928 4218 0 net28
rlabel metal1 1872 2997 1872 2997 0 net29
rlabel metal1 6192 3848 6192 3848 0 net3
rlabel metal2 3312 3885 3312 3885 0 net30
rlabel metal1 5184 10767 5184 10767 0 net31
rlabel metal1 5280 12987 5280 12987 0 net32
rlabel metal1 6912 2997 6912 2997 0 net33
rlabel metal1 7968 3663 7968 3663 0 net34
rlabel metal2 8208 6438 8208 6438 0 net35
rlabel metal1 10176 2997 10176 2997 0 net36
rlabel metal1 8880 10767 8880 10767 0 net37
rlabel metal1 2400 24975 2400 24975 0 net38
rlabel metal1 2448 25567 2448 25567 0 net39
rlabel metal1 3072 6993 3072 6993 0 net4
rlabel metal1 3792 11877 3792 11877 0 net40
rlabel metal1 5088 25567 5088 25567 0 net41
rlabel metal2 5616 16243 5616 16243 0 net42
rlabel metal2 6480 21756 6480 21756 0 net43
rlabel metal2 7824 22200 7824 22200 0 net44
rlabel metal1 7680 20535 7680 20535 0 net45
rlabel metal2 7632 24272 7632 24272 0 net46
rlabel metal2 8496 24420 8496 24420 0 net47
rlabel metal1 1584 5698 1584 5698 0 net5
rlabel metal2 3792 5291 3792 5291 0 net6
rlabel metal1 1968 4995 1968 4995 0 net7
rlabel metal1 3936 12099 3936 12099 0 net8
rlabel metal1 2544 14763 2544 14763 0 net9
<< properties >>
string FIXED_BBOX 0 0 11722 28874
<< end >>
