magic
tech sky130A
magscale 1 2
timestamp 1749385379
<< locali >>
rect 628 2103 659 2137
rect 693 2103 755 2137
rect 789 2103 851 2137
rect 885 2103 947 2137
rect 981 2103 1043 2137
rect 1077 2103 1139 2137
rect 1173 2103 1235 2137
rect 1269 2103 1331 2137
rect 1365 2103 1427 2137
rect 1461 2103 1523 2137
rect 1557 2103 1619 2137
rect 1653 2103 1682 2137
rect 664 1947 698 2103
rect 980 1956 1014 2103
rect 1296 1959 1330 2103
rect 1612 1958 1646 2103
rect 664 -2317 698 -2167
rect 980 -2317 1014 -2169
rect 1296 -2317 1330 -2176
rect 1612 -2317 1646 -2163
rect 628 -2351 659 -2317
rect 693 -2351 755 -2317
rect 789 -2351 851 -2317
rect 885 -2351 947 -2317
rect 981 -2351 1043 -2317
rect 1077 -2351 1139 -2317
rect 1173 -2351 1235 -2317
rect 1269 -2351 1331 -2317
rect 1365 -2351 1427 -2317
rect 1461 -2351 1523 -2317
rect 1557 -2351 1619 -2317
rect 1653 -2351 1682 -2317
<< viali >>
rect 659 2103 693 2137
rect 755 2103 789 2137
rect 851 2103 885 2137
rect 947 2103 981 2137
rect 1043 2103 1077 2137
rect 1139 2103 1173 2137
rect 1235 2103 1269 2137
rect 1331 2103 1365 2137
rect 1427 2103 1461 2137
rect 1523 2103 1557 2137
rect 1619 2103 1653 2137
rect 659 -2351 693 -2317
rect 755 -2351 789 -2317
rect 851 -2351 885 -2317
rect 947 -2351 981 -2317
rect 1043 -2351 1077 -2317
rect 1139 -2351 1173 -2317
rect 1235 -2351 1269 -2317
rect 1331 -2351 1365 -2317
rect 1427 -2351 1461 -2317
rect 1523 -2351 1557 -2317
rect 1619 -2351 1653 -2317
<< metal1 >>
rect 628 2137 1682 2168
rect 628 2103 659 2137
rect 693 2103 755 2137
rect 789 2103 851 2137
rect 885 2103 947 2137
rect 981 2103 1043 2137
rect 1077 2103 1139 2137
rect 1173 2103 1235 2137
rect 1269 2103 1331 2137
rect 1365 2103 1427 2137
rect 1461 2103 1523 2137
rect 1557 2103 1619 2137
rect 1653 2103 1682 2137
rect 628 2072 1682 2103
rect 803 1980 813 2032
rect 865 1980 1445 2032
rect 1497 1980 1507 2032
rect 803 1894 813 1946
rect 865 1894 875 1946
rect 1119 1894 1129 1946
rect 1181 1894 1191 1946
rect 1435 1894 1445 1946
rect 1497 1894 1507 1946
rect 584 -2126 1094 1850
rect 1216 -2126 1726 1850
rect 628 -2317 1682 -2286
rect 628 -2351 659 -2317
rect 693 -2351 755 -2317
rect 789 -2351 851 -2317
rect 885 -2351 947 -2317
rect 981 -2351 1043 -2317
rect 1077 -2351 1139 -2317
rect 1173 -2351 1235 -2317
rect 1269 -2351 1331 -2317
rect 1365 -2351 1427 -2317
rect 1461 -2351 1523 -2317
rect 1557 -2351 1619 -2317
rect 1653 -2351 1682 -2317
rect 628 -2382 1682 -2351
<< via1 >>
rect 813 1980 865 2032
rect 1445 1980 1497 2032
rect 813 1894 865 1946
rect 1129 1894 1181 1946
rect 1445 1894 1497 1946
<< metal2 >>
rect 813 2032 865 2168
rect 813 1946 865 1980
rect 813 1884 865 1894
rect 1129 1946 1181 2168
rect 1129 1884 1181 1894
rect 1445 2032 1497 2042
rect 1445 1946 1497 1980
rect 1445 1884 1497 1894
use sky130_fd_pr__nfet_01v8_9HAEJX  XM10
timestamp 1749384884
transform 1 0 839 0 1 -107
box -211 -2179 211 2179
use sky130_fd_pr__nfet_01v8_WBAE2P  XM11
timestamp 1749384884
transform 1 0 1155 0 1 -107
box -211 -2179 211 2179
use sky130_fd_pr__nfet_01v8_9HAEH6  XM12
timestamp 1749384884
transform 1 0 1471 0 1 -107
box -211 -2179 211 2179
<< labels >>
flabel metal2 813 2116 865 2168 0 FreeSans 400 0 0 0 CK
port 0 nsew
flabel metal2 1129 2114 1181 2166 0 FreeSans 400 0 0 0 VGS
port 1 nsew
flabel viali 659 2103 693 2137 0 FreeSans 400 0 0 0 VSS
port 2 nsew
flabel metal1 1692 1816 1726 1850 0 FreeSans 400 0 0 0 IN
port 3 nsew
flabel metal1 584 1816 618 1850 0 FreeSans 400 0 0 0 OUT
port 4 nsew
<< end >>
