magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect 142 1527 172 1561
rect 206 1527 244 1561
rect 278 1527 316 1561
rect 350 1527 388 1561
rect 422 1527 460 1561
rect 494 1527 532 1561
rect 566 1527 604 1561
rect 638 1527 676 1561
rect 710 1527 748 1561
rect 782 1527 820 1561
rect 854 1527 892 1561
rect 926 1527 964 1561
rect 998 1527 1036 1561
rect 1070 1527 1108 1561
rect 1142 1527 1180 1561
rect 1214 1527 1252 1561
rect 1286 1527 1324 1561
rect 1358 1527 1396 1561
rect 1430 1527 1468 1561
rect 1502 1527 1540 1561
rect 1574 1527 1612 1561
rect 1646 1527 1684 1561
rect 1718 1527 1756 1561
rect 1790 1527 1828 1561
rect 1862 1527 1900 1561
rect 1934 1527 1972 1561
rect 2006 1527 2044 1561
rect 2078 1527 2116 1561
rect 2150 1527 2188 1561
rect 2222 1527 2260 1561
rect 2294 1527 2332 1561
rect 2366 1527 2404 1561
rect 2438 1527 2476 1561
rect 2510 1527 2548 1561
rect 2582 1527 2620 1561
rect 2654 1527 2692 1561
rect 2726 1527 2764 1561
rect 2798 1527 2836 1561
rect 2870 1527 2908 1561
rect 2942 1527 2980 1561
rect 3014 1527 3052 1561
rect 3086 1527 3124 1561
rect 3158 1527 3196 1561
rect 3230 1527 3268 1561
rect 3302 1527 3340 1561
rect 3374 1527 3412 1561
rect 3446 1527 3484 1561
rect 3518 1527 3556 1561
rect 3590 1527 3628 1561
rect 3662 1527 3700 1561
rect 3734 1527 3772 1561
rect 3806 1527 3844 1561
rect 3878 1527 3916 1561
rect 3950 1527 3988 1561
rect 4022 1527 4060 1561
rect 4094 1527 4132 1561
rect 4166 1527 4204 1561
rect 4238 1527 4276 1561
rect 4310 1527 4348 1561
rect 4382 1527 4420 1561
rect 4454 1527 4492 1561
rect 4526 1527 4564 1561
rect 4598 1527 4636 1561
rect 4670 1527 4708 1561
rect 4742 1527 4780 1561
rect 4814 1527 4852 1561
rect 4886 1527 4924 1561
rect 4958 1527 4996 1561
rect 5030 1527 5068 1561
rect 5102 1527 5140 1561
rect 5174 1527 5212 1561
rect 5246 1527 5284 1561
rect 5318 1527 5356 1561
rect 5390 1527 5428 1561
rect 5462 1527 5500 1561
rect 5534 1527 5572 1561
rect 5606 1527 5644 1561
rect 5678 1527 5716 1561
rect 5750 1527 5788 1561
rect 5822 1527 5860 1561
rect 5894 1527 5932 1561
rect 5966 1527 6004 1561
rect 6038 1527 6076 1561
rect 6110 1527 6148 1561
rect 6182 1527 6220 1561
rect 6254 1527 6292 1561
rect 6326 1527 6364 1561
rect 6398 1527 6436 1561
rect 6470 1527 6508 1561
rect 6542 1527 6580 1561
rect 6614 1527 6652 1561
rect 6686 1527 6724 1561
rect 6758 1527 6796 1561
rect 6830 1527 6868 1561
rect 6902 1527 6940 1561
rect 6974 1527 7012 1561
rect 7046 1527 7084 1561
rect 7118 1527 7156 1561
rect 7190 1527 7228 1561
rect 7262 1527 7300 1561
rect 7334 1527 7372 1561
rect 7406 1527 7444 1561
rect 7478 1527 7516 1561
rect 7550 1527 7588 1561
rect 7622 1527 7660 1561
rect 7694 1527 7732 1561
rect 7766 1527 7804 1561
rect 7838 1527 7876 1561
rect 7910 1527 7948 1561
rect 7982 1527 8020 1561
rect 8054 1527 8084 1561
rect 142 -123 154 -89
rect 188 -123 226 -89
rect 260 -123 298 -89
rect 332 -123 370 -89
rect 404 -123 442 -89
rect 476 -123 514 -89
rect 548 -123 586 -89
rect 620 -123 658 -89
rect 692 -123 730 -89
rect 764 -123 802 -89
rect 836 -123 874 -89
rect 908 -123 946 -89
rect 980 -123 1018 -89
rect 1052 -123 1090 -89
rect 1124 -123 1162 -89
rect 1196 -123 1234 -89
rect 1268 -123 1306 -89
rect 1340 -123 1378 -89
rect 1412 -123 1450 -89
rect 1484 -123 1522 -89
rect 1556 -123 1594 -89
rect 1628 -123 1666 -89
rect 1700 -123 1738 -89
rect 1772 -123 1810 -89
rect 1844 -123 1882 -89
rect 1916 -123 1954 -89
rect 1988 -123 2026 -89
rect 2060 -123 2098 -89
rect 2132 -123 2170 -89
rect 2204 -123 2242 -89
rect 2276 -123 2314 -89
rect 2348 -123 2386 -89
rect 2420 -123 2458 -89
rect 2492 -123 2530 -89
rect 2564 -123 2602 -89
rect 2636 -123 2674 -89
rect 2708 -123 2746 -89
rect 2780 -123 2818 -89
rect 2852 -123 2890 -89
rect 2924 -123 2962 -89
rect 2996 -123 3034 -89
rect 3068 -123 3106 -89
rect 3140 -123 3178 -89
rect 3212 -123 3250 -89
rect 3284 -123 3322 -89
rect 3356 -123 3394 -89
rect 3428 -123 3466 -89
rect 3500 -123 3538 -89
rect 3572 -123 3610 -89
rect 3644 -123 3682 -89
rect 3716 -123 3754 -89
rect 3788 -123 3826 -89
rect 3860 -123 3898 -89
rect 3932 -123 3970 -89
rect 4004 -123 4042 -89
rect 4076 -123 4114 -89
rect 4148 -123 4160 -89
<< viali >>
rect 172 1527 206 1561
rect 244 1527 278 1561
rect 316 1527 350 1561
rect 388 1527 422 1561
rect 460 1527 494 1561
rect 532 1527 566 1561
rect 604 1527 638 1561
rect 676 1527 710 1561
rect 748 1527 782 1561
rect 820 1527 854 1561
rect 892 1527 926 1561
rect 964 1527 998 1561
rect 1036 1527 1070 1561
rect 1108 1527 1142 1561
rect 1180 1527 1214 1561
rect 1252 1527 1286 1561
rect 1324 1527 1358 1561
rect 1396 1527 1430 1561
rect 1468 1527 1502 1561
rect 1540 1527 1574 1561
rect 1612 1527 1646 1561
rect 1684 1527 1718 1561
rect 1756 1527 1790 1561
rect 1828 1527 1862 1561
rect 1900 1527 1934 1561
rect 1972 1527 2006 1561
rect 2044 1527 2078 1561
rect 2116 1527 2150 1561
rect 2188 1527 2222 1561
rect 2260 1527 2294 1561
rect 2332 1527 2366 1561
rect 2404 1527 2438 1561
rect 2476 1527 2510 1561
rect 2548 1527 2582 1561
rect 2620 1527 2654 1561
rect 2692 1527 2726 1561
rect 2764 1527 2798 1561
rect 2836 1527 2870 1561
rect 2908 1527 2942 1561
rect 2980 1527 3014 1561
rect 3052 1527 3086 1561
rect 3124 1527 3158 1561
rect 3196 1527 3230 1561
rect 3268 1527 3302 1561
rect 3340 1527 3374 1561
rect 3412 1527 3446 1561
rect 3484 1527 3518 1561
rect 3556 1527 3590 1561
rect 3628 1527 3662 1561
rect 3700 1527 3734 1561
rect 3772 1527 3806 1561
rect 3844 1527 3878 1561
rect 3916 1527 3950 1561
rect 3988 1527 4022 1561
rect 4060 1527 4094 1561
rect 4132 1527 4166 1561
rect 4204 1527 4238 1561
rect 4276 1527 4310 1561
rect 4348 1527 4382 1561
rect 4420 1527 4454 1561
rect 4492 1527 4526 1561
rect 4564 1527 4598 1561
rect 4636 1527 4670 1561
rect 4708 1527 4742 1561
rect 4780 1527 4814 1561
rect 4852 1527 4886 1561
rect 4924 1527 4958 1561
rect 4996 1527 5030 1561
rect 5068 1527 5102 1561
rect 5140 1527 5174 1561
rect 5212 1527 5246 1561
rect 5284 1527 5318 1561
rect 5356 1527 5390 1561
rect 5428 1527 5462 1561
rect 5500 1527 5534 1561
rect 5572 1527 5606 1561
rect 5644 1527 5678 1561
rect 5716 1527 5750 1561
rect 5788 1527 5822 1561
rect 5860 1527 5894 1561
rect 5932 1527 5966 1561
rect 6004 1527 6038 1561
rect 6076 1527 6110 1561
rect 6148 1527 6182 1561
rect 6220 1527 6254 1561
rect 6292 1527 6326 1561
rect 6364 1527 6398 1561
rect 6436 1527 6470 1561
rect 6508 1527 6542 1561
rect 6580 1527 6614 1561
rect 6652 1527 6686 1561
rect 6724 1527 6758 1561
rect 6796 1527 6830 1561
rect 6868 1527 6902 1561
rect 6940 1527 6974 1561
rect 7012 1527 7046 1561
rect 7084 1527 7118 1561
rect 7156 1527 7190 1561
rect 7228 1527 7262 1561
rect 7300 1527 7334 1561
rect 7372 1527 7406 1561
rect 7444 1527 7478 1561
rect 7516 1527 7550 1561
rect 7588 1527 7622 1561
rect 7660 1527 7694 1561
rect 7732 1527 7766 1561
rect 7804 1527 7838 1561
rect 7876 1527 7910 1561
rect 7948 1527 7982 1561
rect 8020 1527 8054 1561
rect 154 -123 188 -89
rect 226 -123 260 -89
rect 298 -123 332 -89
rect 370 -123 404 -89
rect 442 -123 476 -89
rect 514 -123 548 -89
rect 586 -123 620 -89
rect 658 -123 692 -89
rect 730 -123 764 -89
rect 802 -123 836 -89
rect 874 -123 908 -89
rect 946 -123 980 -89
rect 1018 -123 1052 -89
rect 1090 -123 1124 -89
rect 1162 -123 1196 -89
rect 1234 -123 1268 -89
rect 1306 -123 1340 -89
rect 1378 -123 1412 -89
rect 1450 -123 1484 -89
rect 1522 -123 1556 -89
rect 1594 -123 1628 -89
rect 1666 -123 1700 -89
rect 1738 -123 1772 -89
rect 1810 -123 1844 -89
rect 1882 -123 1916 -89
rect 1954 -123 1988 -89
rect 2026 -123 2060 -89
rect 2098 -123 2132 -89
rect 2170 -123 2204 -89
rect 2242 -123 2276 -89
rect 2314 -123 2348 -89
rect 2386 -123 2420 -89
rect 2458 -123 2492 -89
rect 2530 -123 2564 -89
rect 2602 -123 2636 -89
rect 2674 -123 2708 -89
rect 2746 -123 2780 -89
rect 2818 -123 2852 -89
rect 2890 -123 2924 -89
rect 2962 -123 2996 -89
rect 3034 -123 3068 -89
rect 3106 -123 3140 -89
rect 3178 -123 3212 -89
rect 3250 -123 3284 -89
rect 3322 -123 3356 -89
rect 3394 -123 3428 -89
rect 3466 -123 3500 -89
rect 3538 -123 3572 -89
rect 3610 -123 3644 -89
rect 3682 -123 3716 -89
rect 3754 -123 3788 -89
rect 3826 -123 3860 -89
rect 3898 -123 3932 -89
rect 3970 -123 4004 -89
rect 4042 -123 4076 -89
rect 4114 -123 4148 -89
<< metal1 >>
rect 106 1561 8120 1597
rect 106 1527 172 1561
rect 206 1527 244 1561
rect 278 1527 316 1561
rect 350 1527 388 1561
rect 422 1527 460 1561
rect 494 1527 532 1561
rect 566 1527 604 1561
rect 638 1527 676 1561
rect 710 1527 748 1561
rect 782 1527 820 1561
rect 854 1527 892 1561
rect 926 1527 964 1561
rect 998 1527 1036 1561
rect 1070 1527 1108 1561
rect 1142 1527 1180 1561
rect 1214 1527 1252 1561
rect 1286 1527 1324 1561
rect 1358 1527 1396 1561
rect 1430 1527 1468 1561
rect 1502 1527 1540 1561
rect 1574 1527 1612 1561
rect 1646 1527 1684 1561
rect 1718 1527 1756 1561
rect 1790 1527 1828 1561
rect 1862 1527 1900 1561
rect 1934 1527 1972 1561
rect 2006 1527 2044 1561
rect 2078 1527 2116 1561
rect 2150 1527 2188 1561
rect 2222 1527 2260 1561
rect 2294 1527 2332 1561
rect 2366 1527 2404 1561
rect 2438 1527 2476 1561
rect 2510 1527 2548 1561
rect 2582 1527 2620 1561
rect 2654 1527 2692 1561
rect 2726 1527 2764 1561
rect 2798 1527 2836 1561
rect 2870 1527 2908 1561
rect 2942 1527 2980 1561
rect 3014 1527 3052 1561
rect 3086 1527 3124 1561
rect 3158 1527 3196 1561
rect 3230 1527 3268 1561
rect 3302 1527 3340 1561
rect 3374 1527 3412 1561
rect 3446 1527 3484 1561
rect 3518 1527 3556 1561
rect 3590 1527 3628 1561
rect 3662 1527 3700 1561
rect 3734 1527 3772 1561
rect 3806 1527 3844 1561
rect 3878 1527 3916 1561
rect 3950 1527 3988 1561
rect 4022 1527 4060 1561
rect 4094 1527 4132 1561
rect 4166 1527 4204 1561
rect 4238 1527 4276 1561
rect 4310 1527 4348 1561
rect 4382 1527 4420 1561
rect 4454 1527 4492 1561
rect 4526 1527 4564 1561
rect 4598 1527 4636 1561
rect 4670 1527 4708 1561
rect 4742 1527 4780 1561
rect 4814 1527 4852 1561
rect 4886 1527 4924 1561
rect 4958 1527 4996 1561
rect 5030 1527 5068 1561
rect 5102 1527 5140 1561
rect 5174 1527 5212 1561
rect 5246 1527 5284 1561
rect 5318 1527 5356 1561
rect 5390 1527 5428 1561
rect 5462 1527 5500 1561
rect 5534 1527 5572 1561
rect 5606 1527 5644 1561
rect 5678 1527 5716 1561
rect 5750 1527 5788 1561
rect 5822 1527 5860 1561
rect 5894 1527 5932 1561
rect 5966 1527 6004 1561
rect 6038 1527 6076 1561
rect 6110 1527 6148 1561
rect 6182 1527 6220 1561
rect 6254 1527 6292 1561
rect 6326 1527 6364 1561
rect 6398 1527 6436 1561
rect 6470 1527 6508 1561
rect 6542 1527 6580 1561
rect 6614 1527 6652 1561
rect 6686 1527 6724 1561
rect 6758 1527 6796 1561
rect 6830 1527 6868 1561
rect 6902 1527 6940 1561
rect 6974 1527 7012 1561
rect 7046 1527 7084 1561
rect 7118 1527 7156 1561
rect 7190 1527 7228 1561
rect 7262 1527 7300 1561
rect 7334 1527 7372 1561
rect 7406 1527 7444 1561
rect 7478 1527 7516 1561
rect 7550 1527 7588 1561
rect 7622 1527 7660 1561
rect 7694 1527 7732 1561
rect 7766 1527 7804 1561
rect 7838 1527 7876 1561
rect 7910 1527 7948 1561
rect 7982 1527 8020 1561
rect 8054 1527 8120 1561
rect 106 1521 8120 1527
rect 325 1447 7901 1521
rect 106 1377 284 1401
rect 106 1325 176 1377
rect 228 1325 284 1377
rect 106 1301 284 1325
rect 325 1061 7901 1255
rect 106 915 284 1015
rect 106 569 8120 868
rect 106 423 284 523
rect 316 183 3986 377
rect 166 113 284 137
rect 166 61 176 113
rect 228 61 284 113
rect 166 37 284 61
rect 316 -83 3986 -9
rect 106 -89 8120 -83
rect 106 -123 154 -89
rect 188 -123 226 -89
rect 260 -123 298 -89
rect 332 -123 370 -89
rect 404 -123 442 -89
rect 476 -123 514 -89
rect 548 -123 586 -89
rect 620 -123 658 -89
rect 692 -123 730 -89
rect 764 -123 802 -89
rect 836 -123 874 -89
rect 908 -123 946 -89
rect 980 -123 1018 -89
rect 1052 -123 1090 -89
rect 1124 -123 1162 -89
rect 1196 -123 1234 -89
rect 1268 -123 1306 -89
rect 1340 -123 1378 -89
rect 1412 -123 1450 -89
rect 1484 -123 1522 -89
rect 1556 -123 1594 -89
rect 1628 -123 1666 -89
rect 1700 -123 1738 -89
rect 1772 -123 1810 -89
rect 1844 -123 1882 -89
rect 1916 -123 1954 -89
rect 1988 -123 2026 -89
rect 2060 -123 2098 -89
rect 2132 -123 2170 -89
rect 2204 -123 2242 -89
rect 2276 -123 2314 -89
rect 2348 -123 2386 -89
rect 2420 -123 2458 -89
rect 2492 -123 2530 -89
rect 2564 -123 2602 -89
rect 2636 -123 2674 -89
rect 2708 -123 2746 -89
rect 2780 -123 2818 -89
rect 2852 -123 2890 -89
rect 2924 -123 2962 -89
rect 2996 -123 3034 -89
rect 3068 -123 3106 -89
rect 3140 -123 3178 -89
rect 3212 -123 3250 -89
rect 3284 -123 3322 -89
rect 3356 -123 3394 -89
rect 3428 -123 3466 -89
rect 3500 -123 3538 -89
rect 3572 -123 3610 -89
rect 3644 -123 3682 -89
rect 3716 -123 3754 -89
rect 3788 -123 3826 -89
rect 3860 -123 3898 -89
rect 3932 -123 3970 -89
rect 4004 -123 4042 -89
rect 4076 -123 4114 -89
rect 4148 -123 8120 -89
rect 106 -159 8120 -123
<< via1 >>
rect 176 1325 228 1377
rect 176 61 228 113
<< metal2 >>
rect 176 1377 228 1411
rect 176 113 228 1325
rect 176 27 228 61
use sky130_fd_pr__nfet_01v8_DPTN2D  sky130_fd_pr__nfet_01v8_DPTN2D_0
timestamp 1750100919
transform 0 1 2151 -1 0 87
box -236 -2035 236 2035
use sky130_fd_pr__pfet_01v8_D9QHA6  sky130_fd_pr__pfet_01v8_D9QHA6_0
timestamp 1750100919
transform 0 1 4113 -1 0 965
box -246 -4007 246 4007
use sky130_fd_pr__pfet_01v8_D9QHA6  XM1
timestamp 1750100919
transform 0 1 4113 -1 0 1351
box -246 -4007 246 4007
use sky130_fd_pr__nfet_01v8_DPTN2D  XM3
timestamp 1750100919
transform 0 1 2151 -1 0 473
box -236 -2035 236 2035
<< labels >>
flabel metal1 s 117 1553 126 1563 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 118 1345 127 1355 0 FreeSans 500 0 0 0 IN
port 2 nsew
flabel metal1 s 123 958 132 968 0 FreeSans 500 0 0 0 CKB
port 3 nsew
flabel metal1 s 120 467 129 477 0 FreeSans 500 0 0 0 CK
port 4 nsew
flabel metal1 s 121 -124 130 -114 0 FreeSans 500 0 0 0 VSS
port 5 nsew
flabel metal1 s 8079 708 8088 718 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
