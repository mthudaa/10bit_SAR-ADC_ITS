magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect -17 369 -7 403
rect 27 369 65 403
rect 99 369 137 403
rect 171 369 209 403
rect 243 369 281 403
rect 315 369 353 403
rect 387 369 425 403
rect 459 369 497 403
rect 531 369 569 403
rect 603 369 641 403
rect 675 369 713 403
rect 747 369 785 403
rect 819 369 857 403
rect 891 369 929 403
rect 963 369 1001 403
rect 1035 369 1073 403
rect 1107 369 1145 403
rect 1179 369 1217 403
rect 1251 369 1289 403
rect 1323 369 1361 403
rect 1395 369 1433 403
rect 1467 369 1505 403
rect 1539 369 1577 403
rect 1611 369 1649 403
rect 1683 369 1721 403
rect 1755 369 1793 403
rect 1827 369 1865 403
rect 1899 369 1937 403
rect 1971 369 2009 403
rect 2043 369 2081 403
rect 2115 369 2153 403
rect 2187 369 2225 403
rect 2259 369 2297 403
rect 2331 369 2369 403
rect 2403 369 2441 403
rect 2475 369 2513 403
rect 2547 369 2585 403
rect 2619 369 2657 403
rect 2691 369 2729 403
rect 2763 369 2801 403
rect 2835 369 2873 403
rect 2907 369 2945 403
rect 2979 369 3017 403
rect 3051 369 3089 403
rect 3123 369 3161 403
rect 3195 369 3233 403
rect 3267 369 3305 403
rect 3339 369 3377 403
rect 3411 369 3449 403
rect 3483 369 3521 403
rect 3555 369 3593 403
rect 3627 369 3665 403
rect 3699 369 3737 403
rect 3771 369 3809 403
rect 3843 369 3881 403
rect 3915 369 3953 403
rect 3987 369 4025 403
rect 4059 369 4097 403
rect 4131 369 4169 403
rect 4203 369 4241 403
rect 4275 369 4313 403
rect 4347 369 4385 403
rect 4419 369 4457 403
rect 4491 369 4501 403
rect 4607 -17 4645 17
rect 4679 -17 4717 17
rect 4751 -17 4789 17
rect 4823 -17 4861 17
rect 4895 -17 4933 17
rect 4967 -17 5005 17
rect 5039 -17 5077 17
rect 5111 -17 5149 17
rect 5183 -17 5221 17
rect 5255 -17 5293 17
rect 5327 -17 5365 17
rect 5399 -17 5437 17
rect 5471 -17 5509 17
rect 5543 -17 5581 17
rect 5615 -17 5653 17
rect 5687 -17 5725 17
rect 5759 -17 5797 17
rect 5831 -17 5869 17
rect 5903 -17 5941 17
rect 5975 -17 6013 17
rect 6047 -17 6085 17
rect 6119 -17 6157 17
rect 6191 -17 6229 17
rect 6263 -17 6301 17
rect 6335 -17 6373 17
rect 6407 -17 6445 17
rect 6479 -17 6517 17
rect 6551 -17 6589 17
rect 6623 -17 6661 17
rect 6695 -17 6733 17
rect 6767 -17 6805 17
rect 6839 -17 6877 17
<< viali >>
rect -7 369 27 403
rect 65 369 99 403
rect 137 369 171 403
rect 209 369 243 403
rect 281 369 315 403
rect 353 369 387 403
rect 425 369 459 403
rect 497 369 531 403
rect 569 369 603 403
rect 641 369 675 403
rect 713 369 747 403
rect 785 369 819 403
rect 857 369 891 403
rect 929 369 963 403
rect 1001 369 1035 403
rect 1073 369 1107 403
rect 1145 369 1179 403
rect 1217 369 1251 403
rect 1289 369 1323 403
rect 1361 369 1395 403
rect 1433 369 1467 403
rect 1505 369 1539 403
rect 1577 369 1611 403
rect 1649 369 1683 403
rect 1721 369 1755 403
rect 1793 369 1827 403
rect 1865 369 1899 403
rect 1937 369 1971 403
rect 2009 369 2043 403
rect 2081 369 2115 403
rect 2153 369 2187 403
rect 2225 369 2259 403
rect 2297 369 2331 403
rect 2369 369 2403 403
rect 2441 369 2475 403
rect 2513 369 2547 403
rect 2585 369 2619 403
rect 2657 369 2691 403
rect 2729 369 2763 403
rect 2801 369 2835 403
rect 2873 369 2907 403
rect 2945 369 2979 403
rect 3017 369 3051 403
rect 3089 369 3123 403
rect 3161 369 3195 403
rect 3233 369 3267 403
rect 3305 369 3339 403
rect 3377 369 3411 403
rect 3449 369 3483 403
rect 3521 369 3555 403
rect 3593 369 3627 403
rect 3665 369 3699 403
rect 3737 369 3771 403
rect 3809 369 3843 403
rect 3881 369 3915 403
rect 3953 369 3987 403
rect 4025 369 4059 403
rect 4097 369 4131 403
rect 4169 369 4203 403
rect 4241 369 4275 403
rect 4313 369 4347 403
rect 4385 369 4419 403
rect 4457 369 4491 403
rect 4573 -17 4607 17
rect 4645 -17 4679 17
rect 4717 -17 4751 17
rect 4789 -17 4823 17
rect 4861 -17 4895 17
rect 4933 -17 4967 17
rect 5005 -17 5039 17
rect 5077 -17 5111 17
rect 5149 -17 5183 17
rect 5221 -17 5255 17
rect 5293 -17 5327 17
rect 5365 -17 5399 17
rect 5437 -17 5471 17
rect 5509 -17 5543 17
rect 5581 -17 5615 17
rect 5653 -17 5687 17
rect 5725 -17 5759 17
rect 5797 -17 5831 17
rect 5869 -17 5903 17
rect 5941 -17 5975 17
rect 6013 -17 6047 17
rect 6085 -17 6119 17
rect 6157 -17 6191 17
rect 6229 -17 6263 17
rect 6301 -17 6335 17
rect 6373 -17 6407 17
rect 6445 -17 6479 17
rect 6517 -17 6551 17
rect 6589 -17 6623 17
rect 6661 -17 6695 17
rect 6733 -17 6767 17
rect 6805 -17 6839 17
rect 6877 -17 6911 17
<< metal1 >>
rect -53 403 6947 439
rect -53 369 -7 403
rect 27 369 65 403
rect 99 369 137 403
rect 171 369 209 403
rect 243 369 281 403
rect 315 369 353 403
rect 387 369 425 403
rect 459 369 497 403
rect 531 369 569 403
rect 603 369 641 403
rect 675 369 713 403
rect 747 369 785 403
rect 819 369 857 403
rect 891 369 929 403
rect 963 369 1001 403
rect 1035 369 1073 403
rect 1107 369 1145 403
rect 1179 369 1217 403
rect 1251 369 1289 403
rect 1323 369 1361 403
rect 1395 369 1433 403
rect 1467 369 1505 403
rect 1539 369 1577 403
rect 1611 369 1649 403
rect 1683 369 1721 403
rect 1755 369 1793 403
rect 1827 369 1865 403
rect 1899 369 1937 403
rect 1971 369 2009 403
rect 2043 369 2081 403
rect 2115 369 2153 403
rect 2187 369 2225 403
rect 2259 369 2297 403
rect 2331 369 2369 403
rect 2403 369 2441 403
rect 2475 369 2513 403
rect 2547 369 2585 403
rect 2619 369 2657 403
rect 2691 369 2729 403
rect 2763 369 2801 403
rect 2835 369 2873 403
rect 2907 369 2945 403
rect 2979 369 3017 403
rect 3051 369 3089 403
rect 3123 369 3161 403
rect 3195 369 3233 403
rect 3267 369 3305 403
rect 3339 369 3377 403
rect 3411 369 3449 403
rect 3483 369 3521 403
rect 3555 369 3593 403
rect 3627 369 3665 403
rect 3699 369 3737 403
rect 3771 369 3809 403
rect 3843 369 3881 403
rect 3915 369 3953 403
rect 3987 369 4025 403
rect 4059 369 4097 403
rect 4131 369 4169 403
rect 4203 369 4241 403
rect 4275 369 4313 403
rect 4347 369 4385 403
rect 4419 369 4457 403
rect 4491 369 6947 403
rect -53 363 6947 369
rect -53 289 6737 323
rect -53 143 125 243
rect 6769 143 6947 243
rect 166 63 6947 97
rect -53 17 6947 23
rect -53 -17 4573 17
rect 4607 -17 4645 17
rect 4679 -17 4717 17
rect 4751 -17 4789 17
rect 4823 -17 4861 17
rect 4895 -17 4933 17
rect 4967 -17 5005 17
rect 5039 -17 5077 17
rect 5111 -17 5149 17
rect 5183 -17 5221 17
rect 5255 -17 5293 17
rect 5327 -17 5365 17
rect 5399 -17 5437 17
rect 5471 -17 5509 17
rect 5543 -17 5581 17
rect 5615 -17 5653 17
rect 5687 -17 5725 17
rect 5759 -17 5797 17
rect 5831 -17 5869 17
rect 5903 -17 5941 17
rect 5975 -17 6013 17
rect 6047 -17 6085 17
rect 6119 -17 6157 17
rect 6191 -17 6229 17
rect 6263 -17 6301 17
rect 6335 -17 6373 17
rect 6407 -17 6445 17
rect 6479 -17 6517 17
rect 6551 -17 6589 17
rect 6623 -17 6661 17
rect 6695 -17 6733 17
rect 6767 -17 6805 17
rect 6839 -17 6877 17
rect 6911 -17 6947 17
rect -53 -53 6947 -17
use sky130_fd_pr__pfet_01v8_D9QZ56  XM1
timestamp 1750100919
transform 0 1 2242 -1 0 193
box -246 -2295 246 2295
use sky130_fd_pr__nfet_01v8_55NS9E  XM2
timestamp 1750100919
transform 0 1 5742 -1 0 193
box -236 -1195 236 1195
<< labels >>
flabel metal1 s -42 391 -33 401 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s -39 -19 -30 -9 0 FreeSans 500 0 0 0 VSS
port 2 nsew
flabel metal1 s -41 302 -32 312 0 FreeSans 500 0 0 0 IN
port 3 nsew
flabel metal1 s -40 184 -31 194 0 FreeSans 500 0 0 0 SWP
port 4 nsew
flabel metal1 s 6924 187 6933 197 0 FreeSans 500 0 0 0 SWN
port 5 nsew
flabel metal1 s 6927 74 6936 84 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
