magic
tech sky130A
magscale 1 2
timestamp 1748849030
<< metal3 >>
rect -23884 18332 -22712 18360
rect -23884 17508 -22796 18332
rect -22732 17508 -22712 18332
rect -23884 17480 -22712 17508
rect -22472 18332 -21300 18360
rect -22472 17508 -21384 18332
rect -21320 17508 -21300 18332
rect -22472 17480 -21300 17508
rect -21060 18332 -19888 18360
rect -21060 17508 -19972 18332
rect -19908 17508 -19888 18332
rect -21060 17480 -19888 17508
rect -19648 18332 -18476 18360
rect -19648 17508 -18560 18332
rect -18496 17508 -18476 18332
rect -19648 17480 -18476 17508
rect -18236 18332 -17064 18360
rect -18236 17508 -17148 18332
rect -17084 17508 -17064 18332
rect -18236 17480 -17064 17508
rect -16824 18332 -15652 18360
rect -16824 17508 -15736 18332
rect -15672 17508 -15652 18332
rect -16824 17480 -15652 17508
rect -15412 18332 -14240 18360
rect -15412 17508 -14324 18332
rect -14260 17508 -14240 18332
rect -15412 17480 -14240 17508
rect -14000 18332 -12828 18360
rect -14000 17508 -12912 18332
rect -12848 17508 -12828 18332
rect -14000 17480 -12828 17508
rect -12588 18332 -11416 18360
rect -12588 17508 -11500 18332
rect -11436 17508 -11416 18332
rect -12588 17480 -11416 17508
rect -11176 18332 -10004 18360
rect -11176 17508 -10088 18332
rect -10024 17508 -10004 18332
rect -11176 17480 -10004 17508
rect -9764 18332 -8592 18360
rect -9764 17508 -8676 18332
rect -8612 17508 -8592 18332
rect -9764 17480 -8592 17508
rect -8352 18332 -7180 18360
rect -8352 17508 -7264 18332
rect -7200 17508 -7180 18332
rect -8352 17480 -7180 17508
rect -6940 18332 -5768 18360
rect -6940 17508 -5852 18332
rect -5788 17508 -5768 18332
rect -6940 17480 -5768 17508
rect -5528 18332 -4356 18360
rect -5528 17508 -4440 18332
rect -4376 17508 -4356 18332
rect -5528 17480 -4356 17508
rect -4116 18332 -2944 18360
rect -4116 17508 -3028 18332
rect -2964 17508 -2944 18332
rect -4116 17480 -2944 17508
rect -2704 18332 -1532 18360
rect -2704 17508 -1616 18332
rect -1552 17508 -1532 18332
rect -2704 17480 -1532 17508
rect -1292 18332 -120 18360
rect -1292 17508 -204 18332
rect -140 17508 -120 18332
rect -1292 17480 -120 17508
rect 120 18332 1292 18360
rect 120 17508 1208 18332
rect 1272 17508 1292 18332
rect 120 17480 1292 17508
rect 1532 18332 2704 18360
rect 1532 17508 2620 18332
rect 2684 17508 2704 18332
rect 1532 17480 2704 17508
rect 2944 18332 4116 18360
rect 2944 17508 4032 18332
rect 4096 17508 4116 18332
rect 2944 17480 4116 17508
rect 4356 18332 5528 18360
rect 4356 17508 5444 18332
rect 5508 17508 5528 18332
rect 4356 17480 5528 17508
rect 5768 18332 6940 18360
rect 5768 17508 6856 18332
rect 6920 17508 6940 18332
rect 5768 17480 6940 17508
rect 7180 18332 8352 18360
rect 7180 17508 8268 18332
rect 8332 17508 8352 18332
rect 7180 17480 8352 17508
rect 8592 18332 9764 18360
rect 8592 17508 9680 18332
rect 9744 17508 9764 18332
rect 8592 17480 9764 17508
rect 10004 18332 11176 18360
rect 10004 17508 11092 18332
rect 11156 17508 11176 18332
rect 10004 17480 11176 17508
rect 11416 18332 12588 18360
rect 11416 17508 12504 18332
rect 12568 17508 12588 18332
rect 11416 17480 12588 17508
rect 12828 18332 14000 18360
rect 12828 17508 13916 18332
rect 13980 17508 14000 18332
rect 12828 17480 14000 17508
rect 14240 18332 15412 18360
rect 14240 17508 15328 18332
rect 15392 17508 15412 18332
rect 14240 17480 15412 17508
rect 15652 18332 16824 18360
rect 15652 17508 16740 18332
rect 16804 17508 16824 18332
rect 15652 17480 16824 17508
rect 17064 18332 18236 18360
rect 17064 17508 18152 18332
rect 18216 17508 18236 18332
rect 17064 17480 18236 17508
rect 18476 18332 19648 18360
rect 18476 17508 19564 18332
rect 19628 17508 19648 18332
rect 18476 17480 19648 17508
rect 19888 18332 21060 18360
rect 19888 17508 20976 18332
rect 21040 17508 21060 18332
rect 19888 17480 21060 17508
rect 21300 18332 22472 18360
rect 21300 17508 22388 18332
rect 22452 17508 22472 18332
rect 21300 17480 22472 17508
rect 22712 18332 23884 18360
rect 22712 17508 23800 18332
rect 23864 17508 23884 18332
rect 22712 17480 23884 17508
rect -23884 17212 -22712 17240
rect -23884 16388 -22796 17212
rect -22732 16388 -22712 17212
rect -23884 16360 -22712 16388
rect -22472 17212 -21300 17240
rect -22472 16388 -21384 17212
rect -21320 16388 -21300 17212
rect -22472 16360 -21300 16388
rect -21060 17212 -19888 17240
rect -21060 16388 -19972 17212
rect -19908 16388 -19888 17212
rect -21060 16360 -19888 16388
rect -19648 17212 -18476 17240
rect -19648 16388 -18560 17212
rect -18496 16388 -18476 17212
rect -19648 16360 -18476 16388
rect -18236 17212 -17064 17240
rect -18236 16388 -17148 17212
rect -17084 16388 -17064 17212
rect -18236 16360 -17064 16388
rect -16824 17212 -15652 17240
rect -16824 16388 -15736 17212
rect -15672 16388 -15652 17212
rect -16824 16360 -15652 16388
rect -15412 17212 -14240 17240
rect -15412 16388 -14324 17212
rect -14260 16388 -14240 17212
rect -15412 16360 -14240 16388
rect -14000 17212 -12828 17240
rect -14000 16388 -12912 17212
rect -12848 16388 -12828 17212
rect -14000 16360 -12828 16388
rect -12588 17212 -11416 17240
rect -12588 16388 -11500 17212
rect -11436 16388 -11416 17212
rect -12588 16360 -11416 16388
rect -11176 17212 -10004 17240
rect -11176 16388 -10088 17212
rect -10024 16388 -10004 17212
rect -11176 16360 -10004 16388
rect -9764 17212 -8592 17240
rect -9764 16388 -8676 17212
rect -8612 16388 -8592 17212
rect -9764 16360 -8592 16388
rect -8352 17212 -7180 17240
rect -8352 16388 -7264 17212
rect -7200 16388 -7180 17212
rect -8352 16360 -7180 16388
rect -6940 17212 -5768 17240
rect -6940 16388 -5852 17212
rect -5788 16388 -5768 17212
rect -6940 16360 -5768 16388
rect -5528 17212 -4356 17240
rect -5528 16388 -4440 17212
rect -4376 16388 -4356 17212
rect -5528 16360 -4356 16388
rect -4116 17212 -2944 17240
rect -4116 16388 -3028 17212
rect -2964 16388 -2944 17212
rect -4116 16360 -2944 16388
rect -2704 17212 -1532 17240
rect -2704 16388 -1616 17212
rect -1552 16388 -1532 17212
rect -2704 16360 -1532 16388
rect -1292 17212 -120 17240
rect -1292 16388 -204 17212
rect -140 16388 -120 17212
rect -1292 16360 -120 16388
rect 120 17212 1292 17240
rect 120 16388 1208 17212
rect 1272 16388 1292 17212
rect 120 16360 1292 16388
rect 1532 17212 2704 17240
rect 1532 16388 2620 17212
rect 2684 16388 2704 17212
rect 1532 16360 2704 16388
rect 2944 17212 4116 17240
rect 2944 16388 4032 17212
rect 4096 16388 4116 17212
rect 2944 16360 4116 16388
rect 4356 17212 5528 17240
rect 4356 16388 5444 17212
rect 5508 16388 5528 17212
rect 4356 16360 5528 16388
rect 5768 17212 6940 17240
rect 5768 16388 6856 17212
rect 6920 16388 6940 17212
rect 5768 16360 6940 16388
rect 7180 17212 8352 17240
rect 7180 16388 8268 17212
rect 8332 16388 8352 17212
rect 7180 16360 8352 16388
rect 8592 17212 9764 17240
rect 8592 16388 9680 17212
rect 9744 16388 9764 17212
rect 8592 16360 9764 16388
rect 10004 17212 11176 17240
rect 10004 16388 11092 17212
rect 11156 16388 11176 17212
rect 10004 16360 11176 16388
rect 11416 17212 12588 17240
rect 11416 16388 12504 17212
rect 12568 16388 12588 17212
rect 11416 16360 12588 16388
rect 12828 17212 14000 17240
rect 12828 16388 13916 17212
rect 13980 16388 14000 17212
rect 12828 16360 14000 16388
rect 14240 17212 15412 17240
rect 14240 16388 15328 17212
rect 15392 16388 15412 17212
rect 14240 16360 15412 16388
rect 15652 17212 16824 17240
rect 15652 16388 16740 17212
rect 16804 16388 16824 17212
rect 15652 16360 16824 16388
rect 17064 17212 18236 17240
rect 17064 16388 18152 17212
rect 18216 16388 18236 17212
rect 17064 16360 18236 16388
rect 18476 17212 19648 17240
rect 18476 16388 19564 17212
rect 19628 16388 19648 17212
rect 18476 16360 19648 16388
rect 19888 17212 21060 17240
rect 19888 16388 20976 17212
rect 21040 16388 21060 17212
rect 19888 16360 21060 16388
rect 21300 17212 22472 17240
rect 21300 16388 22388 17212
rect 22452 16388 22472 17212
rect 21300 16360 22472 16388
rect 22712 17212 23884 17240
rect 22712 16388 23800 17212
rect 23864 16388 23884 17212
rect 22712 16360 23884 16388
rect -23884 16092 -22712 16120
rect -23884 15268 -22796 16092
rect -22732 15268 -22712 16092
rect -23884 15240 -22712 15268
rect -22472 16092 -21300 16120
rect -22472 15268 -21384 16092
rect -21320 15268 -21300 16092
rect -22472 15240 -21300 15268
rect -21060 16092 -19888 16120
rect -21060 15268 -19972 16092
rect -19908 15268 -19888 16092
rect -21060 15240 -19888 15268
rect -19648 16092 -18476 16120
rect -19648 15268 -18560 16092
rect -18496 15268 -18476 16092
rect -19648 15240 -18476 15268
rect -18236 16092 -17064 16120
rect -18236 15268 -17148 16092
rect -17084 15268 -17064 16092
rect -18236 15240 -17064 15268
rect -16824 16092 -15652 16120
rect -16824 15268 -15736 16092
rect -15672 15268 -15652 16092
rect -16824 15240 -15652 15268
rect -15412 16092 -14240 16120
rect -15412 15268 -14324 16092
rect -14260 15268 -14240 16092
rect -15412 15240 -14240 15268
rect -14000 16092 -12828 16120
rect -14000 15268 -12912 16092
rect -12848 15268 -12828 16092
rect -14000 15240 -12828 15268
rect -12588 16092 -11416 16120
rect -12588 15268 -11500 16092
rect -11436 15268 -11416 16092
rect -12588 15240 -11416 15268
rect -11176 16092 -10004 16120
rect -11176 15268 -10088 16092
rect -10024 15268 -10004 16092
rect -11176 15240 -10004 15268
rect -9764 16092 -8592 16120
rect -9764 15268 -8676 16092
rect -8612 15268 -8592 16092
rect -9764 15240 -8592 15268
rect -8352 16092 -7180 16120
rect -8352 15268 -7264 16092
rect -7200 15268 -7180 16092
rect -8352 15240 -7180 15268
rect -6940 16092 -5768 16120
rect -6940 15268 -5852 16092
rect -5788 15268 -5768 16092
rect -6940 15240 -5768 15268
rect -5528 16092 -4356 16120
rect -5528 15268 -4440 16092
rect -4376 15268 -4356 16092
rect -5528 15240 -4356 15268
rect -4116 16092 -2944 16120
rect -4116 15268 -3028 16092
rect -2964 15268 -2944 16092
rect -4116 15240 -2944 15268
rect -2704 16092 -1532 16120
rect -2704 15268 -1616 16092
rect -1552 15268 -1532 16092
rect -2704 15240 -1532 15268
rect -1292 16092 -120 16120
rect -1292 15268 -204 16092
rect -140 15268 -120 16092
rect -1292 15240 -120 15268
rect 120 16092 1292 16120
rect 120 15268 1208 16092
rect 1272 15268 1292 16092
rect 120 15240 1292 15268
rect 1532 16092 2704 16120
rect 1532 15268 2620 16092
rect 2684 15268 2704 16092
rect 1532 15240 2704 15268
rect 2944 16092 4116 16120
rect 2944 15268 4032 16092
rect 4096 15268 4116 16092
rect 2944 15240 4116 15268
rect 4356 16092 5528 16120
rect 4356 15268 5444 16092
rect 5508 15268 5528 16092
rect 4356 15240 5528 15268
rect 5768 16092 6940 16120
rect 5768 15268 6856 16092
rect 6920 15268 6940 16092
rect 5768 15240 6940 15268
rect 7180 16092 8352 16120
rect 7180 15268 8268 16092
rect 8332 15268 8352 16092
rect 7180 15240 8352 15268
rect 8592 16092 9764 16120
rect 8592 15268 9680 16092
rect 9744 15268 9764 16092
rect 8592 15240 9764 15268
rect 10004 16092 11176 16120
rect 10004 15268 11092 16092
rect 11156 15268 11176 16092
rect 10004 15240 11176 15268
rect 11416 16092 12588 16120
rect 11416 15268 12504 16092
rect 12568 15268 12588 16092
rect 11416 15240 12588 15268
rect 12828 16092 14000 16120
rect 12828 15268 13916 16092
rect 13980 15268 14000 16092
rect 12828 15240 14000 15268
rect 14240 16092 15412 16120
rect 14240 15268 15328 16092
rect 15392 15268 15412 16092
rect 14240 15240 15412 15268
rect 15652 16092 16824 16120
rect 15652 15268 16740 16092
rect 16804 15268 16824 16092
rect 15652 15240 16824 15268
rect 17064 16092 18236 16120
rect 17064 15268 18152 16092
rect 18216 15268 18236 16092
rect 17064 15240 18236 15268
rect 18476 16092 19648 16120
rect 18476 15268 19564 16092
rect 19628 15268 19648 16092
rect 18476 15240 19648 15268
rect 19888 16092 21060 16120
rect 19888 15268 20976 16092
rect 21040 15268 21060 16092
rect 19888 15240 21060 15268
rect 21300 16092 22472 16120
rect 21300 15268 22388 16092
rect 22452 15268 22472 16092
rect 21300 15240 22472 15268
rect 22712 16092 23884 16120
rect 22712 15268 23800 16092
rect 23864 15268 23884 16092
rect 22712 15240 23884 15268
rect -23884 14972 -22712 15000
rect -23884 14148 -22796 14972
rect -22732 14148 -22712 14972
rect -23884 14120 -22712 14148
rect -22472 14972 -21300 15000
rect -22472 14148 -21384 14972
rect -21320 14148 -21300 14972
rect -22472 14120 -21300 14148
rect -21060 14972 -19888 15000
rect -21060 14148 -19972 14972
rect -19908 14148 -19888 14972
rect -21060 14120 -19888 14148
rect -19648 14972 -18476 15000
rect -19648 14148 -18560 14972
rect -18496 14148 -18476 14972
rect -19648 14120 -18476 14148
rect -18236 14972 -17064 15000
rect -18236 14148 -17148 14972
rect -17084 14148 -17064 14972
rect -18236 14120 -17064 14148
rect -16824 14972 -15652 15000
rect -16824 14148 -15736 14972
rect -15672 14148 -15652 14972
rect -16824 14120 -15652 14148
rect -15412 14972 -14240 15000
rect -15412 14148 -14324 14972
rect -14260 14148 -14240 14972
rect -15412 14120 -14240 14148
rect -14000 14972 -12828 15000
rect -14000 14148 -12912 14972
rect -12848 14148 -12828 14972
rect -14000 14120 -12828 14148
rect -12588 14972 -11416 15000
rect -12588 14148 -11500 14972
rect -11436 14148 -11416 14972
rect -12588 14120 -11416 14148
rect -11176 14972 -10004 15000
rect -11176 14148 -10088 14972
rect -10024 14148 -10004 14972
rect -11176 14120 -10004 14148
rect -9764 14972 -8592 15000
rect -9764 14148 -8676 14972
rect -8612 14148 -8592 14972
rect -9764 14120 -8592 14148
rect -8352 14972 -7180 15000
rect -8352 14148 -7264 14972
rect -7200 14148 -7180 14972
rect -8352 14120 -7180 14148
rect -6940 14972 -5768 15000
rect -6940 14148 -5852 14972
rect -5788 14148 -5768 14972
rect -6940 14120 -5768 14148
rect -5528 14972 -4356 15000
rect -5528 14148 -4440 14972
rect -4376 14148 -4356 14972
rect -5528 14120 -4356 14148
rect -4116 14972 -2944 15000
rect -4116 14148 -3028 14972
rect -2964 14148 -2944 14972
rect -4116 14120 -2944 14148
rect -2704 14972 -1532 15000
rect -2704 14148 -1616 14972
rect -1552 14148 -1532 14972
rect -2704 14120 -1532 14148
rect -1292 14972 -120 15000
rect -1292 14148 -204 14972
rect -140 14148 -120 14972
rect -1292 14120 -120 14148
rect 120 14972 1292 15000
rect 120 14148 1208 14972
rect 1272 14148 1292 14972
rect 120 14120 1292 14148
rect 1532 14972 2704 15000
rect 1532 14148 2620 14972
rect 2684 14148 2704 14972
rect 1532 14120 2704 14148
rect 2944 14972 4116 15000
rect 2944 14148 4032 14972
rect 4096 14148 4116 14972
rect 2944 14120 4116 14148
rect 4356 14972 5528 15000
rect 4356 14148 5444 14972
rect 5508 14148 5528 14972
rect 4356 14120 5528 14148
rect 5768 14972 6940 15000
rect 5768 14148 6856 14972
rect 6920 14148 6940 14972
rect 5768 14120 6940 14148
rect 7180 14972 8352 15000
rect 7180 14148 8268 14972
rect 8332 14148 8352 14972
rect 7180 14120 8352 14148
rect 8592 14972 9764 15000
rect 8592 14148 9680 14972
rect 9744 14148 9764 14972
rect 8592 14120 9764 14148
rect 10004 14972 11176 15000
rect 10004 14148 11092 14972
rect 11156 14148 11176 14972
rect 10004 14120 11176 14148
rect 11416 14972 12588 15000
rect 11416 14148 12504 14972
rect 12568 14148 12588 14972
rect 11416 14120 12588 14148
rect 12828 14972 14000 15000
rect 12828 14148 13916 14972
rect 13980 14148 14000 14972
rect 12828 14120 14000 14148
rect 14240 14972 15412 15000
rect 14240 14148 15328 14972
rect 15392 14148 15412 14972
rect 14240 14120 15412 14148
rect 15652 14972 16824 15000
rect 15652 14148 16740 14972
rect 16804 14148 16824 14972
rect 15652 14120 16824 14148
rect 17064 14972 18236 15000
rect 17064 14148 18152 14972
rect 18216 14148 18236 14972
rect 17064 14120 18236 14148
rect 18476 14972 19648 15000
rect 18476 14148 19564 14972
rect 19628 14148 19648 14972
rect 18476 14120 19648 14148
rect 19888 14972 21060 15000
rect 19888 14148 20976 14972
rect 21040 14148 21060 14972
rect 19888 14120 21060 14148
rect 21300 14972 22472 15000
rect 21300 14148 22388 14972
rect 22452 14148 22472 14972
rect 21300 14120 22472 14148
rect 22712 14972 23884 15000
rect 22712 14148 23800 14972
rect 23864 14148 23884 14972
rect 22712 14120 23884 14148
rect -23884 13852 -22712 13880
rect -23884 13028 -22796 13852
rect -22732 13028 -22712 13852
rect -23884 13000 -22712 13028
rect -22472 13852 -21300 13880
rect -22472 13028 -21384 13852
rect -21320 13028 -21300 13852
rect -22472 13000 -21300 13028
rect -21060 13852 -19888 13880
rect -21060 13028 -19972 13852
rect -19908 13028 -19888 13852
rect -21060 13000 -19888 13028
rect -19648 13852 -18476 13880
rect -19648 13028 -18560 13852
rect -18496 13028 -18476 13852
rect -19648 13000 -18476 13028
rect -18236 13852 -17064 13880
rect -18236 13028 -17148 13852
rect -17084 13028 -17064 13852
rect -18236 13000 -17064 13028
rect -16824 13852 -15652 13880
rect -16824 13028 -15736 13852
rect -15672 13028 -15652 13852
rect -16824 13000 -15652 13028
rect -15412 13852 -14240 13880
rect -15412 13028 -14324 13852
rect -14260 13028 -14240 13852
rect -15412 13000 -14240 13028
rect -14000 13852 -12828 13880
rect -14000 13028 -12912 13852
rect -12848 13028 -12828 13852
rect -14000 13000 -12828 13028
rect -12588 13852 -11416 13880
rect -12588 13028 -11500 13852
rect -11436 13028 -11416 13852
rect -12588 13000 -11416 13028
rect -11176 13852 -10004 13880
rect -11176 13028 -10088 13852
rect -10024 13028 -10004 13852
rect -11176 13000 -10004 13028
rect -9764 13852 -8592 13880
rect -9764 13028 -8676 13852
rect -8612 13028 -8592 13852
rect -9764 13000 -8592 13028
rect -8352 13852 -7180 13880
rect -8352 13028 -7264 13852
rect -7200 13028 -7180 13852
rect -8352 13000 -7180 13028
rect -6940 13852 -5768 13880
rect -6940 13028 -5852 13852
rect -5788 13028 -5768 13852
rect -6940 13000 -5768 13028
rect -5528 13852 -4356 13880
rect -5528 13028 -4440 13852
rect -4376 13028 -4356 13852
rect -5528 13000 -4356 13028
rect -4116 13852 -2944 13880
rect -4116 13028 -3028 13852
rect -2964 13028 -2944 13852
rect -4116 13000 -2944 13028
rect -2704 13852 -1532 13880
rect -2704 13028 -1616 13852
rect -1552 13028 -1532 13852
rect -2704 13000 -1532 13028
rect -1292 13852 -120 13880
rect -1292 13028 -204 13852
rect -140 13028 -120 13852
rect -1292 13000 -120 13028
rect 120 13852 1292 13880
rect 120 13028 1208 13852
rect 1272 13028 1292 13852
rect 120 13000 1292 13028
rect 1532 13852 2704 13880
rect 1532 13028 2620 13852
rect 2684 13028 2704 13852
rect 1532 13000 2704 13028
rect 2944 13852 4116 13880
rect 2944 13028 4032 13852
rect 4096 13028 4116 13852
rect 2944 13000 4116 13028
rect 4356 13852 5528 13880
rect 4356 13028 5444 13852
rect 5508 13028 5528 13852
rect 4356 13000 5528 13028
rect 5768 13852 6940 13880
rect 5768 13028 6856 13852
rect 6920 13028 6940 13852
rect 5768 13000 6940 13028
rect 7180 13852 8352 13880
rect 7180 13028 8268 13852
rect 8332 13028 8352 13852
rect 7180 13000 8352 13028
rect 8592 13852 9764 13880
rect 8592 13028 9680 13852
rect 9744 13028 9764 13852
rect 8592 13000 9764 13028
rect 10004 13852 11176 13880
rect 10004 13028 11092 13852
rect 11156 13028 11176 13852
rect 10004 13000 11176 13028
rect 11416 13852 12588 13880
rect 11416 13028 12504 13852
rect 12568 13028 12588 13852
rect 11416 13000 12588 13028
rect 12828 13852 14000 13880
rect 12828 13028 13916 13852
rect 13980 13028 14000 13852
rect 12828 13000 14000 13028
rect 14240 13852 15412 13880
rect 14240 13028 15328 13852
rect 15392 13028 15412 13852
rect 14240 13000 15412 13028
rect 15652 13852 16824 13880
rect 15652 13028 16740 13852
rect 16804 13028 16824 13852
rect 15652 13000 16824 13028
rect 17064 13852 18236 13880
rect 17064 13028 18152 13852
rect 18216 13028 18236 13852
rect 17064 13000 18236 13028
rect 18476 13852 19648 13880
rect 18476 13028 19564 13852
rect 19628 13028 19648 13852
rect 18476 13000 19648 13028
rect 19888 13852 21060 13880
rect 19888 13028 20976 13852
rect 21040 13028 21060 13852
rect 19888 13000 21060 13028
rect 21300 13852 22472 13880
rect 21300 13028 22388 13852
rect 22452 13028 22472 13852
rect 21300 13000 22472 13028
rect 22712 13852 23884 13880
rect 22712 13028 23800 13852
rect 23864 13028 23884 13852
rect 22712 13000 23884 13028
rect -23884 12732 -22712 12760
rect -23884 11908 -22796 12732
rect -22732 11908 -22712 12732
rect -23884 11880 -22712 11908
rect -22472 12732 -21300 12760
rect -22472 11908 -21384 12732
rect -21320 11908 -21300 12732
rect -22472 11880 -21300 11908
rect -21060 12732 -19888 12760
rect -21060 11908 -19972 12732
rect -19908 11908 -19888 12732
rect -21060 11880 -19888 11908
rect -19648 12732 -18476 12760
rect -19648 11908 -18560 12732
rect -18496 11908 -18476 12732
rect -19648 11880 -18476 11908
rect -18236 12732 -17064 12760
rect -18236 11908 -17148 12732
rect -17084 11908 -17064 12732
rect -18236 11880 -17064 11908
rect -16824 12732 -15652 12760
rect -16824 11908 -15736 12732
rect -15672 11908 -15652 12732
rect -16824 11880 -15652 11908
rect -15412 12732 -14240 12760
rect -15412 11908 -14324 12732
rect -14260 11908 -14240 12732
rect -15412 11880 -14240 11908
rect -14000 12732 -12828 12760
rect -14000 11908 -12912 12732
rect -12848 11908 -12828 12732
rect -14000 11880 -12828 11908
rect -12588 12732 -11416 12760
rect -12588 11908 -11500 12732
rect -11436 11908 -11416 12732
rect -12588 11880 -11416 11908
rect -11176 12732 -10004 12760
rect -11176 11908 -10088 12732
rect -10024 11908 -10004 12732
rect -11176 11880 -10004 11908
rect -9764 12732 -8592 12760
rect -9764 11908 -8676 12732
rect -8612 11908 -8592 12732
rect -9764 11880 -8592 11908
rect -8352 12732 -7180 12760
rect -8352 11908 -7264 12732
rect -7200 11908 -7180 12732
rect -8352 11880 -7180 11908
rect -6940 12732 -5768 12760
rect -6940 11908 -5852 12732
rect -5788 11908 -5768 12732
rect -6940 11880 -5768 11908
rect -5528 12732 -4356 12760
rect -5528 11908 -4440 12732
rect -4376 11908 -4356 12732
rect -5528 11880 -4356 11908
rect -4116 12732 -2944 12760
rect -4116 11908 -3028 12732
rect -2964 11908 -2944 12732
rect -4116 11880 -2944 11908
rect -2704 12732 -1532 12760
rect -2704 11908 -1616 12732
rect -1552 11908 -1532 12732
rect -2704 11880 -1532 11908
rect -1292 12732 -120 12760
rect -1292 11908 -204 12732
rect -140 11908 -120 12732
rect -1292 11880 -120 11908
rect 120 12732 1292 12760
rect 120 11908 1208 12732
rect 1272 11908 1292 12732
rect 120 11880 1292 11908
rect 1532 12732 2704 12760
rect 1532 11908 2620 12732
rect 2684 11908 2704 12732
rect 1532 11880 2704 11908
rect 2944 12732 4116 12760
rect 2944 11908 4032 12732
rect 4096 11908 4116 12732
rect 2944 11880 4116 11908
rect 4356 12732 5528 12760
rect 4356 11908 5444 12732
rect 5508 11908 5528 12732
rect 4356 11880 5528 11908
rect 5768 12732 6940 12760
rect 5768 11908 6856 12732
rect 6920 11908 6940 12732
rect 5768 11880 6940 11908
rect 7180 12732 8352 12760
rect 7180 11908 8268 12732
rect 8332 11908 8352 12732
rect 7180 11880 8352 11908
rect 8592 12732 9764 12760
rect 8592 11908 9680 12732
rect 9744 11908 9764 12732
rect 8592 11880 9764 11908
rect 10004 12732 11176 12760
rect 10004 11908 11092 12732
rect 11156 11908 11176 12732
rect 10004 11880 11176 11908
rect 11416 12732 12588 12760
rect 11416 11908 12504 12732
rect 12568 11908 12588 12732
rect 11416 11880 12588 11908
rect 12828 12732 14000 12760
rect 12828 11908 13916 12732
rect 13980 11908 14000 12732
rect 12828 11880 14000 11908
rect 14240 12732 15412 12760
rect 14240 11908 15328 12732
rect 15392 11908 15412 12732
rect 14240 11880 15412 11908
rect 15652 12732 16824 12760
rect 15652 11908 16740 12732
rect 16804 11908 16824 12732
rect 15652 11880 16824 11908
rect 17064 12732 18236 12760
rect 17064 11908 18152 12732
rect 18216 11908 18236 12732
rect 17064 11880 18236 11908
rect 18476 12732 19648 12760
rect 18476 11908 19564 12732
rect 19628 11908 19648 12732
rect 18476 11880 19648 11908
rect 19888 12732 21060 12760
rect 19888 11908 20976 12732
rect 21040 11908 21060 12732
rect 19888 11880 21060 11908
rect 21300 12732 22472 12760
rect 21300 11908 22388 12732
rect 22452 11908 22472 12732
rect 21300 11880 22472 11908
rect 22712 12732 23884 12760
rect 22712 11908 23800 12732
rect 23864 11908 23884 12732
rect 22712 11880 23884 11908
rect -23884 11612 -22712 11640
rect -23884 10788 -22796 11612
rect -22732 10788 -22712 11612
rect -23884 10760 -22712 10788
rect -22472 11612 -21300 11640
rect -22472 10788 -21384 11612
rect -21320 10788 -21300 11612
rect -22472 10760 -21300 10788
rect -21060 11612 -19888 11640
rect -21060 10788 -19972 11612
rect -19908 10788 -19888 11612
rect -21060 10760 -19888 10788
rect -19648 11612 -18476 11640
rect -19648 10788 -18560 11612
rect -18496 10788 -18476 11612
rect -19648 10760 -18476 10788
rect -18236 11612 -17064 11640
rect -18236 10788 -17148 11612
rect -17084 10788 -17064 11612
rect -18236 10760 -17064 10788
rect -16824 11612 -15652 11640
rect -16824 10788 -15736 11612
rect -15672 10788 -15652 11612
rect -16824 10760 -15652 10788
rect -15412 11612 -14240 11640
rect -15412 10788 -14324 11612
rect -14260 10788 -14240 11612
rect -15412 10760 -14240 10788
rect -14000 11612 -12828 11640
rect -14000 10788 -12912 11612
rect -12848 10788 -12828 11612
rect -14000 10760 -12828 10788
rect -12588 11612 -11416 11640
rect -12588 10788 -11500 11612
rect -11436 10788 -11416 11612
rect -12588 10760 -11416 10788
rect -11176 11612 -10004 11640
rect -11176 10788 -10088 11612
rect -10024 10788 -10004 11612
rect -11176 10760 -10004 10788
rect -9764 11612 -8592 11640
rect -9764 10788 -8676 11612
rect -8612 10788 -8592 11612
rect -9764 10760 -8592 10788
rect -8352 11612 -7180 11640
rect -8352 10788 -7264 11612
rect -7200 10788 -7180 11612
rect -8352 10760 -7180 10788
rect -6940 11612 -5768 11640
rect -6940 10788 -5852 11612
rect -5788 10788 -5768 11612
rect -6940 10760 -5768 10788
rect -5528 11612 -4356 11640
rect -5528 10788 -4440 11612
rect -4376 10788 -4356 11612
rect -5528 10760 -4356 10788
rect -4116 11612 -2944 11640
rect -4116 10788 -3028 11612
rect -2964 10788 -2944 11612
rect -4116 10760 -2944 10788
rect -2704 11612 -1532 11640
rect -2704 10788 -1616 11612
rect -1552 10788 -1532 11612
rect -2704 10760 -1532 10788
rect -1292 11612 -120 11640
rect -1292 10788 -204 11612
rect -140 10788 -120 11612
rect -1292 10760 -120 10788
rect 120 11612 1292 11640
rect 120 10788 1208 11612
rect 1272 10788 1292 11612
rect 120 10760 1292 10788
rect 1532 11612 2704 11640
rect 1532 10788 2620 11612
rect 2684 10788 2704 11612
rect 1532 10760 2704 10788
rect 2944 11612 4116 11640
rect 2944 10788 4032 11612
rect 4096 10788 4116 11612
rect 2944 10760 4116 10788
rect 4356 11612 5528 11640
rect 4356 10788 5444 11612
rect 5508 10788 5528 11612
rect 4356 10760 5528 10788
rect 5768 11612 6940 11640
rect 5768 10788 6856 11612
rect 6920 10788 6940 11612
rect 5768 10760 6940 10788
rect 7180 11612 8352 11640
rect 7180 10788 8268 11612
rect 8332 10788 8352 11612
rect 7180 10760 8352 10788
rect 8592 11612 9764 11640
rect 8592 10788 9680 11612
rect 9744 10788 9764 11612
rect 8592 10760 9764 10788
rect 10004 11612 11176 11640
rect 10004 10788 11092 11612
rect 11156 10788 11176 11612
rect 10004 10760 11176 10788
rect 11416 11612 12588 11640
rect 11416 10788 12504 11612
rect 12568 10788 12588 11612
rect 11416 10760 12588 10788
rect 12828 11612 14000 11640
rect 12828 10788 13916 11612
rect 13980 10788 14000 11612
rect 12828 10760 14000 10788
rect 14240 11612 15412 11640
rect 14240 10788 15328 11612
rect 15392 10788 15412 11612
rect 14240 10760 15412 10788
rect 15652 11612 16824 11640
rect 15652 10788 16740 11612
rect 16804 10788 16824 11612
rect 15652 10760 16824 10788
rect 17064 11612 18236 11640
rect 17064 10788 18152 11612
rect 18216 10788 18236 11612
rect 17064 10760 18236 10788
rect 18476 11612 19648 11640
rect 18476 10788 19564 11612
rect 19628 10788 19648 11612
rect 18476 10760 19648 10788
rect 19888 11612 21060 11640
rect 19888 10788 20976 11612
rect 21040 10788 21060 11612
rect 19888 10760 21060 10788
rect 21300 11612 22472 11640
rect 21300 10788 22388 11612
rect 22452 10788 22472 11612
rect 21300 10760 22472 10788
rect 22712 11612 23884 11640
rect 22712 10788 23800 11612
rect 23864 10788 23884 11612
rect 22712 10760 23884 10788
rect -23884 10492 -22712 10520
rect -23884 9668 -22796 10492
rect -22732 9668 -22712 10492
rect -23884 9640 -22712 9668
rect -22472 10492 -21300 10520
rect -22472 9668 -21384 10492
rect -21320 9668 -21300 10492
rect -22472 9640 -21300 9668
rect -21060 10492 -19888 10520
rect -21060 9668 -19972 10492
rect -19908 9668 -19888 10492
rect -21060 9640 -19888 9668
rect -19648 10492 -18476 10520
rect -19648 9668 -18560 10492
rect -18496 9668 -18476 10492
rect -19648 9640 -18476 9668
rect -18236 10492 -17064 10520
rect -18236 9668 -17148 10492
rect -17084 9668 -17064 10492
rect -18236 9640 -17064 9668
rect -16824 10492 -15652 10520
rect -16824 9668 -15736 10492
rect -15672 9668 -15652 10492
rect -16824 9640 -15652 9668
rect -15412 10492 -14240 10520
rect -15412 9668 -14324 10492
rect -14260 9668 -14240 10492
rect -15412 9640 -14240 9668
rect -14000 10492 -12828 10520
rect -14000 9668 -12912 10492
rect -12848 9668 -12828 10492
rect -14000 9640 -12828 9668
rect -12588 10492 -11416 10520
rect -12588 9668 -11500 10492
rect -11436 9668 -11416 10492
rect -12588 9640 -11416 9668
rect -11176 10492 -10004 10520
rect -11176 9668 -10088 10492
rect -10024 9668 -10004 10492
rect -11176 9640 -10004 9668
rect -9764 10492 -8592 10520
rect -9764 9668 -8676 10492
rect -8612 9668 -8592 10492
rect -9764 9640 -8592 9668
rect -8352 10492 -7180 10520
rect -8352 9668 -7264 10492
rect -7200 9668 -7180 10492
rect -8352 9640 -7180 9668
rect -6940 10492 -5768 10520
rect -6940 9668 -5852 10492
rect -5788 9668 -5768 10492
rect -6940 9640 -5768 9668
rect -5528 10492 -4356 10520
rect -5528 9668 -4440 10492
rect -4376 9668 -4356 10492
rect -5528 9640 -4356 9668
rect -4116 10492 -2944 10520
rect -4116 9668 -3028 10492
rect -2964 9668 -2944 10492
rect -4116 9640 -2944 9668
rect -2704 10492 -1532 10520
rect -2704 9668 -1616 10492
rect -1552 9668 -1532 10492
rect -2704 9640 -1532 9668
rect -1292 10492 -120 10520
rect -1292 9668 -204 10492
rect -140 9668 -120 10492
rect -1292 9640 -120 9668
rect 120 10492 1292 10520
rect 120 9668 1208 10492
rect 1272 9668 1292 10492
rect 120 9640 1292 9668
rect 1532 10492 2704 10520
rect 1532 9668 2620 10492
rect 2684 9668 2704 10492
rect 1532 9640 2704 9668
rect 2944 10492 4116 10520
rect 2944 9668 4032 10492
rect 4096 9668 4116 10492
rect 2944 9640 4116 9668
rect 4356 10492 5528 10520
rect 4356 9668 5444 10492
rect 5508 9668 5528 10492
rect 4356 9640 5528 9668
rect 5768 10492 6940 10520
rect 5768 9668 6856 10492
rect 6920 9668 6940 10492
rect 5768 9640 6940 9668
rect 7180 10492 8352 10520
rect 7180 9668 8268 10492
rect 8332 9668 8352 10492
rect 7180 9640 8352 9668
rect 8592 10492 9764 10520
rect 8592 9668 9680 10492
rect 9744 9668 9764 10492
rect 8592 9640 9764 9668
rect 10004 10492 11176 10520
rect 10004 9668 11092 10492
rect 11156 9668 11176 10492
rect 10004 9640 11176 9668
rect 11416 10492 12588 10520
rect 11416 9668 12504 10492
rect 12568 9668 12588 10492
rect 11416 9640 12588 9668
rect 12828 10492 14000 10520
rect 12828 9668 13916 10492
rect 13980 9668 14000 10492
rect 12828 9640 14000 9668
rect 14240 10492 15412 10520
rect 14240 9668 15328 10492
rect 15392 9668 15412 10492
rect 14240 9640 15412 9668
rect 15652 10492 16824 10520
rect 15652 9668 16740 10492
rect 16804 9668 16824 10492
rect 15652 9640 16824 9668
rect 17064 10492 18236 10520
rect 17064 9668 18152 10492
rect 18216 9668 18236 10492
rect 17064 9640 18236 9668
rect 18476 10492 19648 10520
rect 18476 9668 19564 10492
rect 19628 9668 19648 10492
rect 18476 9640 19648 9668
rect 19888 10492 21060 10520
rect 19888 9668 20976 10492
rect 21040 9668 21060 10492
rect 19888 9640 21060 9668
rect 21300 10492 22472 10520
rect 21300 9668 22388 10492
rect 22452 9668 22472 10492
rect 21300 9640 22472 9668
rect 22712 10492 23884 10520
rect 22712 9668 23800 10492
rect 23864 9668 23884 10492
rect 22712 9640 23884 9668
rect -23884 9372 -22712 9400
rect -23884 8548 -22796 9372
rect -22732 8548 -22712 9372
rect -23884 8520 -22712 8548
rect -22472 9372 -21300 9400
rect -22472 8548 -21384 9372
rect -21320 8548 -21300 9372
rect -22472 8520 -21300 8548
rect -21060 9372 -19888 9400
rect -21060 8548 -19972 9372
rect -19908 8548 -19888 9372
rect -21060 8520 -19888 8548
rect -19648 9372 -18476 9400
rect -19648 8548 -18560 9372
rect -18496 8548 -18476 9372
rect -19648 8520 -18476 8548
rect -18236 9372 -17064 9400
rect -18236 8548 -17148 9372
rect -17084 8548 -17064 9372
rect -18236 8520 -17064 8548
rect -16824 9372 -15652 9400
rect -16824 8548 -15736 9372
rect -15672 8548 -15652 9372
rect -16824 8520 -15652 8548
rect -15412 9372 -14240 9400
rect -15412 8548 -14324 9372
rect -14260 8548 -14240 9372
rect -15412 8520 -14240 8548
rect -14000 9372 -12828 9400
rect -14000 8548 -12912 9372
rect -12848 8548 -12828 9372
rect -14000 8520 -12828 8548
rect -12588 9372 -11416 9400
rect -12588 8548 -11500 9372
rect -11436 8548 -11416 9372
rect -12588 8520 -11416 8548
rect -11176 9372 -10004 9400
rect -11176 8548 -10088 9372
rect -10024 8548 -10004 9372
rect -11176 8520 -10004 8548
rect -9764 9372 -8592 9400
rect -9764 8548 -8676 9372
rect -8612 8548 -8592 9372
rect -9764 8520 -8592 8548
rect -8352 9372 -7180 9400
rect -8352 8548 -7264 9372
rect -7200 8548 -7180 9372
rect -8352 8520 -7180 8548
rect -6940 9372 -5768 9400
rect -6940 8548 -5852 9372
rect -5788 8548 -5768 9372
rect -6940 8520 -5768 8548
rect -5528 9372 -4356 9400
rect -5528 8548 -4440 9372
rect -4376 8548 -4356 9372
rect -5528 8520 -4356 8548
rect -4116 9372 -2944 9400
rect -4116 8548 -3028 9372
rect -2964 8548 -2944 9372
rect -4116 8520 -2944 8548
rect -2704 9372 -1532 9400
rect -2704 8548 -1616 9372
rect -1552 8548 -1532 9372
rect -2704 8520 -1532 8548
rect -1292 9372 -120 9400
rect -1292 8548 -204 9372
rect -140 8548 -120 9372
rect -1292 8520 -120 8548
rect 120 9372 1292 9400
rect 120 8548 1208 9372
rect 1272 8548 1292 9372
rect 120 8520 1292 8548
rect 1532 9372 2704 9400
rect 1532 8548 2620 9372
rect 2684 8548 2704 9372
rect 1532 8520 2704 8548
rect 2944 9372 4116 9400
rect 2944 8548 4032 9372
rect 4096 8548 4116 9372
rect 2944 8520 4116 8548
rect 4356 9372 5528 9400
rect 4356 8548 5444 9372
rect 5508 8548 5528 9372
rect 4356 8520 5528 8548
rect 5768 9372 6940 9400
rect 5768 8548 6856 9372
rect 6920 8548 6940 9372
rect 5768 8520 6940 8548
rect 7180 9372 8352 9400
rect 7180 8548 8268 9372
rect 8332 8548 8352 9372
rect 7180 8520 8352 8548
rect 8592 9372 9764 9400
rect 8592 8548 9680 9372
rect 9744 8548 9764 9372
rect 8592 8520 9764 8548
rect 10004 9372 11176 9400
rect 10004 8548 11092 9372
rect 11156 8548 11176 9372
rect 10004 8520 11176 8548
rect 11416 9372 12588 9400
rect 11416 8548 12504 9372
rect 12568 8548 12588 9372
rect 11416 8520 12588 8548
rect 12828 9372 14000 9400
rect 12828 8548 13916 9372
rect 13980 8548 14000 9372
rect 12828 8520 14000 8548
rect 14240 9372 15412 9400
rect 14240 8548 15328 9372
rect 15392 8548 15412 9372
rect 14240 8520 15412 8548
rect 15652 9372 16824 9400
rect 15652 8548 16740 9372
rect 16804 8548 16824 9372
rect 15652 8520 16824 8548
rect 17064 9372 18236 9400
rect 17064 8548 18152 9372
rect 18216 8548 18236 9372
rect 17064 8520 18236 8548
rect 18476 9372 19648 9400
rect 18476 8548 19564 9372
rect 19628 8548 19648 9372
rect 18476 8520 19648 8548
rect 19888 9372 21060 9400
rect 19888 8548 20976 9372
rect 21040 8548 21060 9372
rect 19888 8520 21060 8548
rect 21300 9372 22472 9400
rect 21300 8548 22388 9372
rect 22452 8548 22472 9372
rect 21300 8520 22472 8548
rect 22712 9372 23884 9400
rect 22712 8548 23800 9372
rect 23864 8548 23884 9372
rect 22712 8520 23884 8548
rect -23884 8252 -22712 8280
rect -23884 7428 -22796 8252
rect -22732 7428 -22712 8252
rect -23884 7400 -22712 7428
rect -22472 8252 -21300 8280
rect -22472 7428 -21384 8252
rect -21320 7428 -21300 8252
rect -22472 7400 -21300 7428
rect -21060 8252 -19888 8280
rect -21060 7428 -19972 8252
rect -19908 7428 -19888 8252
rect -21060 7400 -19888 7428
rect -19648 8252 -18476 8280
rect -19648 7428 -18560 8252
rect -18496 7428 -18476 8252
rect -19648 7400 -18476 7428
rect -18236 8252 -17064 8280
rect -18236 7428 -17148 8252
rect -17084 7428 -17064 8252
rect -18236 7400 -17064 7428
rect -16824 8252 -15652 8280
rect -16824 7428 -15736 8252
rect -15672 7428 -15652 8252
rect -16824 7400 -15652 7428
rect -15412 8252 -14240 8280
rect -15412 7428 -14324 8252
rect -14260 7428 -14240 8252
rect -15412 7400 -14240 7428
rect -14000 8252 -12828 8280
rect -14000 7428 -12912 8252
rect -12848 7428 -12828 8252
rect -14000 7400 -12828 7428
rect -12588 8252 -11416 8280
rect -12588 7428 -11500 8252
rect -11436 7428 -11416 8252
rect -12588 7400 -11416 7428
rect -11176 8252 -10004 8280
rect -11176 7428 -10088 8252
rect -10024 7428 -10004 8252
rect -11176 7400 -10004 7428
rect -9764 8252 -8592 8280
rect -9764 7428 -8676 8252
rect -8612 7428 -8592 8252
rect -9764 7400 -8592 7428
rect -8352 8252 -7180 8280
rect -8352 7428 -7264 8252
rect -7200 7428 -7180 8252
rect -8352 7400 -7180 7428
rect -6940 8252 -5768 8280
rect -6940 7428 -5852 8252
rect -5788 7428 -5768 8252
rect -6940 7400 -5768 7428
rect -5528 8252 -4356 8280
rect -5528 7428 -4440 8252
rect -4376 7428 -4356 8252
rect -5528 7400 -4356 7428
rect -4116 8252 -2944 8280
rect -4116 7428 -3028 8252
rect -2964 7428 -2944 8252
rect -4116 7400 -2944 7428
rect -2704 8252 -1532 8280
rect -2704 7428 -1616 8252
rect -1552 7428 -1532 8252
rect -2704 7400 -1532 7428
rect -1292 8252 -120 8280
rect -1292 7428 -204 8252
rect -140 7428 -120 8252
rect -1292 7400 -120 7428
rect 120 8252 1292 8280
rect 120 7428 1208 8252
rect 1272 7428 1292 8252
rect 120 7400 1292 7428
rect 1532 8252 2704 8280
rect 1532 7428 2620 8252
rect 2684 7428 2704 8252
rect 1532 7400 2704 7428
rect 2944 8252 4116 8280
rect 2944 7428 4032 8252
rect 4096 7428 4116 8252
rect 2944 7400 4116 7428
rect 4356 8252 5528 8280
rect 4356 7428 5444 8252
rect 5508 7428 5528 8252
rect 4356 7400 5528 7428
rect 5768 8252 6940 8280
rect 5768 7428 6856 8252
rect 6920 7428 6940 8252
rect 5768 7400 6940 7428
rect 7180 8252 8352 8280
rect 7180 7428 8268 8252
rect 8332 7428 8352 8252
rect 7180 7400 8352 7428
rect 8592 8252 9764 8280
rect 8592 7428 9680 8252
rect 9744 7428 9764 8252
rect 8592 7400 9764 7428
rect 10004 8252 11176 8280
rect 10004 7428 11092 8252
rect 11156 7428 11176 8252
rect 10004 7400 11176 7428
rect 11416 8252 12588 8280
rect 11416 7428 12504 8252
rect 12568 7428 12588 8252
rect 11416 7400 12588 7428
rect 12828 8252 14000 8280
rect 12828 7428 13916 8252
rect 13980 7428 14000 8252
rect 12828 7400 14000 7428
rect 14240 8252 15412 8280
rect 14240 7428 15328 8252
rect 15392 7428 15412 8252
rect 14240 7400 15412 7428
rect 15652 8252 16824 8280
rect 15652 7428 16740 8252
rect 16804 7428 16824 8252
rect 15652 7400 16824 7428
rect 17064 8252 18236 8280
rect 17064 7428 18152 8252
rect 18216 7428 18236 8252
rect 17064 7400 18236 7428
rect 18476 8252 19648 8280
rect 18476 7428 19564 8252
rect 19628 7428 19648 8252
rect 18476 7400 19648 7428
rect 19888 8252 21060 8280
rect 19888 7428 20976 8252
rect 21040 7428 21060 8252
rect 19888 7400 21060 7428
rect 21300 8252 22472 8280
rect 21300 7428 22388 8252
rect 22452 7428 22472 8252
rect 21300 7400 22472 7428
rect 22712 8252 23884 8280
rect 22712 7428 23800 8252
rect 23864 7428 23884 8252
rect 22712 7400 23884 7428
rect -23884 7132 -22712 7160
rect -23884 6308 -22796 7132
rect -22732 6308 -22712 7132
rect -23884 6280 -22712 6308
rect -22472 7132 -21300 7160
rect -22472 6308 -21384 7132
rect -21320 6308 -21300 7132
rect -22472 6280 -21300 6308
rect -21060 7132 -19888 7160
rect -21060 6308 -19972 7132
rect -19908 6308 -19888 7132
rect -21060 6280 -19888 6308
rect -19648 7132 -18476 7160
rect -19648 6308 -18560 7132
rect -18496 6308 -18476 7132
rect -19648 6280 -18476 6308
rect -18236 7132 -17064 7160
rect -18236 6308 -17148 7132
rect -17084 6308 -17064 7132
rect -18236 6280 -17064 6308
rect -16824 7132 -15652 7160
rect -16824 6308 -15736 7132
rect -15672 6308 -15652 7132
rect -16824 6280 -15652 6308
rect -15412 7132 -14240 7160
rect -15412 6308 -14324 7132
rect -14260 6308 -14240 7132
rect -15412 6280 -14240 6308
rect -14000 7132 -12828 7160
rect -14000 6308 -12912 7132
rect -12848 6308 -12828 7132
rect -14000 6280 -12828 6308
rect -12588 7132 -11416 7160
rect -12588 6308 -11500 7132
rect -11436 6308 -11416 7132
rect -12588 6280 -11416 6308
rect -11176 7132 -10004 7160
rect -11176 6308 -10088 7132
rect -10024 6308 -10004 7132
rect -11176 6280 -10004 6308
rect -9764 7132 -8592 7160
rect -9764 6308 -8676 7132
rect -8612 6308 -8592 7132
rect -9764 6280 -8592 6308
rect -8352 7132 -7180 7160
rect -8352 6308 -7264 7132
rect -7200 6308 -7180 7132
rect -8352 6280 -7180 6308
rect -6940 7132 -5768 7160
rect -6940 6308 -5852 7132
rect -5788 6308 -5768 7132
rect -6940 6280 -5768 6308
rect -5528 7132 -4356 7160
rect -5528 6308 -4440 7132
rect -4376 6308 -4356 7132
rect -5528 6280 -4356 6308
rect -4116 7132 -2944 7160
rect -4116 6308 -3028 7132
rect -2964 6308 -2944 7132
rect -4116 6280 -2944 6308
rect -2704 7132 -1532 7160
rect -2704 6308 -1616 7132
rect -1552 6308 -1532 7132
rect -2704 6280 -1532 6308
rect -1292 7132 -120 7160
rect -1292 6308 -204 7132
rect -140 6308 -120 7132
rect -1292 6280 -120 6308
rect 120 7132 1292 7160
rect 120 6308 1208 7132
rect 1272 6308 1292 7132
rect 120 6280 1292 6308
rect 1532 7132 2704 7160
rect 1532 6308 2620 7132
rect 2684 6308 2704 7132
rect 1532 6280 2704 6308
rect 2944 7132 4116 7160
rect 2944 6308 4032 7132
rect 4096 6308 4116 7132
rect 2944 6280 4116 6308
rect 4356 7132 5528 7160
rect 4356 6308 5444 7132
rect 5508 6308 5528 7132
rect 4356 6280 5528 6308
rect 5768 7132 6940 7160
rect 5768 6308 6856 7132
rect 6920 6308 6940 7132
rect 5768 6280 6940 6308
rect 7180 7132 8352 7160
rect 7180 6308 8268 7132
rect 8332 6308 8352 7132
rect 7180 6280 8352 6308
rect 8592 7132 9764 7160
rect 8592 6308 9680 7132
rect 9744 6308 9764 7132
rect 8592 6280 9764 6308
rect 10004 7132 11176 7160
rect 10004 6308 11092 7132
rect 11156 6308 11176 7132
rect 10004 6280 11176 6308
rect 11416 7132 12588 7160
rect 11416 6308 12504 7132
rect 12568 6308 12588 7132
rect 11416 6280 12588 6308
rect 12828 7132 14000 7160
rect 12828 6308 13916 7132
rect 13980 6308 14000 7132
rect 12828 6280 14000 6308
rect 14240 7132 15412 7160
rect 14240 6308 15328 7132
rect 15392 6308 15412 7132
rect 14240 6280 15412 6308
rect 15652 7132 16824 7160
rect 15652 6308 16740 7132
rect 16804 6308 16824 7132
rect 15652 6280 16824 6308
rect 17064 7132 18236 7160
rect 17064 6308 18152 7132
rect 18216 6308 18236 7132
rect 17064 6280 18236 6308
rect 18476 7132 19648 7160
rect 18476 6308 19564 7132
rect 19628 6308 19648 7132
rect 18476 6280 19648 6308
rect 19888 7132 21060 7160
rect 19888 6308 20976 7132
rect 21040 6308 21060 7132
rect 19888 6280 21060 6308
rect 21300 7132 22472 7160
rect 21300 6308 22388 7132
rect 22452 6308 22472 7132
rect 21300 6280 22472 6308
rect 22712 7132 23884 7160
rect 22712 6308 23800 7132
rect 23864 6308 23884 7132
rect 22712 6280 23884 6308
rect -23884 6012 -22712 6040
rect -23884 5188 -22796 6012
rect -22732 5188 -22712 6012
rect -23884 5160 -22712 5188
rect -22472 6012 -21300 6040
rect -22472 5188 -21384 6012
rect -21320 5188 -21300 6012
rect -22472 5160 -21300 5188
rect -21060 6012 -19888 6040
rect -21060 5188 -19972 6012
rect -19908 5188 -19888 6012
rect -21060 5160 -19888 5188
rect -19648 6012 -18476 6040
rect -19648 5188 -18560 6012
rect -18496 5188 -18476 6012
rect -19648 5160 -18476 5188
rect -18236 6012 -17064 6040
rect -18236 5188 -17148 6012
rect -17084 5188 -17064 6012
rect -18236 5160 -17064 5188
rect -16824 6012 -15652 6040
rect -16824 5188 -15736 6012
rect -15672 5188 -15652 6012
rect -16824 5160 -15652 5188
rect -15412 6012 -14240 6040
rect -15412 5188 -14324 6012
rect -14260 5188 -14240 6012
rect -15412 5160 -14240 5188
rect -14000 6012 -12828 6040
rect -14000 5188 -12912 6012
rect -12848 5188 -12828 6012
rect -14000 5160 -12828 5188
rect -12588 6012 -11416 6040
rect -12588 5188 -11500 6012
rect -11436 5188 -11416 6012
rect -12588 5160 -11416 5188
rect -11176 6012 -10004 6040
rect -11176 5188 -10088 6012
rect -10024 5188 -10004 6012
rect -11176 5160 -10004 5188
rect -9764 6012 -8592 6040
rect -9764 5188 -8676 6012
rect -8612 5188 -8592 6012
rect -9764 5160 -8592 5188
rect -8352 6012 -7180 6040
rect -8352 5188 -7264 6012
rect -7200 5188 -7180 6012
rect -8352 5160 -7180 5188
rect -6940 6012 -5768 6040
rect -6940 5188 -5852 6012
rect -5788 5188 -5768 6012
rect -6940 5160 -5768 5188
rect -5528 6012 -4356 6040
rect -5528 5188 -4440 6012
rect -4376 5188 -4356 6012
rect -5528 5160 -4356 5188
rect -4116 6012 -2944 6040
rect -4116 5188 -3028 6012
rect -2964 5188 -2944 6012
rect -4116 5160 -2944 5188
rect -2704 6012 -1532 6040
rect -2704 5188 -1616 6012
rect -1552 5188 -1532 6012
rect -2704 5160 -1532 5188
rect -1292 6012 -120 6040
rect -1292 5188 -204 6012
rect -140 5188 -120 6012
rect -1292 5160 -120 5188
rect 120 6012 1292 6040
rect 120 5188 1208 6012
rect 1272 5188 1292 6012
rect 120 5160 1292 5188
rect 1532 6012 2704 6040
rect 1532 5188 2620 6012
rect 2684 5188 2704 6012
rect 1532 5160 2704 5188
rect 2944 6012 4116 6040
rect 2944 5188 4032 6012
rect 4096 5188 4116 6012
rect 2944 5160 4116 5188
rect 4356 6012 5528 6040
rect 4356 5188 5444 6012
rect 5508 5188 5528 6012
rect 4356 5160 5528 5188
rect 5768 6012 6940 6040
rect 5768 5188 6856 6012
rect 6920 5188 6940 6012
rect 5768 5160 6940 5188
rect 7180 6012 8352 6040
rect 7180 5188 8268 6012
rect 8332 5188 8352 6012
rect 7180 5160 8352 5188
rect 8592 6012 9764 6040
rect 8592 5188 9680 6012
rect 9744 5188 9764 6012
rect 8592 5160 9764 5188
rect 10004 6012 11176 6040
rect 10004 5188 11092 6012
rect 11156 5188 11176 6012
rect 10004 5160 11176 5188
rect 11416 6012 12588 6040
rect 11416 5188 12504 6012
rect 12568 5188 12588 6012
rect 11416 5160 12588 5188
rect 12828 6012 14000 6040
rect 12828 5188 13916 6012
rect 13980 5188 14000 6012
rect 12828 5160 14000 5188
rect 14240 6012 15412 6040
rect 14240 5188 15328 6012
rect 15392 5188 15412 6012
rect 14240 5160 15412 5188
rect 15652 6012 16824 6040
rect 15652 5188 16740 6012
rect 16804 5188 16824 6012
rect 15652 5160 16824 5188
rect 17064 6012 18236 6040
rect 17064 5188 18152 6012
rect 18216 5188 18236 6012
rect 17064 5160 18236 5188
rect 18476 6012 19648 6040
rect 18476 5188 19564 6012
rect 19628 5188 19648 6012
rect 18476 5160 19648 5188
rect 19888 6012 21060 6040
rect 19888 5188 20976 6012
rect 21040 5188 21060 6012
rect 19888 5160 21060 5188
rect 21300 6012 22472 6040
rect 21300 5188 22388 6012
rect 22452 5188 22472 6012
rect 21300 5160 22472 5188
rect 22712 6012 23884 6040
rect 22712 5188 23800 6012
rect 23864 5188 23884 6012
rect 22712 5160 23884 5188
rect -23884 4892 -22712 4920
rect -23884 4068 -22796 4892
rect -22732 4068 -22712 4892
rect -23884 4040 -22712 4068
rect -22472 4892 -21300 4920
rect -22472 4068 -21384 4892
rect -21320 4068 -21300 4892
rect -22472 4040 -21300 4068
rect -21060 4892 -19888 4920
rect -21060 4068 -19972 4892
rect -19908 4068 -19888 4892
rect -21060 4040 -19888 4068
rect -19648 4892 -18476 4920
rect -19648 4068 -18560 4892
rect -18496 4068 -18476 4892
rect -19648 4040 -18476 4068
rect -18236 4892 -17064 4920
rect -18236 4068 -17148 4892
rect -17084 4068 -17064 4892
rect -18236 4040 -17064 4068
rect -16824 4892 -15652 4920
rect -16824 4068 -15736 4892
rect -15672 4068 -15652 4892
rect -16824 4040 -15652 4068
rect -15412 4892 -14240 4920
rect -15412 4068 -14324 4892
rect -14260 4068 -14240 4892
rect -15412 4040 -14240 4068
rect -14000 4892 -12828 4920
rect -14000 4068 -12912 4892
rect -12848 4068 -12828 4892
rect -14000 4040 -12828 4068
rect -12588 4892 -11416 4920
rect -12588 4068 -11500 4892
rect -11436 4068 -11416 4892
rect -12588 4040 -11416 4068
rect -11176 4892 -10004 4920
rect -11176 4068 -10088 4892
rect -10024 4068 -10004 4892
rect -11176 4040 -10004 4068
rect -9764 4892 -8592 4920
rect -9764 4068 -8676 4892
rect -8612 4068 -8592 4892
rect -9764 4040 -8592 4068
rect -8352 4892 -7180 4920
rect -8352 4068 -7264 4892
rect -7200 4068 -7180 4892
rect -8352 4040 -7180 4068
rect -6940 4892 -5768 4920
rect -6940 4068 -5852 4892
rect -5788 4068 -5768 4892
rect -6940 4040 -5768 4068
rect -5528 4892 -4356 4920
rect -5528 4068 -4440 4892
rect -4376 4068 -4356 4892
rect -5528 4040 -4356 4068
rect -4116 4892 -2944 4920
rect -4116 4068 -3028 4892
rect -2964 4068 -2944 4892
rect -4116 4040 -2944 4068
rect -2704 4892 -1532 4920
rect -2704 4068 -1616 4892
rect -1552 4068 -1532 4892
rect -2704 4040 -1532 4068
rect -1292 4892 -120 4920
rect -1292 4068 -204 4892
rect -140 4068 -120 4892
rect -1292 4040 -120 4068
rect 120 4892 1292 4920
rect 120 4068 1208 4892
rect 1272 4068 1292 4892
rect 120 4040 1292 4068
rect 1532 4892 2704 4920
rect 1532 4068 2620 4892
rect 2684 4068 2704 4892
rect 1532 4040 2704 4068
rect 2944 4892 4116 4920
rect 2944 4068 4032 4892
rect 4096 4068 4116 4892
rect 2944 4040 4116 4068
rect 4356 4892 5528 4920
rect 4356 4068 5444 4892
rect 5508 4068 5528 4892
rect 4356 4040 5528 4068
rect 5768 4892 6940 4920
rect 5768 4068 6856 4892
rect 6920 4068 6940 4892
rect 5768 4040 6940 4068
rect 7180 4892 8352 4920
rect 7180 4068 8268 4892
rect 8332 4068 8352 4892
rect 7180 4040 8352 4068
rect 8592 4892 9764 4920
rect 8592 4068 9680 4892
rect 9744 4068 9764 4892
rect 8592 4040 9764 4068
rect 10004 4892 11176 4920
rect 10004 4068 11092 4892
rect 11156 4068 11176 4892
rect 10004 4040 11176 4068
rect 11416 4892 12588 4920
rect 11416 4068 12504 4892
rect 12568 4068 12588 4892
rect 11416 4040 12588 4068
rect 12828 4892 14000 4920
rect 12828 4068 13916 4892
rect 13980 4068 14000 4892
rect 12828 4040 14000 4068
rect 14240 4892 15412 4920
rect 14240 4068 15328 4892
rect 15392 4068 15412 4892
rect 14240 4040 15412 4068
rect 15652 4892 16824 4920
rect 15652 4068 16740 4892
rect 16804 4068 16824 4892
rect 15652 4040 16824 4068
rect 17064 4892 18236 4920
rect 17064 4068 18152 4892
rect 18216 4068 18236 4892
rect 17064 4040 18236 4068
rect 18476 4892 19648 4920
rect 18476 4068 19564 4892
rect 19628 4068 19648 4892
rect 18476 4040 19648 4068
rect 19888 4892 21060 4920
rect 19888 4068 20976 4892
rect 21040 4068 21060 4892
rect 19888 4040 21060 4068
rect 21300 4892 22472 4920
rect 21300 4068 22388 4892
rect 22452 4068 22472 4892
rect 21300 4040 22472 4068
rect 22712 4892 23884 4920
rect 22712 4068 23800 4892
rect 23864 4068 23884 4892
rect 22712 4040 23884 4068
rect -23884 3772 -22712 3800
rect -23884 2948 -22796 3772
rect -22732 2948 -22712 3772
rect -23884 2920 -22712 2948
rect -22472 3772 -21300 3800
rect -22472 2948 -21384 3772
rect -21320 2948 -21300 3772
rect -22472 2920 -21300 2948
rect -21060 3772 -19888 3800
rect -21060 2948 -19972 3772
rect -19908 2948 -19888 3772
rect -21060 2920 -19888 2948
rect -19648 3772 -18476 3800
rect -19648 2948 -18560 3772
rect -18496 2948 -18476 3772
rect -19648 2920 -18476 2948
rect -18236 3772 -17064 3800
rect -18236 2948 -17148 3772
rect -17084 2948 -17064 3772
rect -18236 2920 -17064 2948
rect -16824 3772 -15652 3800
rect -16824 2948 -15736 3772
rect -15672 2948 -15652 3772
rect -16824 2920 -15652 2948
rect -15412 3772 -14240 3800
rect -15412 2948 -14324 3772
rect -14260 2948 -14240 3772
rect -15412 2920 -14240 2948
rect -14000 3772 -12828 3800
rect -14000 2948 -12912 3772
rect -12848 2948 -12828 3772
rect -14000 2920 -12828 2948
rect -12588 3772 -11416 3800
rect -12588 2948 -11500 3772
rect -11436 2948 -11416 3772
rect -12588 2920 -11416 2948
rect -11176 3772 -10004 3800
rect -11176 2948 -10088 3772
rect -10024 2948 -10004 3772
rect -11176 2920 -10004 2948
rect -9764 3772 -8592 3800
rect -9764 2948 -8676 3772
rect -8612 2948 -8592 3772
rect -9764 2920 -8592 2948
rect -8352 3772 -7180 3800
rect -8352 2948 -7264 3772
rect -7200 2948 -7180 3772
rect -8352 2920 -7180 2948
rect -6940 3772 -5768 3800
rect -6940 2948 -5852 3772
rect -5788 2948 -5768 3772
rect -6940 2920 -5768 2948
rect -5528 3772 -4356 3800
rect -5528 2948 -4440 3772
rect -4376 2948 -4356 3772
rect -5528 2920 -4356 2948
rect -4116 3772 -2944 3800
rect -4116 2948 -3028 3772
rect -2964 2948 -2944 3772
rect -4116 2920 -2944 2948
rect -2704 3772 -1532 3800
rect -2704 2948 -1616 3772
rect -1552 2948 -1532 3772
rect -2704 2920 -1532 2948
rect -1292 3772 -120 3800
rect -1292 2948 -204 3772
rect -140 2948 -120 3772
rect -1292 2920 -120 2948
rect 120 3772 1292 3800
rect 120 2948 1208 3772
rect 1272 2948 1292 3772
rect 120 2920 1292 2948
rect 1532 3772 2704 3800
rect 1532 2948 2620 3772
rect 2684 2948 2704 3772
rect 1532 2920 2704 2948
rect 2944 3772 4116 3800
rect 2944 2948 4032 3772
rect 4096 2948 4116 3772
rect 2944 2920 4116 2948
rect 4356 3772 5528 3800
rect 4356 2948 5444 3772
rect 5508 2948 5528 3772
rect 4356 2920 5528 2948
rect 5768 3772 6940 3800
rect 5768 2948 6856 3772
rect 6920 2948 6940 3772
rect 5768 2920 6940 2948
rect 7180 3772 8352 3800
rect 7180 2948 8268 3772
rect 8332 2948 8352 3772
rect 7180 2920 8352 2948
rect 8592 3772 9764 3800
rect 8592 2948 9680 3772
rect 9744 2948 9764 3772
rect 8592 2920 9764 2948
rect 10004 3772 11176 3800
rect 10004 2948 11092 3772
rect 11156 2948 11176 3772
rect 10004 2920 11176 2948
rect 11416 3772 12588 3800
rect 11416 2948 12504 3772
rect 12568 2948 12588 3772
rect 11416 2920 12588 2948
rect 12828 3772 14000 3800
rect 12828 2948 13916 3772
rect 13980 2948 14000 3772
rect 12828 2920 14000 2948
rect 14240 3772 15412 3800
rect 14240 2948 15328 3772
rect 15392 2948 15412 3772
rect 14240 2920 15412 2948
rect 15652 3772 16824 3800
rect 15652 2948 16740 3772
rect 16804 2948 16824 3772
rect 15652 2920 16824 2948
rect 17064 3772 18236 3800
rect 17064 2948 18152 3772
rect 18216 2948 18236 3772
rect 17064 2920 18236 2948
rect 18476 3772 19648 3800
rect 18476 2948 19564 3772
rect 19628 2948 19648 3772
rect 18476 2920 19648 2948
rect 19888 3772 21060 3800
rect 19888 2948 20976 3772
rect 21040 2948 21060 3772
rect 19888 2920 21060 2948
rect 21300 3772 22472 3800
rect 21300 2948 22388 3772
rect 22452 2948 22472 3772
rect 21300 2920 22472 2948
rect 22712 3772 23884 3800
rect 22712 2948 23800 3772
rect 23864 2948 23884 3772
rect 22712 2920 23884 2948
rect -23884 2652 -22712 2680
rect -23884 1828 -22796 2652
rect -22732 1828 -22712 2652
rect -23884 1800 -22712 1828
rect -22472 2652 -21300 2680
rect -22472 1828 -21384 2652
rect -21320 1828 -21300 2652
rect -22472 1800 -21300 1828
rect -21060 2652 -19888 2680
rect -21060 1828 -19972 2652
rect -19908 1828 -19888 2652
rect -21060 1800 -19888 1828
rect -19648 2652 -18476 2680
rect -19648 1828 -18560 2652
rect -18496 1828 -18476 2652
rect -19648 1800 -18476 1828
rect -18236 2652 -17064 2680
rect -18236 1828 -17148 2652
rect -17084 1828 -17064 2652
rect -18236 1800 -17064 1828
rect -16824 2652 -15652 2680
rect -16824 1828 -15736 2652
rect -15672 1828 -15652 2652
rect -16824 1800 -15652 1828
rect -15412 2652 -14240 2680
rect -15412 1828 -14324 2652
rect -14260 1828 -14240 2652
rect -15412 1800 -14240 1828
rect -14000 2652 -12828 2680
rect -14000 1828 -12912 2652
rect -12848 1828 -12828 2652
rect -14000 1800 -12828 1828
rect -12588 2652 -11416 2680
rect -12588 1828 -11500 2652
rect -11436 1828 -11416 2652
rect -12588 1800 -11416 1828
rect -11176 2652 -10004 2680
rect -11176 1828 -10088 2652
rect -10024 1828 -10004 2652
rect -11176 1800 -10004 1828
rect -9764 2652 -8592 2680
rect -9764 1828 -8676 2652
rect -8612 1828 -8592 2652
rect -9764 1800 -8592 1828
rect -8352 2652 -7180 2680
rect -8352 1828 -7264 2652
rect -7200 1828 -7180 2652
rect -8352 1800 -7180 1828
rect -6940 2652 -5768 2680
rect -6940 1828 -5852 2652
rect -5788 1828 -5768 2652
rect -6940 1800 -5768 1828
rect -5528 2652 -4356 2680
rect -5528 1828 -4440 2652
rect -4376 1828 -4356 2652
rect -5528 1800 -4356 1828
rect -4116 2652 -2944 2680
rect -4116 1828 -3028 2652
rect -2964 1828 -2944 2652
rect -4116 1800 -2944 1828
rect -2704 2652 -1532 2680
rect -2704 1828 -1616 2652
rect -1552 1828 -1532 2652
rect -2704 1800 -1532 1828
rect -1292 2652 -120 2680
rect -1292 1828 -204 2652
rect -140 1828 -120 2652
rect -1292 1800 -120 1828
rect 120 2652 1292 2680
rect 120 1828 1208 2652
rect 1272 1828 1292 2652
rect 120 1800 1292 1828
rect 1532 2652 2704 2680
rect 1532 1828 2620 2652
rect 2684 1828 2704 2652
rect 1532 1800 2704 1828
rect 2944 2652 4116 2680
rect 2944 1828 4032 2652
rect 4096 1828 4116 2652
rect 2944 1800 4116 1828
rect 4356 2652 5528 2680
rect 4356 1828 5444 2652
rect 5508 1828 5528 2652
rect 4356 1800 5528 1828
rect 5768 2652 6940 2680
rect 5768 1828 6856 2652
rect 6920 1828 6940 2652
rect 5768 1800 6940 1828
rect 7180 2652 8352 2680
rect 7180 1828 8268 2652
rect 8332 1828 8352 2652
rect 7180 1800 8352 1828
rect 8592 2652 9764 2680
rect 8592 1828 9680 2652
rect 9744 1828 9764 2652
rect 8592 1800 9764 1828
rect 10004 2652 11176 2680
rect 10004 1828 11092 2652
rect 11156 1828 11176 2652
rect 10004 1800 11176 1828
rect 11416 2652 12588 2680
rect 11416 1828 12504 2652
rect 12568 1828 12588 2652
rect 11416 1800 12588 1828
rect 12828 2652 14000 2680
rect 12828 1828 13916 2652
rect 13980 1828 14000 2652
rect 12828 1800 14000 1828
rect 14240 2652 15412 2680
rect 14240 1828 15328 2652
rect 15392 1828 15412 2652
rect 14240 1800 15412 1828
rect 15652 2652 16824 2680
rect 15652 1828 16740 2652
rect 16804 1828 16824 2652
rect 15652 1800 16824 1828
rect 17064 2652 18236 2680
rect 17064 1828 18152 2652
rect 18216 1828 18236 2652
rect 17064 1800 18236 1828
rect 18476 2652 19648 2680
rect 18476 1828 19564 2652
rect 19628 1828 19648 2652
rect 18476 1800 19648 1828
rect 19888 2652 21060 2680
rect 19888 1828 20976 2652
rect 21040 1828 21060 2652
rect 19888 1800 21060 1828
rect 21300 2652 22472 2680
rect 21300 1828 22388 2652
rect 22452 1828 22472 2652
rect 21300 1800 22472 1828
rect 22712 2652 23884 2680
rect 22712 1828 23800 2652
rect 23864 1828 23884 2652
rect 22712 1800 23884 1828
rect -23884 1532 -22712 1560
rect -23884 708 -22796 1532
rect -22732 708 -22712 1532
rect -23884 680 -22712 708
rect -22472 1532 -21300 1560
rect -22472 708 -21384 1532
rect -21320 708 -21300 1532
rect -22472 680 -21300 708
rect -21060 1532 -19888 1560
rect -21060 708 -19972 1532
rect -19908 708 -19888 1532
rect -21060 680 -19888 708
rect -19648 1532 -18476 1560
rect -19648 708 -18560 1532
rect -18496 708 -18476 1532
rect -19648 680 -18476 708
rect -18236 1532 -17064 1560
rect -18236 708 -17148 1532
rect -17084 708 -17064 1532
rect -18236 680 -17064 708
rect -16824 1532 -15652 1560
rect -16824 708 -15736 1532
rect -15672 708 -15652 1532
rect -16824 680 -15652 708
rect -15412 1532 -14240 1560
rect -15412 708 -14324 1532
rect -14260 708 -14240 1532
rect -15412 680 -14240 708
rect -14000 1532 -12828 1560
rect -14000 708 -12912 1532
rect -12848 708 -12828 1532
rect -14000 680 -12828 708
rect -12588 1532 -11416 1560
rect -12588 708 -11500 1532
rect -11436 708 -11416 1532
rect -12588 680 -11416 708
rect -11176 1532 -10004 1560
rect -11176 708 -10088 1532
rect -10024 708 -10004 1532
rect -11176 680 -10004 708
rect -9764 1532 -8592 1560
rect -9764 708 -8676 1532
rect -8612 708 -8592 1532
rect -9764 680 -8592 708
rect -8352 1532 -7180 1560
rect -8352 708 -7264 1532
rect -7200 708 -7180 1532
rect -8352 680 -7180 708
rect -6940 1532 -5768 1560
rect -6940 708 -5852 1532
rect -5788 708 -5768 1532
rect -6940 680 -5768 708
rect -5528 1532 -4356 1560
rect -5528 708 -4440 1532
rect -4376 708 -4356 1532
rect -5528 680 -4356 708
rect -4116 1532 -2944 1560
rect -4116 708 -3028 1532
rect -2964 708 -2944 1532
rect -4116 680 -2944 708
rect -2704 1532 -1532 1560
rect -2704 708 -1616 1532
rect -1552 708 -1532 1532
rect -2704 680 -1532 708
rect -1292 1532 -120 1560
rect -1292 708 -204 1532
rect -140 708 -120 1532
rect -1292 680 -120 708
rect 120 1532 1292 1560
rect 120 708 1208 1532
rect 1272 708 1292 1532
rect 120 680 1292 708
rect 1532 1532 2704 1560
rect 1532 708 2620 1532
rect 2684 708 2704 1532
rect 1532 680 2704 708
rect 2944 1532 4116 1560
rect 2944 708 4032 1532
rect 4096 708 4116 1532
rect 2944 680 4116 708
rect 4356 1532 5528 1560
rect 4356 708 5444 1532
rect 5508 708 5528 1532
rect 4356 680 5528 708
rect 5768 1532 6940 1560
rect 5768 708 6856 1532
rect 6920 708 6940 1532
rect 5768 680 6940 708
rect 7180 1532 8352 1560
rect 7180 708 8268 1532
rect 8332 708 8352 1532
rect 7180 680 8352 708
rect 8592 1532 9764 1560
rect 8592 708 9680 1532
rect 9744 708 9764 1532
rect 8592 680 9764 708
rect 10004 1532 11176 1560
rect 10004 708 11092 1532
rect 11156 708 11176 1532
rect 10004 680 11176 708
rect 11416 1532 12588 1560
rect 11416 708 12504 1532
rect 12568 708 12588 1532
rect 11416 680 12588 708
rect 12828 1532 14000 1560
rect 12828 708 13916 1532
rect 13980 708 14000 1532
rect 12828 680 14000 708
rect 14240 1532 15412 1560
rect 14240 708 15328 1532
rect 15392 708 15412 1532
rect 14240 680 15412 708
rect 15652 1532 16824 1560
rect 15652 708 16740 1532
rect 16804 708 16824 1532
rect 15652 680 16824 708
rect 17064 1532 18236 1560
rect 17064 708 18152 1532
rect 18216 708 18236 1532
rect 17064 680 18236 708
rect 18476 1532 19648 1560
rect 18476 708 19564 1532
rect 19628 708 19648 1532
rect 18476 680 19648 708
rect 19888 1532 21060 1560
rect 19888 708 20976 1532
rect 21040 708 21060 1532
rect 19888 680 21060 708
rect 21300 1532 22472 1560
rect 21300 708 22388 1532
rect 22452 708 22472 1532
rect 21300 680 22472 708
rect 22712 1532 23884 1560
rect 22712 708 23800 1532
rect 23864 708 23884 1532
rect 22712 680 23884 708
rect -23884 412 -22712 440
rect -23884 -412 -22796 412
rect -22732 -412 -22712 412
rect -23884 -440 -22712 -412
rect -22472 412 -21300 440
rect -22472 -412 -21384 412
rect -21320 -412 -21300 412
rect -22472 -440 -21300 -412
rect -21060 412 -19888 440
rect -21060 -412 -19972 412
rect -19908 -412 -19888 412
rect -21060 -440 -19888 -412
rect -19648 412 -18476 440
rect -19648 -412 -18560 412
rect -18496 -412 -18476 412
rect -19648 -440 -18476 -412
rect -18236 412 -17064 440
rect -18236 -412 -17148 412
rect -17084 -412 -17064 412
rect -18236 -440 -17064 -412
rect -16824 412 -15652 440
rect -16824 -412 -15736 412
rect -15672 -412 -15652 412
rect -16824 -440 -15652 -412
rect -15412 412 -14240 440
rect -15412 -412 -14324 412
rect -14260 -412 -14240 412
rect -15412 -440 -14240 -412
rect -14000 412 -12828 440
rect -14000 -412 -12912 412
rect -12848 -412 -12828 412
rect -14000 -440 -12828 -412
rect -12588 412 -11416 440
rect -12588 -412 -11500 412
rect -11436 -412 -11416 412
rect -12588 -440 -11416 -412
rect -11176 412 -10004 440
rect -11176 -412 -10088 412
rect -10024 -412 -10004 412
rect -11176 -440 -10004 -412
rect -9764 412 -8592 440
rect -9764 -412 -8676 412
rect -8612 -412 -8592 412
rect -9764 -440 -8592 -412
rect -8352 412 -7180 440
rect -8352 -412 -7264 412
rect -7200 -412 -7180 412
rect -8352 -440 -7180 -412
rect -6940 412 -5768 440
rect -6940 -412 -5852 412
rect -5788 -412 -5768 412
rect -6940 -440 -5768 -412
rect -5528 412 -4356 440
rect -5528 -412 -4440 412
rect -4376 -412 -4356 412
rect -5528 -440 -4356 -412
rect -4116 412 -2944 440
rect -4116 -412 -3028 412
rect -2964 -412 -2944 412
rect -4116 -440 -2944 -412
rect -2704 412 -1532 440
rect -2704 -412 -1616 412
rect -1552 -412 -1532 412
rect -2704 -440 -1532 -412
rect -1292 412 -120 440
rect -1292 -412 -204 412
rect -140 -412 -120 412
rect -1292 -440 -120 -412
rect 120 412 1292 440
rect 120 -412 1208 412
rect 1272 -412 1292 412
rect 120 -440 1292 -412
rect 1532 412 2704 440
rect 1532 -412 2620 412
rect 2684 -412 2704 412
rect 1532 -440 2704 -412
rect 2944 412 4116 440
rect 2944 -412 4032 412
rect 4096 -412 4116 412
rect 2944 -440 4116 -412
rect 4356 412 5528 440
rect 4356 -412 5444 412
rect 5508 -412 5528 412
rect 4356 -440 5528 -412
rect 5768 412 6940 440
rect 5768 -412 6856 412
rect 6920 -412 6940 412
rect 5768 -440 6940 -412
rect 7180 412 8352 440
rect 7180 -412 8268 412
rect 8332 -412 8352 412
rect 7180 -440 8352 -412
rect 8592 412 9764 440
rect 8592 -412 9680 412
rect 9744 -412 9764 412
rect 8592 -440 9764 -412
rect 10004 412 11176 440
rect 10004 -412 11092 412
rect 11156 -412 11176 412
rect 10004 -440 11176 -412
rect 11416 412 12588 440
rect 11416 -412 12504 412
rect 12568 -412 12588 412
rect 11416 -440 12588 -412
rect 12828 412 14000 440
rect 12828 -412 13916 412
rect 13980 -412 14000 412
rect 12828 -440 14000 -412
rect 14240 412 15412 440
rect 14240 -412 15328 412
rect 15392 -412 15412 412
rect 14240 -440 15412 -412
rect 15652 412 16824 440
rect 15652 -412 16740 412
rect 16804 -412 16824 412
rect 15652 -440 16824 -412
rect 17064 412 18236 440
rect 17064 -412 18152 412
rect 18216 -412 18236 412
rect 17064 -440 18236 -412
rect 18476 412 19648 440
rect 18476 -412 19564 412
rect 19628 -412 19648 412
rect 18476 -440 19648 -412
rect 19888 412 21060 440
rect 19888 -412 20976 412
rect 21040 -412 21060 412
rect 19888 -440 21060 -412
rect 21300 412 22472 440
rect 21300 -412 22388 412
rect 22452 -412 22472 412
rect 21300 -440 22472 -412
rect 22712 412 23884 440
rect 22712 -412 23800 412
rect 23864 -412 23884 412
rect 22712 -440 23884 -412
rect -23884 -708 -22712 -680
rect -23884 -1532 -22796 -708
rect -22732 -1532 -22712 -708
rect -23884 -1560 -22712 -1532
rect -22472 -708 -21300 -680
rect -22472 -1532 -21384 -708
rect -21320 -1532 -21300 -708
rect -22472 -1560 -21300 -1532
rect -21060 -708 -19888 -680
rect -21060 -1532 -19972 -708
rect -19908 -1532 -19888 -708
rect -21060 -1560 -19888 -1532
rect -19648 -708 -18476 -680
rect -19648 -1532 -18560 -708
rect -18496 -1532 -18476 -708
rect -19648 -1560 -18476 -1532
rect -18236 -708 -17064 -680
rect -18236 -1532 -17148 -708
rect -17084 -1532 -17064 -708
rect -18236 -1560 -17064 -1532
rect -16824 -708 -15652 -680
rect -16824 -1532 -15736 -708
rect -15672 -1532 -15652 -708
rect -16824 -1560 -15652 -1532
rect -15412 -708 -14240 -680
rect -15412 -1532 -14324 -708
rect -14260 -1532 -14240 -708
rect -15412 -1560 -14240 -1532
rect -14000 -708 -12828 -680
rect -14000 -1532 -12912 -708
rect -12848 -1532 -12828 -708
rect -14000 -1560 -12828 -1532
rect -12588 -708 -11416 -680
rect -12588 -1532 -11500 -708
rect -11436 -1532 -11416 -708
rect -12588 -1560 -11416 -1532
rect -11176 -708 -10004 -680
rect -11176 -1532 -10088 -708
rect -10024 -1532 -10004 -708
rect -11176 -1560 -10004 -1532
rect -9764 -708 -8592 -680
rect -9764 -1532 -8676 -708
rect -8612 -1532 -8592 -708
rect -9764 -1560 -8592 -1532
rect -8352 -708 -7180 -680
rect -8352 -1532 -7264 -708
rect -7200 -1532 -7180 -708
rect -8352 -1560 -7180 -1532
rect -6940 -708 -5768 -680
rect -6940 -1532 -5852 -708
rect -5788 -1532 -5768 -708
rect -6940 -1560 -5768 -1532
rect -5528 -708 -4356 -680
rect -5528 -1532 -4440 -708
rect -4376 -1532 -4356 -708
rect -5528 -1560 -4356 -1532
rect -4116 -708 -2944 -680
rect -4116 -1532 -3028 -708
rect -2964 -1532 -2944 -708
rect -4116 -1560 -2944 -1532
rect -2704 -708 -1532 -680
rect -2704 -1532 -1616 -708
rect -1552 -1532 -1532 -708
rect -2704 -1560 -1532 -1532
rect -1292 -708 -120 -680
rect -1292 -1532 -204 -708
rect -140 -1532 -120 -708
rect -1292 -1560 -120 -1532
rect 120 -708 1292 -680
rect 120 -1532 1208 -708
rect 1272 -1532 1292 -708
rect 120 -1560 1292 -1532
rect 1532 -708 2704 -680
rect 1532 -1532 2620 -708
rect 2684 -1532 2704 -708
rect 1532 -1560 2704 -1532
rect 2944 -708 4116 -680
rect 2944 -1532 4032 -708
rect 4096 -1532 4116 -708
rect 2944 -1560 4116 -1532
rect 4356 -708 5528 -680
rect 4356 -1532 5444 -708
rect 5508 -1532 5528 -708
rect 4356 -1560 5528 -1532
rect 5768 -708 6940 -680
rect 5768 -1532 6856 -708
rect 6920 -1532 6940 -708
rect 5768 -1560 6940 -1532
rect 7180 -708 8352 -680
rect 7180 -1532 8268 -708
rect 8332 -1532 8352 -708
rect 7180 -1560 8352 -1532
rect 8592 -708 9764 -680
rect 8592 -1532 9680 -708
rect 9744 -1532 9764 -708
rect 8592 -1560 9764 -1532
rect 10004 -708 11176 -680
rect 10004 -1532 11092 -708
rect 11156 -1532 11176 -708
rect 10004 -1560 11176 -1532
rect 11416 -708 12588 -680
rect 11416 -1532 12504 -708
rect 12568 -1532 12588 -708
rect 11416 -1560 12588 -1532
rect 12828 -708 14000 -680
rect 12828 -1532 13916 -708
rect 13980 -1532 14000 -708
rect 12828 -1560 14000 -1532
rect 14240 -708 15412 -680
rect 14240 -1532 15328 -708
rect 15392 -1532 15412 -708
rect 14240 -1560 15412 -1532
rect 15652 -708 16824 -680
rect 15652 -1532 16740 -708
rect 16804 -1532 16824 -708
rect 15652 -1560 16824 -1532
rect 17064 -708 18236 -680
rect 17064 -1532 18152 -708
rect 18216 -1532 18236 -708
rect 17064 -1560 18236 -1532
rect 18476 -708 19648 -680
rect 18476 -1532 19564 -708
rect 19628 -1532 19648 -708
rect 18476 -1560 19648 -1532
rect 19888 -708 21060 -680
rect 19888 -1532 20976 -708
rect 21040 -1532 21060 -708
rect 19888 -1560 21060 -1532
rect 21300 -708 22472 -680
rect 21300 -1532 22388 -708
rect 22452 -1532 22472 -708
rect 21300 -1560 22472 -1532
rect 22712 -708 23884 -680
rect 22712 -1532 23800 -708
rect 23864 -1532 23884 -708
rect 22712 -1560 23884 -1532
rect -23884 -1828 -22712 -1800
rect -23884 -2652 -22796 -1828
rect -22732 -2652 -22712 -1828
rect -23884 -2680 -22712 -2652
rect -22472 -1828 -21300 -1800
rect -22472 -2652 -21384 -1828
rect -21320 -2652 -21300 -1828
rect -22472 -2680 -21300 -2652
rect -21060 -1828 -19888 -1800
rect -21060 -2652 -19972 -1828
rect -19908 -2652 -19888 -1828
rect -21060 -2680 -19888 -2652
rect -19648 -1828 -18476 -1800
rect -19648 -2652 -18560 -1828
rect -18496 -2652 -18476 -1828
rect -19648 -2680 -18476 -2652
rect -18236 -1828 -17064 -1800
rect -18236 -2652 -17148 -1828
rect -17084 -2652 -17064 -1828
rect -18236 -2680 -17064 -2652
rect -16824 -1828 -15652 -1800
rect -16824 -2652 -15736 -1828
rect -15672 -2652 -15652 -1828
rect -16824 -2680 -15652 -2652
rect -15412 -1828 -14240 -1800
rect -15412 -2652 -14324 -1828
rect -14260 -2652 -14240 -1828
rect -15412 -2680 -14240 -2652
rect -14000 -1828 -12828 -1800
rect -14000 -2652 -12912 -1828
rect -12848 -2652 -12828 -1828
rect -14000 -2680 -12828 -2652
rect -12588 -1828 -11416 -1800
rect -12588 -2652 -11500 -1828
rect -11436 -2652 -11416 -1828
rect -12588 -2680 -11416 -2652
rect -11176 -1828 -10004 -1800
rect -11176 -2652 -10088 -1828
rect -10024 -2652 -10004 -1828
rect -11176 -2680 -10004 -2652
rect -9764 -1828 -8592 -1800
rect -9764 -2652 -8676 -1828
rect -8612 -2652 -8592 -1828
rect -9764 -2680 -8592 -2652
rect -8352 -1828 -7180 -1800
rect -8352 -2652 -7264 -1828
rect -7200 -2652 -7180 -1828
rect -8352 -2680 -7180 -2652
rect -6940 -1828 -5768 -1800
rect -6940 -2652 -5852 -1828
rect -5788 -2652 -5768 -1828
rect -6940 -2680 -5768 -2652
rect -5528 -1828 -4356 -1800
rect -5528 -2652 -4440 -1828
rect -4376 -2652 -4356 -1828
rect -5528 -2680 -4356 -2652
rect -4116 -1828 -2944 -1800
rect -4116 -2652 -3028 -1828
rect -2964 -2652 -2944 -1828
rect -4116 -2680 -2944 -2652
rect -2704 -1828 -1532 -1800
rect -2704 -2652 -1616 -1828
rect -1552 -2652 -1532 -1828
rect -2704 -2680 -1532 -2652
rect -1292 -1828 -120 -1800
rect -1292 -2652 -204 -1828
rect -140 -2652 -120 -1828
rect -1292 -2680 -120 -2652
rect 120 -1828 1292 -1800
rect 120 -2652 1208 -1828
rect 1272 -2652 1292 -1828
rect 120 -2680 1292 -2652
rect 1532 -1828 2704 -1800
rect 1532 -2652 2620 -1828
rect 2684 -2652 2704 -1828
rect 1532 -2680 2704 -2652
rect 2944 -1828 4116 -1800
rect 2944 -2652 4032 -1828
rect 4096 -2652 4116 -1828
rect 2944 -2680 4116 -2652
rect 4356 -1828 5528 -1800
rect 4356 -2652 5444 -1828
rect 5508 -2652 5528 -1828
rect 4356 -2680 5528 -2652
rect 5768 -1828 6940 -1800
rect 5768 -2652 6856 -1828
rect 6920 -2652 6940 -1828
rect 5768 -2680 6940 -2652
rect 7180 -1828 8352 -1800
rect 7180 -2652 8268 -1828
rect 8332 -2652 8352 -1828
rect 7180 -2680 8352 -2652
rect 8592 -1828 9764 -1800
rect 8592 -2652 9680 -1828
rect 9744 -2652 9764 -1828
rect 8592 -2680 9764 -2652
rect 10004 -1828 11176 -1800
rect 10004 -2652 11092 -1828
rect 11156 -2652 11176 -1828
rect 10004 -2680 11176 -2652
rect 11416 -1828 12588 -1800
rect 11416 -2652 12504 -1828
rect 12568 -2652 12588 -1828
rect 11416 -2680 12588 -2652
rect 12828 -1828 14000 -1800
rect 12828 -2652 13916 -1828
rect 13980 -2652 14000 -1828
rect 12828 -2680 14000 -2652
rect 14240 -1828 15412 -1800
rect 14240 -2652 15328 -1828
rect 15392 -2652 15412 -1828
rect 14240 -2680 15412 -2652
rect 15652 -1828 16824 -1800
rect 15652 -2652 16740 -1828
rect 16804 -2652 16824 -1828
rect 15652 -2680 16824 -2652
rect 17064 -1828 18236 -1800
rect 17064 -2652 18152 -1828
rect 18216 -2652 18236 -1828
rect 17064 -2680 18236 -2652
rect 18476 -1828 19648 -1800
rect 18476 -2652 19564 -1828
rect 19628 -2652 19648 -1828
rect 18476 -2680 19648 -2652
rect 19888 -1828 21060 -1800
rect 19888 -2652 20976 -1828
rect 21040 -2652 21060 -1828
rect 19888 -2680 21060 -2652
rect 21300 -1828 22472 -1800
rect 21300 -2652 22388 -1828
rect 22452 -2652 22472 -1828
rect 21300 -2680 22472 -2652
rect 22712 -1828 23884 -1800
rect 22712 -2652 23800 -1828
rect 23864 -2652 23884 -1828
rect 22712 -2680 23884 -2652
rect -23884 -2948 -22712 -2920
rect -23884 -3772 -22796 -2948
rect -22732 -3772 -22712 -2948
rect -23884 -3800 -22712 -3772
rect -22472 -2948 -21300 -2920
rect -22472 -3772 -21384 -2948
rect -21320 -3772 -21300 -2948
rect -22472 -3800 -21300 -3772
rect -21060 -2948 -19888 -2920
rect -21060 -3772 -19972 -2948
rect -19908 -3772 -19888 -2948
rect -21060 -3800 -19888 -3772
rect -19648 -2948 -18476 -2920
rect -19648 -3772 -18560 -2948
rect -18496 -3772 -18476 -2948
rect -19648 -3800 -18476 -3772
rect -18236 -2948 -17064 -2920
rect -18236 -3772 -17148 -2948
rect -17084 -3772 -17064 -2948
rect -18236 -3800 -17064 -3772
rect -16824 -2948 -15652 -2920
rect -16824 -3772 -15736 -2948
rect -15672 -3772 -15652 -2948
rect -16824 -3800 -15652 -3772
rect -15412 -2948 -14240 -2920
rect -15412 -3772 -14324 -2948
rect -14260 -3772 -14240 -2948
rect -15412 -3800 -14240 -3772
rect -14000 -2948 -12828 -2920
rect -14000 -3772 -12912 -2948
rect -12848 -3772 -12828 -2948
rect -14000 -3800 -12828 -3772
rect -12588 -2948 -11416 -2920
rect -12588 -3772 -11500 -2948
rect -11436 -3772 -11416 -2948
rect -12588 -3800 -11416 -3772
rect -11176 -2948 -10004 -2920
rect -11176 -3772 -10088 -2948
rect -10024 -3772 -10004 -2948
rect -11176 -3800 -10004 -3772
rect -9764 -2948 -8592 -2920
rect -9764 -3772 -8676 -2948
rect -8612 -3772 -8592 -2948
rect -9764 -3800 -8592 -3772
rect -8352 -2948 -7180 -2920
rect -8352 -3772 -7264 -2948
rect -7200 -3772 -7180 -2948
rect -8352 -3800 -7180 -3772
rect -6940 -2948 -5768 -2920
rect -6940 -3772 -5852 -2948
rect -5788 -3772 -5768 -2948
rect -6940 -3800 -5768 -3772
rect -5528 -2948 -4356 -2920
rect -5528 -3772 -4440 -2948
rect -4376 -3772 -4356 -2948
rect -5528 -3800 -4356 -3772
rect -4116 -2948 -2944 -2920
rect -4116 -3772 -3028 -2948
rect -2964 -3772 -2944 -2948
rect -4116 -3800 -2944 -3772
rect -2704 -2948 -1532 -2920
rect -2704 -3772 -1616 -2948
rect -1552 -3772 -1532 -2948
rect -2704 -3800 -1532 -3772
rect -1292 -2948 -120 -2920
rect -1292 -3772 -204 -2948
rect -140 -3772 -120 -2948
rect -1292 -3800 -120 -3772
rect 120 -2948 1292 -2920
rect 120 -3772 1208 -2948
rect 1272 -3772 1292 -2948
rect 120 -3800 1292 -3772
rect 1532 -2948 2704 -2920
rect 1532 -3772 2620 -2948
rect 2684 -3772 2704 -2948
rect 1532 -3800 2704 -3772
rect 2944 -2948 4116 -2920
rect 2944 -3772 4032 -2948
rect 4096 -3772 4116 -2948
rect 2944 -3800 4116 -3772
rect 4356 -2948 5528 -2920
rect 4356 -3772 5444 -2948
rect 5508 -3772 5528 -2948
rect 4356 -3800 5528 -3772
rect 5768 -2948 6940 -2920
rect 5768 -3772 6856 -2948
rect 6920 -3772 6940 -2948
rect 5768 -3800 6940 -3772
rect 7180 -2948 8352 -2920
rect 7180 -3772 8268 -2948
rect 8332 -3772 8352 -2948
rect 7180 -3800 8352 -3772
rect 8592 -2948 9764 -2920
rect 8592 -3772 9680 -2948
rect 9744 -3772 9764 -2948
rect 8592 -3800 9764 -3772
rect 10004 -2948 11176 -2920
rect 10004 -3772 11092 -2948
rect 11156 -3772 11176 -2948
rect 10004 -3800 11176 -3772
rect 11416 -2948 12588 -2920
rect 11416 -3772 12504 -2948
rect 12568 -3772 12588 -2948
rect 11416 -3800 12588 -3772
rect 12828 -2948 14000 -2920
rect 12828 -3772 13916 -2948
rect 13980 -3772 14000 -2948
rect 12828 -3800 14000 -3772
rect 14240 -2948 15412 -2920
rect 14240 -3772 15328 -2948
rect 15392 -3772 15412 -2948
rect 14240 -3800 15412 -3772
rect 15652 -2948 16824 -2920
rect 15652 -3772 16740 -2948
rect 16804 -3772 16824 -2948
rect 15652 -3800 16824 -3772
rect 17064 -2948 18236 -2920
rect 17064 -3772 18152 -2948
rect 18216 -3772 18236 -2948
rect 17064 -3800 18236 -3772
rect 18476 -2948 19648 -2920
rect 18476 -3772 19564 -2948
rect 19628 -3772 19648 -2948
rect 18476 -3800 19648 -3772
rect 19888 -2948 21060 -2920
rect 19888 -3772 20976 -2948
rect 21040 -3772 21060 -2948
rect 19888 -3800 21060 -3772
rect 21300 -2948 22472 -2920
rect 21300 -3772 22388 -2948
rect 22452 -3772 22472 -2948
rect 21300 -3800 22472 -3772
rect 22712 -2948 23884 -2920
rect 22712 -3772 23800 -2948
rect 23864 -3772 23884 -2948
rect 22712 -3800 23884 -3772
rect -23884 -4068 -22712 -4040
rect -23884 -4892 -22796 -4068
rect -22732 -4892 -22712 -4068
rect -23884 -4920 -22712 -4892
rect -22472 -4068 -21300 -4040
rect -22472 -4892 -21384 -4068
rect -21320 -4892 -21300 -4068
rect -22472 -4920 -21300 -4892
rect -21060 -4068 -19888 -4040
rect -21060 -4892 -19972 -4068
rect -19908 -4892 -19888 -4068
rect -21060 -4920 -19888 -4892
rect -19648 -4068 -18476 -4040
rect -19648 -4892 -18560 -4068
rect -18496 -4892 -18476 -4068
rect -19648 -4920 -18476 -4892
rect -18236 -4068 -17064 -4040
rect -18236 -4892 -17148 -4068
rect -17084 -4892 -17064 -4068
rect -18236 -4920 -17064 -4892
rect -16824 -4068 -15652 -4040
rect -16824 -4892 -15736 -4068
rect -15672 -4892 -15652 -4068
rect -16824 -4920 -15652 -4892
rect -15412 -4068 -14240 -4040
rect -15412 -4892 -14324 -4068
rect -14260 -4892 -14240 -4068
rect -15412 -4920 -14240 -4892
rect -14000 -4068 -12828 -4040
rect -14000 -4892 -12912 -4068
rect -12848 -4892 -12828 -4068
rect -14000 -4920 -12828 -4892
rect -12588 -4068 -11416 -4040
rect -12588 -4892 -11500 -4068
rect -11436 -4892 -11416 -4068
rect -12588 -4920 -11416 -4892
rect -11176 -4068 -10004 -4040
rect -11176 -4892 -10088 -4068
rect -10024 -4892 -10004 -4068
rect -11176 -4920 -10004 -4892
rect -9764 -4068 -8592 -4040
rect -9764 -4892 -8676 -4068
rect -8612 -4892 -8592 -4068
rect -9764 -4920 -8592 -4892
rect -8352 -4068 -7180 -4040
rect -8352 -4892 -7264 -4068
rect -7200 -4892 -7180 -4068
rect -8352 -4920 -7180 -4892
rect -6940 -4068 -5768 -4040
rect -6940 -4892 -5852 -4068
rect -5788 -4892 -5768 -4068
rect -6940 -4920 -5768 -4892
rect -5528 -4068 -4356 -4040
rect -5528 -4892 -4440 -4068
rect -4376 -4892 -4356 -4068
rect -5528 -4920 -4356 -4892
rect -4116 -4068 -2944 -4040
rect -4116 -4892 -3028 -4068
rect -2964 -4892 -2944 -4068
rect -4116 -4920 -2944 -4892
rect -2704 -4068 -1532 -4040
rect -2704 -4892 -1616 -4068
rect -1552 -4892 -1532 -4068
rect -2704 -4920 -1532 -4892
rect -1292 -4068 -120 -4040
rect -1292 -4892 -204 -4068
rect -140 -4892 -120 -4068
rect -1292 -4920 -120 -4892
rect 120 -4068 1292 -4040
rect 120 -4892 1208 -4068
rect 1272 -4892 1292 -4068
rect 120 -4920 1292 -4892
rect 1532 -4068 2704 -4040
rect 1532 -4892 2620 -4068
rect 2684 -4892 2704 -4068
rect 1532 -4920 2704 -4892
rect 2944 -4068 4116 -4040
rect 2944 -4892 4032 -4068
rect 4096 -4892 4116 -4068
rect 2944 -4920 4116 -4892
rect 4356 -4068 5528 -4040
rect 4356 -4892 5444 -4068
rect 5508 -4892 5528 -4068
rect 4356 -4920 5528 -4892
rect 5768 -4068 6940 -4040
rect 5768 -4892 6856 -4068
rect 6920 -4892 6940 -4068
rect 5768 -4920 6940 -4892
rect 7180 -4068 8352 -4040
rect 7180 -4892 8268 -4068
rect 8332 -4892 8352 -4068
rect 7180 -4920 8352 -4892
rect 8592 -4068 9764 -4040
rect 8592 -4892 9680 -4068
rect 9744 -4892 9764 -4068
rect 8592 -4920 9764 -4892
rect 10004 -4068 11176 -4040
rect 10004 -4892 11092 -4068
rect 11156 -4892 11176 -4068
rect 10004 -4920 11176 -4892
rect 11416 -4068 12588 -4040
rect 11416 -4892 12504 -4068
rect 12568 -4892 12588 -4068
rect 11416 -4920 12588 -4892
rect 12828 -4068 14000 -4040
rect 12828 -4892 13916 -4068
rect 13980 -4892 14000 -4068
rect 12828 -4920 14000 -4892
rect 14240 -4068 15412 -4040
rect 14240 -4892 15328 -4068
rect 15392 -4892 15412 -4068
rect 14240 -4920 15412 -4892
rect 15652 -4068 16824 -4040
rect 15652 -4892 16740 -4068
rect 16804 -4892 16824 -4068
rect 15652 -4920 16824 -4892
rect 17064 -4068 18236 -4040
rect 17064 -4892 18152 -4068
rect 18216 -4892 18236 -4068
rect 17064 -4920 18236 -4892
rect 18476 -4068 19648 -4040
rect 18476 -4892 19564 -4068
rect 19628 -4892 19648 -4068
rect 18476 -4920 19648 -4892
rect 19888 -4068 21060 -4040
rect 19888 -4892 20976 -4068
rect 21040 -4892 21060 -4068
rect 19888 -4920 21060 -4892
rect 21300 -4068 22472 -4040
rect 21300 -4892 22388 -4068
rect 22452 -4892 22472 -4068
rect 21300 -4920 22472 -4892
rect 22712 -4068 23884 -4040
rect 22712 -4892 23800 -4068
rect 23864 -4892 23884 -4068
rect 22712 -4920 23884 -4892
rect -23884 -5188 -22712 -5160
rect -23884 -6012 -22796 -5188
rect -22732 -6012 -22712 -5188
rect -23884 -6040 -22712 -6012
rect -22472 -5188 -21300 -5160
rect -22472 -6012 -21384 -5188
rect -21320 -6012 -21300 -5188
rect -22472 -6040 -21300 -6012
rect -21060 -5188 -19888 -5160
rect -21060 -6012 -19972 -5188
rect -19908 -6012 -19888 -5188
rect -21060 -6040 -19888 -6012
rect -19648 -5188 -18476 -5160
rect -19648 -6012 -18560 -5188
rect -18496 -6012 -18476 -5188
rect -19648 -6040 -18476 -6012
rect -18236 -5188 -17064 -5160
rect -18236 -6012 -17148 -5188
rect -17084 -6012 -17064 -5188
rect -18236 -6040 -17064 -6012
rect -16824 -5188 -15652 -5160
rect -16824 -6012 -15736 -5188
rect -15672 -6012 -15652 -5188
rect -16824 -6040 -15652 -6012
rect -15412 -5188 -14240 -5160
rect -15412 -6012 -14324 -5188
rect -14260 -6012 -14240 -5188
rect -15412 -6040 -14240 -6012
rect -14000 -5188 -12828 -5160
rect -14000 -6012 -12912 -5188
rect -12848 -6012 -12828 -5188
rect -14000 -6040 -12828 -6012
rect -12588 -5188 -11416 -5160
rect -12588 -6012 -11500 -5188
rect -11436 -6012 -11416 -5188
rect -12588 -6040 -11416 -6012
rect -11176 -5188 -10004 -5160
rect -11176 -6012 -10088 -5188
rect -10024 -6012 -10004 -5188
rect -11176 -6040 -10004 -6012
rect -9764 -5188 -8592 -5160
rect -9764 -6012 -8676 -5188
rect -8612 -6012 -8592 -5188
rect -9764 -6040 -8592 -6012
rect -8352 -5188 -7180 -5160
rect -8352 -6012 -7264 -5188
rect -7200 -6012 -7180 -5188
rect -8352 -6040 -7180 -6012
rect -6940 -5188 -5768 -5160
rect -6940 -6012 -5852 -5188
rect -5788 -6012 -5768 -5188
rect -6940 -6040 -5768 -6012
rect -5528 -5188 -4356 -5160
rect -5528 -6012 -4440 -5188
rect -4376 -6012 -4356 -5188
rect -5528 -6040 -4356 -6012
rect -4116 -5188 -2944 -5160
rect -4116 -6012 -3028 -5188
rect -2964 -6012 -2944 -5188
rect -4116 -6040 -2944 -6012
rect -2704 -5188 -1532 -5160
rect -2704 -6012 -1616 -5188
rect -1552 -6012 -1532 -5188
rect -2704 -6040 -1532 -6012
rect -1292 -5188 -120 -5160
rect -1292 -6012 -204 -5188
rect -140 -6012 -120 -5188
rect -1292 -6040 -120 -6012
rect 120 -5188 1292 -5160
rect 120 -6012 1208 -5188
rect 1272 -6012 1292 -5188
rect 120 -6040 1292 -6012
rect 1532 -5188 2704 -5160
rect 1532 -6012 2620 -5188
rect 2684 -6012 2704 -5188
rect 1532 -6040 2704 -6012
rect 2944 -5188 4116 -5160
rect 2944 -6012 4032 -5188
rect 4096 -6012 4116 -5188
rect 2944 -6040 4116 -6012
rect 4356 -5188 5528 -5160
rect 4356 -6012 5444 -5188
rect 5508 -6012 5528 -5188
rect 4356 -6040 5528 -6012
rect 5768 -5188 6940 -5160
rect 5768 -6012 6856 -5188
rect 6920 -6012 6940 -5188
rect 5768 -6040 6940 -6012
rect 7180 -5188 8352 -5160
rect 7180 -6012 8268 -5188
rect 8332 -6012 8352 -5188
rect 7180 -6040 8352 -6012
rect 8592 -5188 9764 -5160
rect 8592 -6012 9680 -5188
rect 9744 -6012 9764 -5188
rect 8592 -6040 9764 -6012
rect 10004 -5188 11176 -5160
rect 10004 -6012 11092 -5188
rect 11156 -6012 11176 -5188
rect 10004 -6040 11176 -6012
rect 11416 -5188 12588 -5160
rect 11416 -6012 12504 -5188
rect 12568 -6012 12588 -5188
rect 11416 -6040 12588 -6012
rect 12828 -5188 14000 -5160
rect 12828 -6012 13916 -5188
rect 13980 -6012 14000 -5188
rect 12828 -6040 14000 -6012
rect 14240 -5188 15412 -5160
rect 14240 -6012 15328 -5188
rect 15392 -6012 15412 -5188
rect 14240 -6040 15412 -6012
rect 15652 -5188 16824 -5160
rect 15652 -6012 16740 -5188
rect 16804 -6012 16824 -5188
rect 15652 -6040 16824 -6012
rect 17064 -5188 18236 -5160
rect 17064 -6012 18152 -5188
rect 18216 -6012 18236 -5188
rect 17064 -6040 18236 -6012
rect 18476 -5188 19648 -5160
rect 18476 -6012 19564 -5188
rect 19628 -6012 19648 -5188
rect 18476 -6040 19648 -6012
rect 19888 -5188 21060 -5160
rect 19888 -6012 20976 -5188
rect 21040 -6012 21060 -5188
rect 19888 -6040 21060 -6012
rect 21300 -5188 22472 -5160
rect 21300 -6012 22388 -5188
rect 22452 -6012 22472 -5188
rect 21300 -6040 22472 -6012
rect 22712 -5188 23884 -5160
rect 22712 -6012 23800 -5188
rect 23864 -6012 23884 -5188
rect 22712 -6040 23884 -6012
rect -23884 -6308 -22712 -6280
rect -23884 -7132 -22796 -6308
rect -22732 -7132 -22712 -6308
rect -23884 -7160 -22712 -7132
rect -22472 -6308 -21300 -6280
rect -22472 -7132 -21384 -6308
rect -21320 -7132 -21300 -6308
rect -22472 -7160 -21300 -7132
rect -21060 -6308 -19888 -6280
rect -21060 -7132 -19972 -6308
rect -19908 -7132 -19888 -6308
rect -21060 -7160 -19888 -7132
rect -19648 -6308 -18476 -6280
rect -19648 -7132 -18560 -6308
rect -18496 -7132 -18476 -6308
rect -19648 -7160 -18476 -7132
rect -18236 -6308 -17064 -6280
rect -18236 -7132 -17148 -6308
rect -17084 -7132 -17064 -6308
rect -18236 -7160 -17064 -7132
rect -16824 -6308 -15652 -6280
rect -16824 -7132 -15736 -6308
rect -15672 -7132 -15652 -6308
rect -16824 -7160 -15652 -7132
rect -15412 -6308 -14240 -6280
rect -15412 -7132 -14324 -6308
rect -14260 -7132 -14240 -6308
rect -15412 -7160 -14240 -7132
rect -14000 -6308 -12828 -6280
rect -14000 -7132 -12912 -6308
rect -12848 -7132 -12828 -6308
rect -14000 -7160 -12828 -7132
rect -12588 -6308 -11416 -6280
rect -12588 -7132 -11500 -6308
rect -11436 -7132 -11416 -6308
rect -12588 -7160 -11416 -7132
rect -11176 -6308 -10004 -6280
rect -11176 -7132 -10088 -6308
rect -10024 -7132 -10004 -6308
rect -11176 -7160 -10004 -7132
rect -9764 -6308 -8592 -6280
rect -9764 -7132 -8676 -6308
rect -8612 -7132 -8592 -6308
rect -9764 -7160 -8592 -7132
rect -8352 -6308 -7180 -6280
rect -8352 -7132 -7264 -6308
rect -7200 -7132 -7180 -6308
rect -8352 -7160 -7180 -7132
rect -6940 -6308 -5768 -6280
rect -6940 -7132 -5852 -6308
rect -5788 -7132 -5768 -6308
rect -6940 -7160 -5768 -7132
rect -5528 -6308 -4356 -6280
rect -5528 -7132 -4440 -6308
rect -4376 -7132 -4356 -6308
rect -5528 -7160 -4356 -7132
rect -4116 -6308 -2944 -6280
rect -4116 -7132 -3028 -6308
rect -2964 -7132 -2944 -6308
rect -4116 -7160 -2944 -7132
rect -2704 -6308 -1532 -6280
rect -2704 -7132 -1616 -6308
rect -1552 -7132 -1532 -6308
rect -2704 -7160 -1532 -7132
rect -1292 -6308 -120 -6280
rect -1292 -7132 -204 -6308
rect -140 -7132 -120 -6308
rect -1292 -7160 -120 -7132
rect 120 -6308 1292 -6280
rect 120 -7132 1208 -6308
rect 1272 -7132 1292 -6308
rect 120 -7160 1292 -7132
rect 1532 -6308 2704 -6280
rect 1532 -7132 2620 -6308
rect 2684 -7132 2704 -6308
rect 1532 -7160 2704 -7132
rect 2944 -6308 4116 -6280
rect 2944 -7132 4032 -6308
rect 4096 -7132 4116 -6308
rect 2944 -7160 4116 -7132
rect 4356 -6308 5528 -6280
rect 4356 -7132 5444 -6308
rect 5508 -7132 5528 -6308
rect 4356 -7160 5528 -7132
rect 5768 -6308 6940 -6280
rect 5768 -7132 6856 -6308
rect 6920 -7132 6940 -6308
rect 5768 -7160 6940 -7132
rect 7180 -6308 8352 -6280
rect 7180 -7132 8268 -6308
rect 8332 -7132 8352 -6308
rect 7180 -7160 8352 -7132
rect 8592 -6308 9764 -6280
rect 8592 -7132 9680 -6308
rect 9744 -7132 9764 -6308
rect 8592 -7160 9764 -7132
rect 10004 -6308 11176 -6280
rect 10004 -7132 11092 -6308
rect 11156 -7132 11176 -6308
rect 10004 -7160 11176 -7132
rect 11416 -6308 12588 -6280
rect 11416 -7132 12504 -6308
rect 12568 -7132 12588 -6308
rect 11416 -7160 12588 -7132
rect 12828 -6308 14000 -6280
rect 12828 -7132 13916 -6308
rect 13980 -7132 14000 -6308
rect 12828 -7160 14000 -7132
rect 14240 -6308 15412 -6280
rect 14240 -7132 15328 -6308
rect 15392 -7132 15412 -6308
rect 14240 -7160 15412 -7132
rect 15652 -6308 16824 -6280
rect 15652 -7132 16740 -6308
rect 16804 -7132 16824 -6308
rect 15652 -7160 16824 -7132
rect 17064 -6308 18236 -6280
rect 17064 -7132 18152 -6308
rect 18216 -7132 18236 -6308
rect 17064 -7160 18236 -7132
rect 18476 -6308 19648 -6280
rect 18476 -7132 19564 -6308
rect 19628 -7132 19648 -6308
rect 18476 -7160 19648 -7132
rect 19888 -6308 21060 -6280
rect 19888 -7132 20976 -6308
rect 21040 -7132 21060 -6308
rect 19888 -7160 21060 -7132
rect 21300 -6308 22472 -6280
rect 21300 -7132 22388 -6308
rect 22452 -7132 22472 -6308
rect 21300 -7160 22472 -7132
rect 22712 -6308 23884 -6280
rect 22712 -7132 23800 -6308
rect 23864 -7132 23884 -6308
rect 22712 -7160 23884 -7132
rect -23884 -7428 -22712 -7400
rect -23884 -8252 -22796 -7428
rect -22732 -8252 -22712 -7428
rect -23884 -8280 -22712 -8252
rect -22472 -7428 -21300 -7400
rect -22472 -8252 -21384 -7428
rect -21320 -8252 -21300 -7428
rect -22472 -8280 -21300 -8252
rect -21060 -7428 -19888 -7400
rect -21060 -8252 -19972 -7428
rect -19908 -8252 -19888 -7428
rect -21060 -8280 -19888 -8252
rect -19648 -7428 -18476 -7400
rect -19648 -8252 -18560 -7428
rect -18496 -8252 -18476 -7428
rect -19648 -8280 -18476 -8252
rect -18236 -7428 -17064 -7400
rect -18236 -8252 -17148 -7428
rect -17084 -8252 -17064 -7428
rect -18236 -8280 -17064 -8252
rect -16824 -7428 -15652 -7400
rect -16824 -8252 -15736 -7428
rect -15672 -8252 -15652 -7428
rect -16824 -8280 -15652 -8252
rect -15412 -7428 -14240 -7400
rect -15412 -8252 -14324 -7428
rect -14260 -8252 -14240 -7428
rect -15412 -8280 -14240 -8252
rect -14000 -7428 -12828 -7400
rect -14000 -8252 -12912 -7428
rect -12848 -8252 -12828 -7428
rect -14000 -8280 -12828 -8252
rect -12588 -7428 -11416 -7400
rect -12588 -8252 -11500 -7428
rect -11436 -8252 -11416 -7428
rect -12588 -8280 -11416 -8252
rect -11176 -7428 -10004 -7400
rect -11176 -8252 -10088 -7428
rect -10024 -8252 -10004 -7428
rect -11176 -8280 -10004 -8252
rect -9764 -7428 -8592 -7400
rect -9764 -8252 -8676 -7428
rect -8612 -8252 -8592 -7428
rect -9764 -8280 -8592 -8252
rect -8352 -7428 -7180 -7400
rect -8352 -8252 -7264 -7428
rect -7200 -8252 -7180 -7428
rect -8352 -8280 -7180 -8252
rect -6940 -7428 -5768 -7400
rect -6940 -8252 -5852 -7428
rect -5788 -8252 -5768 -7428
rect -6940 -8280 -5768 -8252
rect -5528 -7428 -4356 -7400
rect -5528 -8252 -4440 -7428
rect -4376 -8252 -4356 -7428
rect -5528 -8280 -4356 -8252
rect -4116 -7428 -2944 -7400
rect -4116 -8252 -3028 -7428
rect -2964 -8252 -2944 -7428
rect -4116 -8280 -2944 -8252
rect -2704 -7428 -1532 -7400
rect -2704 -8252 -1616 -7428
rect -1552 -8252 -1532 -7428
rect -2704 -8280 -1532 -8252
rect -1292 -7428 -120 -7400
rect -1292 -8252 -204 -7428
rect -140 -8252 -120 -7428
rect -1292 -8280 -120 -8252
rect 120 -7428 1292 -7400
rect 120 -8252 1208 -7428
rect 1272 -8252 1292 -7428
rect 120 -8280 1292 -8252
rect 1532 -7428 2704 -7400
rect 1532 -8252 2620 -7428
rect 2684 -8252 2704 -7428
rect 1532 -8280 2704 -8252
rect 2944 -7428 4116 -7400
rect 2944 -8252 4032 -7428
rect 4096 -8252 4116 -7428
rect 2944 -8280 4116 -8252
rect 4356 -7428 5528 -7400
rect 4356 -8252 5444 -7428
rect 5508 -8252 5528 -7428
rect 4356 -8280 5528 -8252
rect 5768 -7428 6940 -7400
rect 5768 -8252 6856 -7428
rect 6920 -8252 6940 -7428
rect 5768 -8280 6940 -8252
rect 7180 -7428 8352 -7400
rect 7180 -8252 8268 -7428
rect 8332 -8252 8352 -7428
rect 7180 -8280 8352 -8252
rect 8592 -7428 9764 -7400
rect 8592 -8252 9680 -7428
rect 9744 -8252 9764 -7428
rect 8592 -8280 9764 -8252
rect 10004 -7428 11176 -7400
rect 10004 -8252 11092 -7428
rect 11156 -8252 11176 -7428
rect 10004 -8280 11176 -8252
rect 11416 -7428 12588 -7400
rect 11416 -8252 12504 -7428
rect 12568 -8252 12588 -7428
rect 11416 -8280 12588 -8252
rect 12828 -7428 14000 -7400
rect 12828 -8252 13916 -7428
rect 13980 -8252 14000 -7428
rect 12828 -8280 14000 -8252
rect 14240 -7428 15412 -7400
rect 14240 -8252 15328 -7428
rect 15392 -8252 15412 -7428
rect 14240 -8280 15412 -8252
rect 15652 -7428 16824 -7400
rect 15652 -8252 16740 -7428
rect 16804 -8252 16824 -7428
rect 15652 -8280 16824 -8252
rect 17064 -7428 18236 -7400
rect 17064 -8252 18152 -7428
rect 18216 -8252 18236 -7428
rect 17064 -8280 18236 -8252
rect 18476 -7428 19648 -7400
rect 18476 -8252 19564 -7428
rect 19628 -8252 19648 -7428
rect 18476 -8280 19648 -8252
rect 19888 -7428 21060 -7400
rect 19888 -8252 20976 -7428
rect 21040 -8252 21060 -7428
rect 19888 -8280 21060 -8252
rect 21300 -7428 22472 -7400
rect 21300 -8252 22388 -7428
rect 22452 -8252 22472 -7428
rect 21300 -8280 22472 -8252
rect 22712 -7428 23884 -7400
rect 22712 -8252 23800 -7428
rect 23864 -8252 23884 -7428
rect 22712 -8280 23884 -8252
rect -23884 -8548 -22712 -8520
rect -23884 -9372 -22796 -8548
rect -22732 -9372 -22712 -8548
rect -23884 -9400 -22712 -9372
rect -22472 -8548 -21300 -8520
rect -22472 -9372 -21384 -8548
rect -21320 -9372 -21300 -8548
rect -22472 -9400 -21300 -9372
rect -21060 -8548 -19888 -8520
rect -21060 -9372 -19972 -8548
rect -19908 -9372 -19888 -8548
rect -21060 -9400 -19888 -9372
rect -19648 -8548 -18476 -8520
rect -19648 -9372 -18560 -8548
rect -18496 -9372 -18476 -8548
rect -19648 -9400 -18476 -9372
rect -18236 -8548 -17064 -8520
rect -18236 -9372 -17148 -8548
rect -17084 -9372 -17064 -8548
rect -18236 -9400 -17064 -9372
rect -16824 -8548 -15652 -8520
rect -16824 -9372 -15736 -8548
rect -15672 -9372 -15652 -8548
rect -16824 -9400 -15652 -9372
rect -15412 -8548 -14240 -8520
rect -15412 -9372 -14324 -8548
rect -14260 -9372 -14240 -8548
rect -15412 -9400 -14240 -9372
rect -14000 -8548 -12828 -8520
rect -14000 -9372 -12912 -8548
rect -12848 -9372 -12828 -8548
rect -14000 -9400 -12828 -9372
rect -12588 -8548 -11416 -8520
rect -12588 -9372 -11500 -8548
rect -11436 -9372 -11416 -8548
rect -12588 -9400 -11416 -9372
rect -11176 -8548 -10004 -8520
rect -11176 -9372 -10088 -8548
rect -10024 -9372 -10004 -8548
rect -11176 -9400 -10004 -9372
rect -9764 -8548 -8592 -8520
rect -9764 -9372 -8676 -8548
rect -8612 -9372 -8592 -8548
rect -9764 -9400 -8592 -9372
rect -8352 -8548 -7180 -8520
rect -8352 -9372 -7264 -8548
rect -7200 -9372 -7180 -8548
rect -8352 -9400 -7180 -9372
rect -6940 -8548 -5768 -8520
rect -6940 -9372 -5852 -8548
rect -5788 -9372 -5768 -8548
rect -6940 -9400 -5768 -9372
rect -5528 -8548 -4356 -8520
rect -5528 -9372 -4440 -8548
rect -4376 -9372 -4356 -8548
rect -5528 -9400 -4356 -9372
rect -4116 -8548 -2944 -8520
rect -4116 -9372 -3028 -8548
rect -2964 -9372 -2944 -8548
rect -4116 -9400 -2944 -9372
rect -2704 -8548 -1532 -8520
rect -2704 -9372 -1616 -8548
rect -1552 -9372 -1532 -8548
rect -2704 -9400 -1532 -9372
rect -1292 -8548 -120 -8520
rect -1292 -9372 -204 -8548
rect -140 -9372 -120 -8548
rect -1292 -9400 -120 -9372
rect 120 -8548 1292 -8520
rect 120 -9372 1208 -8548
rect 1272 -9372 1292 -8548
rect 120 -9400 1292 -9372
rect 1532 -8548 2704 -8520
rect 1532 -9372 2620 -8548
rect 2684 -9372 2704 -8548
rect 1532 -9400 2704 -9372
rect 2944 -8548 4116 -8520
rect 2944 -9372 4032 -8548
rect 4096 -9372 4116 -8548
rect 2944 -9400 4116 -9372
rect 4356 -8548 5528 -8520
rect 4356 -9372 5444 -8548
rect 5508 -9372 5528 -8548
rect 4356 -9400 5528 -9372
rect 5768 -8548 6940 -8520
rect 5768 -9372 6856 -8548
rect 6920 -9372 6940 -8548
rect 5768 -9400 6940 -9372
rect 7180 -8548 8352 -8520
rect 7180 -9372 8268 -8548
rect 8332 -9372 8352 -8548
rect 7180 -9400 8352 -9372
rect 8592 -8548 9764 -8520
rect 8592 -9372 9680 -8548
rect 9744 -9372 9764 -8548
rect 8592 -9400 9764 -9372
rect 10004 -8548 11176 -8520
rect 10004 -9372 11092 -8548
rect 11156 -9372 11176 -8548
rect 10004 -9400 11176 -9372
rect 11416 -8548 12588 -8520
rect 11416 -9372 12504 -8548
rect 12568 -9372 12588 -8548
rect 11416 -9400 12588 -9372
rect 12828 -8548 14000 -8520
rect 12828 -9372 13916 -8548
rect 13980 -9372 14000 -8548
rect 12828 -9400 14000 -9372
rect 14240 -8548 15412 -8520
rect 14240 -9372 15328 -8548
rect 15392 -9372 15412 -8548
rect 14240 -9400 15412 -9372
rect 15652 -8548 16824 -8520
rect 15652 -9372 16740 -8548
rect 16804 -9372 16824 -8548
rect 15652 -9400 16824 -9372
rect 17064 -8548 18236 -8520
rect 17064 -9372 18152 -8548
rect 18216 -9372 18236 -8548
rect 17064 -9400 18236 -9372
rect 18476 -8548 19648 -8520
rect 18476 -9372 19564 -8548
rect 19628 -9372 19648 -8548
rect 18476 -9400 19648 -9372
rect 19888 -8548 21060 -8520
rect 19888 -9372 20976 -8548
rect 21040 -9372 21060 -8548
rect 19888 -9400 21060 -9372
rect 21300 -8548 22472 -8520
rect 21300 -9372 22388 -8548
rect 22452 -9372 22472 -8548
rect 21300 -9400 22472 -9372
rect 22712 -8548 23884 -8520
rect 22712 -9372 23800 -8548
rect 23864 -9372 23884 -8548
rect 22712 -9400 23884 -9372
rect -23884 -9668 -22712 -9640
rect -23884 -10492 -22796 -9668
rect -22732 -10492 -22712 -9668
rect -23884 -10520 -22712 -10492
rect -22472 -9668 -21300 -9640
rect -22472 -10492 -21384 -9668
rect -21320 -10492 -21300 -9668
rect -22472 -10520 -21300 -10492
rect -21060 -9668 -19888 -9640
rect -21060 -10492 -19972 -9668
rect -19908 -10492 -19888 -9668
rect -21060 -10520 -19888 -10492
rect -19648 -9668 -18476 -9640
rect -19648 -10492 -18560 -9668
rect -18496 -10492 -18476 -9668
rect -19648 -10520 -18476 -10492
rect -18236 -9668 -17064 -9640
rect -18236 -10492 -17148 -9668
rect -17084 -10492 -17064 -9668
rect -18236 -10520 -17064 -10492
rect -16824 -9668 -15652 -9640
rect -16824 -10492 -15736 -9668
rect -15672 -10492 -15652 -9668
rect -16824 -10520 -15652 -10492
rect -15412 -9668 -14240 -9640
rect -15412 -10492 -14324 -9668
rect -14260 -10492 -14240 -9668
rect -15412 -10520 -14240 -10492
rect -14000 -9668 -12828 -9640
rect -14000 -10492 -12912 -9668
rect -12848 -10492 -12828 -9668
rect -14000 -10520 -12828 -10492
rect -12588 -9668 -11416 -9640
rect -12588 -10492 -11500 -9668
rect -11436 -10492 -11416 -9668
rect -12588 -10520 -11416 -10492
rect -11176 -9668 -10004 -9640
rect -11176 -10492 -10088 -9668
rect -10024 -10492 -10004 -9668
rect -11176 -10520 -10004 -10492
rect -9764 -9668 -8592 -9640
rect -9764 -10492 -8676 -9668
rect -8612 -10492 -8592 -9668
rect -9764 -10520 -8592 -10492
rect -8352 -9668 -7180 -9640
rect -8352 -10492 -7264 -9668
rect -7200 -10492 -7180 -9668
rect -8352 -10520 -7180 -10492
rect -6940 -9668 -5768 -9640
rect -6940 -10492 -5852 -9668
rect -5788 -10492 -5768 -9668
rect -6940 -10520 -5768 -10492
rect -5528 -9668 -4356 -9640
rect -5528 -10492 -4440 -9668
rect -4376 -10492 -4356 -9668
rect -5528 -10520 -4356 -10492
rect -4116 -9668 -2944 -9640
rect -4116 -10492 -3028 -9668
rect -2964 -10492 -2944 -9668
rect -4116 -10520 -2944 -10492
rect -2704 -9668 -1532 -9640
rect -2704 -10492 -1616 -9668
rect -1552 -10492 -1532 -9668
rect -2704 -10520 -1532 -10492
rect -1292 -9668 -120 -9640
rect -1292 -10492 -204 -9668
rect -140 -10492 -120 -9668
rect -1292 -10520 -120 -10492
rect 120 -9668 1292 -9640
rect 120 -10492 1208 -9668
rect 1272 -10492 1292 -9668
rect 120 -10520 1292 -10492
rect 1532 -9668 2704 -9640
rect 1532 -10492 2620 -9668
rect 2684 -10492 2704 -9668
rect 1532 -10520 2704 -10492
rect 2944 -9668 4116 -9640
rect 2944 -10492 4032 -9668
rect 4096 -10492 4116 -9668
rect 2944 -10520 4116 -10492
rect 4356 -9668 5528 -9640
rect 4356 -10492 5444 -9668
rect 5508 -10492 5528 -9668
rect 4356 -10520 5528 -10492
rect 5768 -9668 6940 -9640
rect 5768 -10492 6856 -9668
rect 6920 -10492 6940 -9668
rect 5768 -10520 6940 -10492
rect 7180 -9668 8352 -9640
rect 7180 -10492 8268 -9668
rect 8332 -10492 8352 -9668
rect 7180 -10520 8352 -10492
rect 8592 -9668 9764 -9640
rect 8592 -10492 9680 -9668
rect 9744 -10492 9764 -9668
rect 8592 -10520 9764 -10492
rect 10004 -9668 11176 -9640
rect 10004 -10492 11092 -9668
rect 11156 -10492 11176 -9668
rect 10004 -10520 11176 -10492
rect 11416 -9668 12588 -9640
rect 11416 -10492 12504 -9668
rect 12568 -10492 12588 -9668
rect 11416 -10520 12588 -10492
rect 12828 -9668 14000 -9640
rect 12828 -10492 13916 -9668
rect 13980 -10492 14000 -9668
rect 12828 -10520 14000 -10492
rect 14240 -9668 15412 -9640
rect 14240 -10492 15328 -9668
rect 15392 -10492 15412 -9668
rect 14240 -10520 15412 -10492
rect 15652 -9668 16824 -9640
rect 15652 -10492 16740 -9668
rect 16804 -10492 16824 -9668
rect 15652 -10520 16824 -10492
rect 17064 -9668 18236 -9640
rect 17064 -10492 18152 -9668
rect 18216 -10492 18236 -9668
rect 17064 -10520 18236 -10492
rect 18476 -9668 19648 -9640
rect 18476 -10492 19564 -9668
rect 19628 -10492 19648 -9668
rect 18476 -10520 19648 -10492
rect 19888 -9668 21060 -9640
rect 19888 -10492 20976 -9668
rect 21040 -10492 21060 -9668
rect 19888 -10520 21060 -10492
rect 21300 -9668 22472 -9640
rect 21300 -10492 22388 -9668
rect 22452 -10492 22472 -9668
rect 21300 -10520 22472 -10492
rect 22712 -9668 23884 -9640
rect 22712 -10492 23800 -9668
rect 23864 -10492 23884 -9668
rect 22712 -10520 23884 -10492
rect -23884 -10788 -22712 -10760
rect -23884 -11612 -22796 -10788
rect -22732 -11612 -22712 -10788
rect -23884 -11640 -22712 -11612
rect -22472 -10788 -21300 -10760
rect -22472 -11612 -21384 -10788
rect -21320 -11612 -21300 -10788
rect -22472 -11640 -21300 -11612
rect -21060 -10788 -19888 -10760
rect -21060 -11612 -19972 -10788
rect -19908 -11612 -19888 -10788
rect -21060 -11640 -19888 -11612
rect -19648 -10788 -18476 -10760
rect -19648 -11612 -18560 -10788
rect -18496 -11612 -18476 -10788
rect -19648 -11640 -18476 -11612
rect -18236 -10788 -17064 -10760
rect -18236 -11612 -17148 -10788
rect -17084 -11612 -17064 -10788
rect -18236 -11640 -17064 -11612
rect -16824 -10788 -15652 -10760
rect -16824 -11612 -15736 -10788
rect -15672 -11612 -15652 -10788
rect -16824 -11640 -15652 -11612
rect -15412 -10788 -14240 -10760
rect -15412 -11612 -14324 -10788
rect -14260 -11612 -14240 -10788
rect -15412 -11640 -14240 -11612
rect -14000 -10788 -12828 -10760
rect -14000 -11612 -12912 -10788
rect -12848 -11612 -12828 -10788
rect -14000 -11640 -12828 -11612
rect -12588 -10788 -11416 -10760
rect -12588 -11612 -11500 -10788
rect -11436 -11612 -11416 -10788
rect -12588 -11640 -11416 -11612
rect -11176 -10788 -10004 -10760
rect -11176 -11612 -10088 -10788
rect -10024 -11612 -10004 -10788
rect -11176 -11640 -10004 -11612
rect -9764 -10788 -8592 -10760
rect -9764 -11612 -8676 -10788
rect -8612 -11612 -8592 -10788
rect -9764 -11640 -8592 -11612
rect -8352 -10788 -7180 -10760
rect -8352 -11612 -7264 -10788
rect -7200 -11612 -7180 -10788
rect -8352 -11640 -7180 -11612
rect -6940 -10788 -5768 -10760
rect -6940 -11612 -5852 -10788
rect -5788 -11612 -5768 -10788
rect -6940 -11640 -5768 -11612
rect -5528 -10788 -4356 -10760
rect -5528 -11612 -4440 -10788
rect -4376 -11612 -4356 -10788
rect -5528 -11640 -4356 -11612
rect -4116 -10788 -2944 -10760
rect -4116 -11612 -3028 -10788
rect -2964 -11612 -2944 -10788
rect -4116 -11640 -2944 -11612
rect -2704 -10788 -1532 -10760
rect -2704 -11612 -1616 -10788
rect -1552 -11612 -1532 -10788
rect -2704 -11640 -1532 -11612
rect -1292 -10788 -120 -10760
rect -1292 -11612 -204 -10788
rect -140 -11612 -120 -10788
rect -1292 -11640 -120 -11612
rect 120 -10788 1292 -10760
rect 120 -11612 1208 -10788
rect 1272 -11612 1292 -10788
rect 120 -11640 1292 -11612
rect 1532 -10788 2704 -10760
rect 1532 -11612 2620 -10788
rect 2684 -11612 2704 -10788
rect 1532 -11640 2704 -11612
rect 2944 -10788 4116 -10760
rect 2944 -11612 4032 -10788
rect 4096 -11612 4116 -10788
rect 2944 -11640 4116 -11612
rect 4356 -10788 5528 -10760
rect 4356 -11612 5444 -10788
rect 5508 -11612 5528 -10788
rect 4356 -11640 5528 -11612
rect 5768 -10788 6940 -10760
rect 5768 -11612 6856 -10788
rect 6920 -11612 6940 -10788
rect 5768 -11640 6940 -11612
rect 7180 -10788 8352 -10760
rect 7180 -11612 8268 -10788
rect 8332 -11612 8352 -10788
rect 7180 -11640 8352 -11612
rect 8592 -10788 9764 -10760
rect 8592 -11612 9680 -10788
rect 9744 -11612 9764 -10788
rect 8592 -11640 9764 -11612
rect 10004 -10788 11176 -10760
rect 10004 -11612 11092 -10788
rect 11156 -11612 11176 -10788
rect 10004 -11640 11176 -11612
rect 11416 -10788 12588 -10760
rect 11416 -11612 12504 -10788
rect 12568 -11612 12588 -10788
rect 11416 -11640 12588 -11612
rect 12828 -10788 14000 -10760
rect 12828 -11612 13916 -10788
rect 13980 -11612 14000 -10788
rect 12828 -11640 14000 -11612
rect 14240 -10788 15412 -10760
rect 14240 -11612 15328 -10788
rect 15392 -11612 15412 -10788
rect 14240 -11640 15412 -11612
rect 15652 -10788 16824 -10760
rect 15652 -11612 16740 -10788
rect 16804 -11612 16824 -10788
rect 15652 -11640 16824 -11612
rect 17064 -10788 18236 -10760
rect 17064 -11612 18152 -10788
rect 18216 -11612 18236 -10788
rect 17064 -11640 18236 -11612
rect 18476 -10788 19648 -10760
rect 18476 -11612 19564 -10788
rect 19628 -11612 19648 -10788
rect 18476 -11640 19648 -11612
rect 19888 -10788 21060 -10760
rect 19888 -11612 20976 -10788
rect 21040 -11612 21060 -10788
rect 19888 -11640 21060 -11612
rect 21300 -10788 22472 -10760
rect 21300 -11612 22388 -10788
rect 22452 -11612 22472 -10788
rect 21300 -11640 22472 -11612
rect 22712 -10788 23884 -10760
rect 22712 -11612 23800 -10788
rect 23864 -11612 23884 -10788
rect 22712 -11640 23884 -11612
rect -23884 -11908 -22712 -11880
rect -23884 -12732 -22796 -11908
rect -22732 -12732 -22712 -11908
rect -23884 -12760 -22712 -12732
rect -22472 -11908 -21300 -11880
rect -22472 -12732 -21384 -11908
rect -21320 -12732 -21300 -11908
rect -22472 -12760 -21300 -12732
rect -21060 -11908 -19888 -11880
rect -21060 -12732 -19972 -11908
rect -19908 -12732 -19888 -11908
rect -21060 -12760 -19888 -12732
rect -19648 -11908 -18476 -11880
rect -19648 -12732 -18560 -11908
rect -18496 -12732 -18476 -11908
rect -19648 -12760 -18476 -12732
rect -18236 -11908 -17064 -11880
rect -18236 -12732 -17148 -11908
rect -17084 -12732 -17064 -11908
rect -18236 -12760 -17064 -12732
rect -16824 -11908 -15652 -11880
rect -16824 -12732 -15736 -11908
rect -15672 -12732 -15652 -11908
rect -16824 -12760 -15652 -12732
rect -15412 -11908 -14240 -11880
rect -15412 -12732 -14324 -11908
rect -14260 -12732 -14240 -11908
rect -15412 -12760 -14240 -12732
rect -14000 -11908 -12828 -11880
rect -14000 -12732 -12912 -11908
rect -12848 -12732 -12828 -11908
rect -14000 -12760 -12828 -12732
rect -12588 -11908 -11416 -11880
rect -12588 -12732 -11500 -11908
rect -11436 -12732 -11416 -11908
rect -12588 -12760 -11416 -12732
rect -11176 -11908 -10004 -11880
rect -11176 -12732 -10088 -11908
rect -10024 -12732 -10004 -11908
rect -11176 -12760 -10004 -12732
rect -9764 -11908 -8592 -11880
rect -9764 -12732 -8676 -11908
rect -8612 -12732 -8592 -11908
rect -9764 -12760 -8592 -12732
rect -8352 -11908 -7180 -11880
rect -8352 -12732 -7264 -11908
rect -7200 -12732 -7180 -11908
rect -8352 -12760 -7180 -12732
rect -6940 -11908 -5768 -11880
rect -6940 -12732 -5852 -11908
rect -5788 -12732 -5768 -11908
rect -6940 -12760 -5768 -12732
rect -5528 -11908 -4356 -11880
rect -5528 -12732 -4440 -11908
rect -4376 -12732 -4356 -11908
rect -5528 -12760 -4356 -12732
rect -4116 -11908 -2944 -11880
rect -4116 -12732 -3028 -11908
rect -2964 -12732 -2944 -11908
rect -4116 -12760 -2944 -12732
rect -2704 -11908 -1532 -11880
rect -2704 -12732 -1616 -11908
rect -1552 -12732 -1532 -11908
rect -2704 -12760 -1532 -12732
rect -1292 -11908 -120 -11880
rect -1292 -12732 -204 -11908
rect -140 -12732 -120 -11908
rect -1292 -12760 -120 -12732
rect 120 -11908 1292 -11880
rect 120 -12732 1208 -11908
rect 1272 -12732 1292 -11908
rect 120 -12760 1292 -12732
rect 1532 -11908 2704 -11880
rect 1532 -12732 2620 -11908
rect 2684 -12732 2704 -11908
rect 1532 -12760 2704 -12732
rect 2944 -11908 4116 -11880
rect 2944 -12732 4032 -11908
rect 4096 -12732 4116 -11908
rect 2944 -12760 4116 -12732
rect 4356 -11908 5528 -11880
rect 4356 -12732 5444 -11908
rect 5508 -12732 5528 -11908
rect 4356 -12760 5528 -12732
rect 5768 -11908 6940 -11880
rect 5768 -12732 6856 -11908
rect 6920 -12732 6940 -11908
rect 5768 -12760 6940 -12732
rect 7180 -11908 8352 -11880
rect 7180 -12732 8268 -11908
rect 8332 -12732 8352 -11908
rect 7180 -12760 8352 -12732
rect 8592 -11908 9764 -11880
rect 8592 -12732 9680 -11908
rect 9744 -12732 9764 -11908
rect 8592 -12760 9764 -12732
rect 10004 -11908 11176 -11880
rect 10004 -12732 11092 -11908
rect 11156 -12732 11176 -11908
rect 10004 -12760 11176 -12732
rect 11416 -11908 12588 -11880
rect 11416 -12732 12504 -11908
rect 12568 -12732 12588 -11908
rect 11416 -12760 12588 -12732
rect 12828 -11908 14000 -11880
rect 12828 -12732 13916 -11908
rect 13980 -12732 14000 -11908
rect 12828 -12760 14000 -12732
rect 14240 -11908 15412 -11880
rect 14240 -12732 15328 -11908
rect 15392 -12732 15412 -11908
rect 14240 -12760 15412 -12732
rect 15652 -11908 16824 -11880
rect 15652 -12732 16740 -11908
rect 16804 -12732 16824 -11908
rect 15652 -12760 16824 -12732
rect 17064 -11908 18236 -11880
rect 17064 -12732 18152 -11908
rect 18216 -12732 18236 -11908
rect 17064 -12760 18236 -12732
rect 18476 -11908 19648 -11880
rect 18476 -12732 19564 -11908
rect 19628 -12732 19648 -11908
rect 18476 -12760 19648 -12732
rect 19888 -11908 21060 -11880
rect 19888 -12732 20976 -11908
rect 21040 -12732 21060 -11908
rect 19888 -12760 21060 -12732
rect 21300 -11908 22472 -11880
rect 21300 -12732 22388 -11908
rect 22452 -12732 22472 -11908
rect 21300 -12760 22472 -12732
rect 22712 -11908 23884 -11880
rect 22712 -12732 23800 -11908
rect 23864 -12732 23884 -11908
rect 22712 -12760 23884 -12732
rect -23884 -13028 -22712 -13000
rect -23884 -13852 -22796 -13028
rect -22732 -13852 -22712 -13028
rect -23884 -13880 -22712 -13852
rect -22472 -13028 -21300 -13000
rect -22472 -13852 -21384 -13028
rect -21320 -13852 -21300 -13028
rect -22472 -13880 -21300 -13852
rect -21060 -13028 -19888 -13000
rect -21060 -13852 -19972 -13028
rect -19908 -13852 -19888 -13028
rect -21060 -13880 -19888 -13852
rect -19648 -13028 -18476 -13000
rect -19648 -13852 -18560 -13028
rect -18496 -13852 -18476 -13028
rect -19648 -13880 -18476 -13852
rect -18236 -13028 -17064 -13000
rect -18236 -13852 -17148 -13028
rect -17084 -13852 -17064 -13028
rect -18236 -13880 -17064 -13852
rect -16824 -13028 -15652 -13000
rect -16824 -13852 -15736 -13028
rect -15672 -13852 -15652 -13028
rect -16824 -13880 -15652 -13852
rect -15412 -13028 -14240 -13000
rect -15412 -13852 -14324 -13028
rect -14260 -13852 -14240 -13028
rect -15412 -13880 -14240 -13852
rect -14000 -13028 -12828 -13000
rect -14000 -13852 -12912 -13028
rect -12848 -13852 -12828 -13028
rect -14000 -13880 -12828 -13852
rect -12588 -13028 -11416 -13000
rect -12588 -13852 -11500 -13028
rect -11436 -13852 -11416 -13028
rect -12588 -13880 -11416 -13852
rect -11176 -13028 -10004 -13000
rect -11176 -13852 -10088 -13028
rect -10024 -13852 -10004 -13028
rect -11176 -13880 -10004 -13852
rect -9764 -13028 -8592 -13000
rect -9764 -13852 -8676 -13028
rect -8612 -13852 -8592 -13028
rect -9764 -13880 -8592 -13852
rect -8352 -13028 -7180 -13000
rect -8352 -13852 -7264 -13028
rect -7200 -13852 -7180 -13028
rect -8352 -13880 -7180 -13852
rect -6940 -13028 -5768 -13000
rect -6940 -13852 -5852 -13028
rect -5788 -13852 -5768 -13028
rect -6940 -13880 -5768 -13852
rect -5528 -13028 -4356 -13000
rect -5528 -13852 -4440 -13028
rect -4376 -13852 -4356 -13028
rect -5528 -13880 -4356 -13852
rect -4116 -13028 -2944 -13000
rect -4116 -13852 -3028 -13028
rect -2964 -13852 -2944 -13028
rect -4116 -13880 -2944 -13852
rect -2704 -13028 -1532 -13000
rect -2704 -13852 -1616 -13028
rect -1552 -13852 -1532 -13028
rect -2704 -13880 -1532 -13852
rect -1292 -13028 -120 -13000
rect -1292 -13852 -204 -13028
rect -140 -13852 -120 -13028
rect -1292 -13880 -120 -13852
rect 120 -13028 1292 -13000
rect 120 -13852 1208 -13028
rect 1272 -13852 1292 -13028
rect 120 -13880 1292 -13852
rect 1532 -13028 2704 -13000
rect 1532 -13852 2620 -13028
rect 2684 -13852 2704 -13028
rect 1532 -13880 2704 -13852
rect 2944 -13028 4116 -13000
rect 2944 -13852 4032 -13028
rect 4096 -13852 4116 -13028
rect 2944 -13880 4116 -13852
rect 4356 -13028 5528 -13000
rect 4356 -13852 5444 -13028
rect 5508 -13852 5528 -13028
rect 4356 -13880 5528 -13852
rect 5768 -13028 6940 -13000
rect 5768 -13852 6856 -13028
rect 6920 -13852 6940 -13028
rect 5768 -13880 6940 -13852
rect 7180 -13028 8352 -13000
rect 7180 -13852 8268 -13028
rect 8332 -13852 8352 -13028
rect 7180 -13880 8352 -13852
rect 8592 -13028 9764 -13000
rect 8592 -13852 9680 -13028
rect 9744 -13852 9764 -13028
rect 8592 -13880 9764 -13852
rect 10004 -13028 11176 -13000
rect 10004 -13852 11092 -13028
rect 11156 -13852 11176 -13028
rect 10004 -13880 11176 -13852
rect 11416 -13028 12588 -13000
rect 11416 -13852 12504 -13028
rect 12568 -13852 12588 -13028
rect 11416 -13880 12588 -13852
rect 12828 -13028 14000 -13000
rect 12828 -13852 13916 -13028
rect 13980 -13852 14000 -13028
rect 12828 -13880 14000 -13852
rect 14240 -13028 15412 -13000
rect 14240 -13852 15328 -13028
rect 15392 -13852 15412 -13028
rect 14240 -13880 15412 -13852
rect 15652 -13028 16824 -13000
rect 15652 -13852 16740 -13028
rect 16804 -13852 16824 -13028
rect 15652 -13880 16824 -13852
rect 17064 -13028 18236 -13000
rect 17064 -13852 18152 -13028
rect 18216 -13852 18236 -13028
rect 17064 -13880 18236 -13852
rect 18476 -13028 19648 -13000
rect 18476 -13852 19564 -13028
rect 19628 -13852 19648 -13028
rect 18476 -13880 19648 -13852
rect 19888 -13028 21060 -13000
rect 19888 -13852 20976 -13028
rect 21040 -13852 21060 -13028
rect 19888 -13880 21060 -13852
rect 21300 -13028 22472 -13000
rect 21300 -13852 22388 -13028
rect 22452 -13852 22472 -13028
rect 21300 -13880 22472 -13852
rect 22712 -13028 23884 -13000
rect 22712 -13852 23800 -13028
rect 23864 -13852 23884 -13028
rect 22712 -13880 23884 -13852
rect -23884 -14148 -22712 -14120
rect -23884 -14972 -22796 -14148
rect -22732 -14972 -22712 -14148
rect -23884 -15000 -22712 -14972
rect -22472 -14148 -21300 -14120
rect -22472 -14972 -21384 -14148
rect -21320 -14972 -21300 -14148
rect -22472 -15000 -21300 -14972
rect -21060 -14148 -19888 -14120
rect -21060 -14972 -19972 -14148
rect -19908 -14972 -19888 -14148
rect -21060 -15000 -19888 -14972
rect -19648 -14148 -18476 -14120
rect -19648 -14972 -18560 -14148
rect -18496 -14972 -18476 -14148
rect -19648 -15000 -18476 -14972
rect -18236 -14148 -17064 -14120
rect -18236 -14972 -17148 -14148
rect -17084 -14972 -17064 -14148
rect -18236 -15000 -17064 -14972
rect -16824 -14148 -15652 -14120
rect -16824 -14972 -15736 -14148
rect -15672 -14972 -15652 -14148
rect -16824 -15000 -15652 -14972
rect -15412 -14148 -14240 -14120
rect -15412 -14972 -14324 -14148
rect -14260 -14972 -14240 -14148
rect -15412 -15000 -14240 -14972
rect -14000 -14148 -12828 -14120
rect -14000 -14972 -12912 -14148
rect -12848 -14972 -12828 -14148
rect -14000 -15000 -12828 -14972
rect -12588 -14148 -11416 -14120
rect -12588 -14972 -11500 -14148
rect -11436 -14972 -11416 -14148
rect -12588 -15000 -11416 -14972
rect -11176 -14148 -10004 -14120
rect -11176 -14972 -10088 -14148
rect -10024 -14972 -10004 -14148
rect -11176 -15000 -10004 -14972
rect -9764 -14148 -8592 -14120
rect -9764 -14972 -8676 -14148
rect -8612 -14972 -8592 -14148
rect -9764 -15000 -8592 -14972
rect -8352 -14148 -7180 -14120
rect -8352 -14972 -7264 -14148
rect -7200 -14972 -7180 -14148
rect -8352 -15000 -7180 -14972
rect -6940 -14148 -5768 -14120
rect -6940 -14972 -5852 -14148
rect -5788 -14972 -5768 -14148
rect -6940 -15000 -5768 -14972
rect -5528 -14148 -4356 -14120
rect -5528 -14972 -4440 -14148
rect -4376 -14972 -4356 -14148
rect -5528 -15000 -4356 -14972
rect -4116 -14148 -2944 -14120
rect -4116 -14972 -3028 -14148
rect -2964 -14972 -2944 -14148
rect -4116 -15000 -2944 -14972
rect -2704 -14148 -1532 -14120
rect -2704 -14972 -1616 -14148
rect -1552 -14972 -1532 -14148
rect -2704 -15000 -1532 -14972
rect -1292 -14148 -120 -14120
rect -1292 -14972 -204 -14148
rect -140 -14972 -120 -14148
rect -1292 -15000 -120 -14972
rect 120 -14148 1292 -14120
rect 120 -14972 1208 -14148
rect 1272 -14972 1292 -14148
rect 120 -15000 1292 -14972
rect 1532 -14148 2704 -14120
rect 1532 -14972 2620 -14148
rect 2684 -14972 2704 -14148
rect 1532 -15000 2704 -14972
rect 2944 -14148 4116 -14120
rect 2944 -14972 4032 -14148
rect 4096 -14972 4116 -14148
rect 2944 -15000 4116 -14972
rect 4356 -14148 5528 -14120
rect 4356 -14972 5444 -14148
rect 5508 -14972 5528 -14148
rect 4356 -15000 5528 -14972
rect 5768 -14148 6940 -14120
rect 5768 -14972 6856 -14148
rect 6920 -14972 6940 -14148
rect 5768 -15000 6940 -14972
rect 7180 -14148 8352 -14120
rect 7180 -14972 8268 -14148
rect 8332 -14972 8352 -14148
rect 7180 -15000 8352 -14972
rect 8592 -14148 9764 -14120
rect 8592 -14972 9680 -14148
rect 9744 -14972 9764 -14148
rect 8592 -15000 9764 -14972
rect 10004 -14148 11176 -14120
rect 10004 -14972 11092 -14148
rect 11156 -14972 11176 -14148
rect 10004 -15000 11176 -14972
rect 11416 -14148 12588 -14120
rect 11416 -14972 12504 -14148
rect 12568 -14972 12588 -14148
rect 11416 -15000 12588 -14972
rect 12828 -14148 14000 -14120
rect 12828 -14972 13916 -14148
rect 13980 -14972 14000 -14148
rect 12828 -15000 14000 -14972
rect 14240 -14148 15412 -14120
rect 14240 -14972 15328 -14148
rect 15392 -14972 15412 -14148
rect 14240 -15000 15412 -14972
rect 15652 -14148 16824 -14120
rect 15652 -14972 16740 -14148
rect 16804 -14972 16824 -14148
rect 15652 -15000 16824 -14972
rect 17064 -14148 18236 -14120
rect 17064 -14972 18152 -14148
rect 18216 -14972 18236 -14148
rect 17064 -15000 18236 -14972
rect 18476 -14148 19648 -14120
rect 18476 -14972 19564 -14148
rect 19628 -14972 19648 -14148
rect 18476 -15000 19648 -14972
rect 19888 -14148 21060 -14120
rect 19888 -14972 20976 -14148
rect 21040 -14972 21060 -14148
rect 19888 -15000 21060 -14972
rect 21300 -14148 22472 -14120
rect 21300 -14972 22388 -14148
rect 22452 -14972 22472 -14148
rect 21300 -15000 22472 -14972
rect 22712 -14148 23884 -14120
rect 22712 -14972 23800 -14148
rect 23864 -14972 23884 -14148
rect 22712 -15000 23884 -14972
rect -23884 -15268 -22712 -15240
rect -23884 -16092 -22796 -15268
rect -22732 -16092 -22712 -15268
rect -23884 -16120 -22712 -16092
rect -22472 -15268 -21300 -15240
rect -22472 -16092 -21384 -15268
rect -21320 -16092 -21300 -15268
rect -22472 -16120 -21300 -16092
rect -21060 -15268 -19888 -15240
rect -21060 -16092 -19972 -15268
rect -19908 -16092 -19888 -15268
rect -21060 -16120 -19888 -16092
rect -19648 -15268 -18476 -15240
rect -19648 -16092 -18560 -15268
rect -18496 -16092 -18476 -15268
rect -19648 -16120 -18476 -16092
rect -18236 -15268 -17064 -15240
rect -18236 -16092 -17148 -15268
rect -17084 -16092 -17064 -15268
rect -18236 -16120 -17064 -16092
rect -16824 -15268 -15652 -15240
rect -16824 -16092 -15736 -15268
rect -15672 -16092 -15652 -15268
rect -16824 -16120 -15652 -16092
rect -15412 -15268 -14240 -15240
rect -15412 -16092 -14324 -15268
rect -14260 -16092 -14240 -15268
rect -15412 -16120 -14240 -16092
rect -14000 -15268 -12828 -15240
rect -14000 -16092 -12912 -15268
rect -12848 -16092 -12828 -15268
rect -14000 -16120 -12828 -16092
rect -12588 -15268 -11416 -15240
rect -12588 -16092 -11500 -15268
rect -11436 -16092 -11416 -15268
rect -12588 -16120 -11416 -16092
rect -11176 -15268 -10004 -15240
rect -11176 -16092 -10088 -15268
rect -10024 -16092 -10004 -15268
rect -11176 -16120 -10004 -16092
rect -9764 -15268 -8592 -15240
rect -9764 -16092 -8676 -15268
rect -8612 -16092 -8592 -15268
rect -9764 -16120 -8592 -16092
rect -8352 -15268 -7180 -15240
rect -8352 -16092 -7264 -15268
rect -7200 -16092 -7180 -15268
rect -8352 -16120 -7180 -16092
rect -6940 -15268 -5768 -15240
rect -6940 -16092 -5852 -15268
rect -5788 -16092 -5768 -15268
rect -6940 -16120 -5768 -16092
rect -5528 -15268 -4356 -15240
rect -5528 -16092 -4440 -15268
rect -4376 -16092 -4356 -15268
rect -5528 -16120 -4356 -16092
rect -4116 -15268 -2944 -15240
rect -4116 -16092 -3028 -15268
rect -2964 -16092 -2944 -15268
rect -4116 -16120 -2944 -16092
rect -2704 -15268 -1532 -15240
rect -2704 -16092 -1616 -15268
rect -1552 -16092 -1532 -15268
rect -2704 -16120 -1532 -16092
rect -1292 -15268 -120 -15240
rect -1292 -16092 -204 -15268
rect -140 -16092 -120 -15268
rect -1292 -16120 -120 -16092
rect 120 -15268 1292 -15240
rect 120 -16092 1208 -15268
rect 1272 -16092 1292 -15268
rect 120 -16120 1292 -16092
rect 1532 -15268 2704 -15240
rect 1532 -16092 2620 -15268
rect 2684 -16092 2704 -15268
rect 1532 -16120 2704 -16092
rect 2944 -15268 4116 -15240
rect 2944 -16092 4032 -15268
rect 4096 -16092 4116 -15268
rect 2944 -16120 4116 -16092
rect 4356 -15268 5528 -15240
rect 4356 -16092 5444 -15268
rect 5508 -16092 5528 -15268
rect 4356 -16120 5528 -16092
rect 5768 -15268 6940 -15240
rect 5768 -16092 6856 -15268
rect 6920 -16092 6940 -15268
rect 5768 -16120 6940 -16092
rect 7180 -15268 8352 -15240
rect 7180 -16092 8268 -15268
rect 8332 -16092 8352 -15268
rect 7180 -16120 8352 -16092
rect 8592 -15268 9764 -15240
rect 8592 -16092 9680 -15268
rect 9744 -16092 9764 -15268
rect 8592 -16120 9764 -16092
rect 10004 -15268 11176 -15240
rect 10004 -16092 11092 -15268
rect 11156 -16092 11176 -15268
rect 10004 -16120 11176 -16092
rect 11416 -15268 12588 -15240
rect 11416 -16092 12504 -15268
rect 12568 -16092 12588 -15268
rect 11416 -16120 12588 -16092
rect 12828 -15268 14000 -15240
rect 12828 -16092 13916 -15268
rect 13980 -16092 14000 -15268
rect 12828 -16120 14000 -16092
rect 14240 -15268 15412 -15240
rect 14240 -16092 15328 -15268
rect 15392 -16092 15412 -15268
rect 14240 -16120 15412 -16092
rect 15652 -15268 16824 -15240
rect 15652 -16092 16740 -15268
rect 16804 -16092 16824 -15268
rect 15652 -16120 16824 -16092
rect 17064 -15268 18236 -15240
rect 17064 -16092 18152 -15268
rect 18216 -16092 18236 -15268
rect 17064 -16120 18236 -16092
rect 18476 -15268 19648 -15240
rect 18476 -16092 19564 -15268
rect 19628 -16092 19648 -15268
rect 18476 -16120 19648 -16092
rect 19888 -15268 21060 -15240
rect 19888 -16092 20976 -15268
rect 21040 -16092 21060 -15268
rect 19888 -16120 21060 -16092
rect 21300 -15268 22472 -15240
rect 21300 -16092 22388 -15268
rect 22452 -16092 22472 -15268
rect 21300 -16120 22472 -16092
rect 22712 -15268 23884 -15240
rect 22712 -16092 23800 -15268
rect 23864 -16092 23884 -15268
rect 22712 -16120 23884 -16092
rect -23884 -16388 -22712 -16360
rect -23884 -17212 -22796 -16388
rect -22732 -17212 -22712 -16388
rect -23884 -17240 -22712 -17212
rect -22472 -16388 -21300 -16360
rect -22472 -17212 -21384 -16388
rect -21320 -17212 -21300 -16388
rect -22472 -17240 -21300 -17212
rect -21060 -16388 -19888 -16360
rect -21060 -17212 -19972 -16388
rect -19908 -17212 -19888 -16388
rect -21060 -17240 -19888 -17212
rect -19648 -16388 -18476 -16360
rect -19648 -17212 -18560 -16388
rect -18496 -17212 -18476 -16388
rect -19648 -17240 -18476 -17212
rect -18236 -16388 -17064 -16360
rect -18236 -17212 -17148 -16388
rect -17084 -17212 -17064 -16388
rect -18236 -17240 -17064 -17212
rect -16824 -16388 -15652 -16360
rect -16824 -17212 -15736 -16388
rect -15672 -17212 -15652 -16388
rect -16824 -17240 -15652 -17212
rect -15412 -16388 -14240 -16360
rect -15412 -17212 -14324 -16388
rect -14260 -17212 -14240 -16388
rect -15412 -17240 -14240 -17212
rect -14000 -16388 -12828 -16360
rect -14000 -17212 -12912 -16388
rect -12848 -17212 -12828 -16388
rect -14000 -17240 -12828 -17212
rect -12588 -16388 -11416 -16360
rect -12588 -17212 -11500 -16388
rect -11436 -17212 -11416 -16388
rect -12588 -17240 -11416 -17212
rect -11176 -16388 -10004 -16360
rect -11176 -17212 -10088 -16388
rect -10024 -17212 -10004 -16388
rect -11176 -17240 -10004 -17212
rect -9764 -16388 -8592 -16360
rect -9764 -17212 -8676 -16388
rect -8612 -17212 -8592 -16388
rect -9764 -17240 -8592 -17212
rect -8352 -16388 -7180 -16360
rect -8352 -17212 -7264 -16388
rect -7200 -17212 -7180 -16388
rect -8352 -17240 -7180 -17212
rect -6940 -16388 -5768 -16360
rect -6940 -17212 -5852 -16388
rect -5788 -17212 -5768 -16388
rect -6940 -17240 -5768 -17212
rect -5528 -16388 -4356 -16360
rect -5528 -17212 -4440 -16388
rect -4376 -17212 -4356 -16388
rect -5528 -17240 -4356 -17212
rect -4116 -16388 -2944 -16360
rect -4116 -17212 -3028 -16388
rect -2964 -17212 -2944 -16388
rect -4116 -17240 -2944 -17212
rect -2704 -16388 -1532 -16360
rect -2704 -17212 -1616 -16388
rect -1552 -17212 -1532 -16388
rect -2704 -17240 -1532 -17212
rect -1292 -16388 -120 -16360
rect -1292 -17212 -204 -16388
rect -140 -17212 -120 -16388
rect -1292 -17240 -120 -17212
rect 120 -16388 1292 -16360
rect 120 -17212 1208 -16388
rect 1272 -17212 1292 -16388
rect 120 -17240 1292 -17212
rect 1532 -16388 2704 -16360
rect 1532 -17212 2620 -16388
rect 2684 -17212 2704 -16388
rect 1532 -17240 2704 -17212
rect 2944 -16388 4116 -16360
rect 2944 -17212 4032 -16388
rect 4096 -17212 4116 -16388
rect 2944 -17240 4116 -17212
rect 4356 -16388 5528 -16360
rect 4356 -17212 5444 -16388
rect 5508 -17212 5528 -16388
rect 4356 -17240 5528 -17212
rect 5768 -16388 6940 -16360
rect 5768 -17212 6856 -16388
rect 6920 -17212 6940 -16388
rect 5768 -17240 6940 -17212
rect 7180 -16388 8352 -16360
rect 7180 -17212 8268 -16388
rect 8332 -17212 8352 -16388
rect 7180 -17240 8352 -17212
rect 8592 -16388 9764 -16360
rect 8592 -17212 9680 -16388
rect 9744 -17212 9764 -16388
rect 8592 -17240 9764 -17212
rect 10004 -16388 11176 -16360
rect 10004 -17212 11092 -16388
rect 11156 -17212 11176 -16388
rect 10004 -17240 11176 -17212
rect 11416 -16388 12588 -16360
rect 11416 -17212 12504 -16388
rect 12568 -17212 12588 -16388
rect 11416 -17240 12588 -17212
rect 12828 -16388 14000 -16360
rect 12828 -17212 13916 -16388
rect 13980 -17212 14000 -16388
rect 12828 -17240 14000 -17212
rect 14240 -16388 15412 -16360
rect 14240 -17212 15328 -16388
rect 15392 -17212 15412 -16388
rect 14240 -17240 15412 -17212
rect 15652 -16388 16824 -16360
rect 15652 -17212 16740 -16388
rect 16804 -17212 16824 -16388
rect 15652 -17240 16824 -17212
rect 17064 -16388 18236 -16360
rect 17064 -17212 18152 -16388
rect 18216 -17212 18236 -16388
rect 17064 -17240 18236 -17212
rect 18476 -16388 19648 -16360
rect 18476 -17212 19564 -16388
rect 19628 -17212 19648 -16388
rect 18476 -17240 19648 -17212
rect 19888 -16388 21060 -16360
rect 19888 -17212 20976 -16388
rect 21040 -17212 21060 -16388
rect 19888 -17240 21060 -17212
rect 21300 -16388 22472 -16360
rect 21300 -17212 22388 -16388
rect 22452 -17212 22472 -16388
rect 21300 -17240 22472 -17212
rect 22712 -16388 23884 -16360
rect 22712 -17212 23800 -16388
rect 23864 -17212 23884 -16388
rect 22712 -17240 23884 -17212
rect -23884 -17508 -22712 -17480
rect -23884 -18332 -22796 -17508
rect -22732 -18332 -22712 -17508
rect -23884 -18360 -22712 -18332
rect -22472 -17508 -21300 -17480
rect -22472 -18332 -21384 -17508
rect -21320 -18332 -21300 -17508
rect -22472 -18360 -21300 -18332
rect -21060 -17508 -19888 -17480
rect -21060 -18332 -19972 -17508
rect -19908 -18332 -19888 -17508
rect -21060 -18360 -19888 -18332
rect -19648 -17508 -18476 -17480
rect -19648 -18332 -18560 -17508
rect -18496 -18332 -18476 -17508
rect -19648 -18360 -18476 -18332
rect -18236 -17508 -17064 -17480
rect -18236 -18332 -17148 -17508
rect -17084 -18332 -17064 -17508
rect -18236 -18360 -17064 -18332
rect -16824 -17508 -15652 -17480
rect -16824 -18332 -15736 -17508
rect -15672 -18332 -15652 -17508
rect -16824 -18360 -15652 -18332
rect -15412 -17508 -14240 -17480
rect -15412 -18332 -14324 -17508
rect -14260 -18332 -14240 -17508
rect -15412 -18360 -14240 -18332
rect -14000 -17508 -12828 -17480
rect -14000 -18332 -12912 -17508
rect -12848 -18332 -12828 -17508
rect -14000 -18360 -12828 -18332
rect -12588 -17508 -11416 -17480
rect -12588 -18332 -11500 -17508
rect -11436 -18332 -11416 -17508
rect -12588 -18360 -11416 -18332
rect -11176 -17508 -10004 -17480
rect -11176 -18332 -10088 -17508
rect -10024 -18332 -10004 -17508
rect -11176 -18360 -10004 -18332
rect -9764 -17508 -8592 -17480
rect -9764 -18332 -8676 -17508
rect -8612 -18332 -8592 -17508
rect -9764 -18360 -8592 -18332
rect -8352 -17508 -7180 -17480
rect -8352 -18332 -7264 -17508
rect -7200 -18332 -7180 -17508
rect -8352 -18360 -7180 -18332
rect -6940 -17508 -5768 -17480
rect -6940 -18332 -5852 -17508
rect -5788 -18332 -5768 -17508
rect -6940 -18360 -5768 -18332
rect -5528 -17508 -4356 -17480
rect -5528 -18332 -4440 -17508
rect -4376 -18332 -4356 -17508
rect -5528 -18360 -4356 -18332
rect -4116 -17508 -2944 -17480
rect -4116 -18332 -3028 -17508
rect -2964 -18332 -2944 -17508
rect -4116 -18360 -2944 -18332
rect -2704 -17508 -1532 -17480
rect -2704 -18332 -1616 -17508
rect -1552 -18332 -1532 -17508
rect -2704 -18360 -1532 -18332
rect -1292 -17508 -120 -17480
rect -1292 -18332 -204 -17508
rect -140 -18332 -120 -17508
rect -1292 -18360 -120 -18332
rect 120 -17508 1292 -17480
rect 120 -18332 1208 -17508
rect 1272 -18332 1292 -17508
rect 120 -18360 1292 -18332
rect 1532 -17508 2704 -17480
rect 1532 -18332 2620 -17508
rect 2684 -18332 2704 -17508
rect 1532 -18360 2704 -18332
rect 2944 -17508 4116 -17480
rect 2944 -18332 4032 -17508
rect 4096 -18332 4116 -17508
rect 2944 -18360 4116 -18332
rect 4356 -17508 5528 -17480
rect 4356 -18332 5444 -17508
rect 5508 -18332 5528 -17508
rect 4356 -18360 5528 -18332
rect 5768 -17508 6940 -17480
rect 5768 -18332 6856 -17508
rect 6920 -18332 6940 -17508
rect 5768 -18360 6940 -18332
rect 7180 -17508 8352 -17480
rect 7180 -18332 8268 -17508
rect 8332 -18332 8352 -17508
rect 7180 -18360 8352 -18332
rect 8592 -17508 9764 -17480
rect 8592 -18332 9680 -17508
rect 9744 -18332 9764 -17508
rect 8592 -18360 9764 -18332
rect 10004 -17508 11176 -17480
rect 10004 -18332 11092 -17508
rect 11156 -18332 11176 -17508
rect 10004 -18360 11176 -18332
rect 11416 -17508 12588 -17480
rect 11416 -18332 12504 -17508
rect 12568 -18332 12588 -17508
rect 11416 -18360 12588 -18332
rect 12828 -17508 14000 -17480
rect 12828 -18332 13916 -17508
rect 13980 -18332 14000 -17508
rect 12828 -18360 14000 -18332
rect 14240 -17508 15412 -17480
rect 14240 -18332 15328 -17508
rect 15392 -18332 15412 -17508
rect 14240 -18360 15412 -18332
rect 15652 -17508 16824 -17480
rect 15652 -18332 16740 -17508
rect 16804 -18332 16824 -17508
rect 15652 -18360 16824 -18332
rect 17064 -17508 18236 -17480
rect 17064 -18332 18152 -17508
rect 18216 -18332 18236 -17508
rect 17064 -18360 18236 -18332
rect 18476 -17508 19648 -17480
rect 18476 -18332 19564 -17508
rect 19628 -18332 19648 -17508
rect 18476 -18360 19648 -18332
rect 19888 -17508 21060 -17480
rect 19888 -18332 20976 -17508
rect 21040 -18332 21060 -17508
rect 19888 -18360 21060 -18332
rect 21300 -17508 22472 -17480
rect 21300 -18332 22388 -17508
rect 22452 -18332 22472 -17508
rect 21300 -18360 22472 -18332
rect 22712 -17508 23884 -17480
rect 22712 -18332 23800 -17508
rect 23864 -18332 23884 -17508
rect 22712 -18360 23884 -18332
<< via3 >>
rect -22796 17508 -22732 18332
rect -21384 17508 -21320 18332
rect -19972 17508 -19908 18332
rect -18560 17508 -18496 18332
rect -17148 17508 -17084 18332
rect -15736 17508 -15672 18332
rect -14324 17508 -14260 18332
rect -12912 17508 -12848 18332
rect -11500 17508 -11436 18332
rect -10088 17508 -10024 18332
rect -8676 17508 -8612 18332
rect -7264 17508 -7200 18332
rect -5852 17508 -5788 18332
rect -4440 17508 -4376 18332
rect -3028 17508 -2964 18332
rect -1616 17508 -1552 18332
rect -204 17508 -140 18332
rect 1208 17508 1272 18332
rect 2620 17508 2684 18332
rect 4032 17508 4096 18332
rect 5444 17508 5508 18332
rect 6856 17508 6920 18332
rect 8268 17508 8332 18332
rect 9680 17508 9744 18332
rect 11092 17508 11156 18332
rect 12504 17508 12568 18332
rect 13916 17508 13980 18332
rect 15328 17508 15392 18332
rect 16740 17508 16804 18332
rect 18152 17508 18216 18332
rect 19564 17508 19628 18332
rect 20976 17508 21040 18332
rect 22388 17508 22452 18332
rect 23800 17508 23864 18332
rect -22796 16388 -22732 17212
rect -21384 16388 -21320 17212
rect -19972 16388 -19908 17212
rect -18560 16388 -18496 17212
rect -17148 16388 -17084 17212
rect -15736 16388 -15672 17212
rect -14324 16388 -14260 17212
rect -12912 16388 -12848 17212
rect -11500 16388 -11436 17212
rect -10088 16388 -10024 17212
rect -8676 16388 -8612 17212
rect -7264 16388 -7200 17212
rect -5852 16388 -5788 17212
rect -4440 16388 -4376 17212
rect -3028 16388 -2964 17212
rect -1616 16388 -1552 17212
rect -204 16388 -140 17212
rect 1208 16388 1272 17212
rect 2620 16388 2684 17212
rect 4032 16388 4096 17212
rect 5444 16388 5508 17212
rect 6856 16388 6920 17212
rect 8268 16388 8332 17212
rect 9680 16388 9744 17212
rect 11092 16388 11156 17212
rect 12504 16388 12568 17212
rect 13916 16388 13980 17212
rect 15328 16388 15392 17212
rect 16740 16388 16804 17212
rect 18152 16388 18216 17212
rect 19564 16388 19628 17212
rect 20976 16388 21040 17212
rect 22388 16388 22452 17212
rect 23800 16388 23864 17212
rect -22796 15268 -22732 16092
rect -21384 15268 -21320 16092
rect -19972 15268 -19908 16092
rect -18560 15268 -18496 16092
rect -17148 15268 -17084 16092
rect -15736 15268 -15672 16092
rect -14324 15268 -14260 16092
rect -12912 15268 -12848 16092
rect -11500 15268 -11436 16092
rect -10088 15268 -10024 16092
rect -8676 15268 -8612 16092
rect -7264 15268 -7200 16092
rect -5852 15268 -5788 16092
rect -4440 15268 -4376 16092
rect -3028 15268 -2964 16092
rect -1616 15268 -1552 16092
rect -204 15268 -140 16092
rect 1208 15268 1272 16092
rect 2620 15268 2684 16092
rect 4032 15268 4096 16092
rect 5444 15268 5508 16092
rect 6856 15268 6920 16092
rect 8268 15268 8332 16092
rect 9680 15268 9744 16092
rect 11092 15268 11156 16092
rect 12504 15268 12568 16092
rect 13916 15268 13980 16092
rect 15328 15268 15392 16092
rect 16740 15268 16804 16092
rect 18152 15268 18216 16092
rect 19564 15268 19628 16092
rect 20976 15268 21040 16092
rect 22388 15268 22452 16092
rect 23800 15268 23864 16092
rect -22796 14148 -22732 14972
rect -21384 14148 -21320 14972
rect -19972 14148 -19908 14972
rect -18560 14148 -18496 14972
rect -17148 14148 -17084 14972
rect -15736 14148 -15672 14972
rect -14324 14148 -14260 14972
rect -12912 14148 -12848 14972
rect -11500 14148 -11436 14972
rect -10088 14148 -10024 14972
rect -8676 14148 -8612 14972
rect -7264 14148 -7200 14972
rect -5852 14148 -5788 14972
rect -4440 14148 -4376 14972
rect -3028 14148 -2964 14972
rect -1616 14148 -1552 14972
rect -204 14148 -140 14972
rect 1208 14148 1272 14972
rect 2620 14148 2684 14972
rect 4032 14148 4096 14972
rect 5444 14148 5508 14972
rect 6856 14148 6920 14972
rect 8268 14148 8332 14972
rect 9680 14148 9744 14972
rect 11092 14148 11156 14972
rect 12504 14148 12568 14972
rect 13916 14148 13980 14972
rect 15328 14148 15392 14972
rect 16740 14148 16804 14972
rect 18152 14148 18216 14972
rect 19564 14148 19628 14972
rect 20976 14148 21040 14972
rect 22388 14148 22452 14972
rect 23800 14148 23864 14972
rect -22796 13028 -22732 13852
rect -21384 13028 -21320 13852
rect -19972 13028 -19908 13852
rect -18560 13028 -18496 13852
rect -17148 13028 -17084 13852
rect -15736 13028 -15672 13852
rect -14324 13028 -14260 13852
rect -12912 13028 -12848 13852
rect -11500 13028 -11436 13852
rect -10088 13028 -10024 13852
rect -8676 13028 -8612 13852
rect -7264 13028 -7200 13852
rect -5852 13028 -5788 13852
rect -4440 13028 -4376 13852
rect -3028 13028 -2964 13852
rect -1616 13028 -1552 13852
rect -204 13028 -140 13852
rect 1208 13028 1272 13852
rect 2620 13028 2684 13852
rect 4032 13028 4096 13852
rect 5444 13028 5508 13852
rect 6856 13028 6920 13852
rect 8268 13028 8332 13852
rect 9680 13028 9744 13852
rect 11092 13028 11156 13852
rect 12504 13028 12568 13852
rect 13916 13028 13980 13852
rect 15328 13028 15392 13852
rect 16740 13028 16804 13852
rect 18152 13028 18216 13852
rect 19564 13028 19628 13852
rect 20976 13028 21040 13852
rect 22388 13028 22452 13852
rect 23800 13028 23864 13852
rect -22796 11908 -22732 12732
rect -21384 11908 -21320 12732
rect -19972 11908 -19908 12732
rect -18560 11908 -18496 12732
rect -17148 11908 -17084 12732
rect -15736 11908 -15672 12732
rect -14324 11908 -14260 12732
rect -12912 11908 -12848 12732
rect -11500 11908 -11436 12732
rect -10088 11908 -10024 12732
rect -8676 11908 -8612 12732
rect -7264 11908 -7200 12732
rect -5852 11908 -5788 12732
rect -4440 11908 -4376 12732
rect -3028 11908 -2964 12732
rect -1616 11908 -1552 12732
rect -204 11908 -140 12732
rect 1208 11908 1272 12732
rect 2620 11908 2684 12732
rect 4032 11908 4096 12732
rect 5444 11908 5508 12732
rect 6856 11908 6920 12732
rect 8268 11908 8332 12732
rect 9680 11908 9744 12732
rect 11092 11908 11156 12732
rect 12504 11908 12568 12732
rect 13916 11908 13980 12732
rect 15328 11908 15392 12732
rect 16740 11908 16804 12732
rect 18152 11908 18216 12732
rect 19564 11908 19628 12732
rect 20976 11908 21040 12732
rect 22388 11908 22452 12732
rect 23800 11908 23864 12732
rect -22796 10788 -22732 11612
rect -21384 10788 -21320 11612
rect -19972 10788 -19908 11612
rect -18560 10788 -18496 11612
rect -17148 10788 -17084 11612
rect -15736 10788 -15672 11612
rect -14324 10788 -14260 11612
rect -12912 10788 -12848 11612
rect -11500 10788 -11436 11612
rect -10088 10788 -10024 11612
rect -8676 10788 -8612 11612
rect -7264 10788 -7200 11612
rect -5852 10788 -5788 11612
rect -4440 10788 -4376 11612
rect -3028 10788 -2964 11612
rect -1616 10788 -1552 11612
rect -204 10788 -140 11612
rect 1208 10788 1272 11612
rect 2620 10788 2684 11612
rect 4032 10788 4096 11612
rect 5444 10788 5508 11612
rect 6856 10788 6920 11612
rect 8268 10788 8332 11612
rect 9680 10788 9744 11612
rect 11092 10788 11156 11612
rect 12504 10788 12568 11612
rect 13916 10788 13980 11612
rect 15328 10788 15392 11612
rect 16740 10788 16804 11612
rect 18152 10788 18216 11612
rect 19564 10788 19628 11612
rect 20976 10788 21040 11612
rect 22388 10788 22452 11612
rect 23800 10788 23864 11612
rect -22796 9668 -22732 10492
rect -21384 9668 -21320 10492
rect -19972 9668 -19908 10492
rect -18560 9668 -18496 10492
rect -17148 9668 -17084 10492
rect -15736 9668 -15672 10492
rect -14324 9668 -14260 10492
rect -12912 9668 -12848 10492
rect -11500 9668 -11436 10492
rect -10088 9668 -10024 10492
rect -8676 9668 -8612 10492
rect -7264 9668 -7200 10492
rect -5852 9668 -5788 10492
rect -4440 9668 -4376 10492
rect -3028 9668 -2964 10492
rect -1616 9668 -1552 10492
rect -204 9668 -140 10492
rect 1208 9668 1272 10492
rect 2620 9668 2684 10492
rect 4032 9668 4096 10492
rect 5444 9668 5508 10492
rect 6856 9668 6920 10492
rect 8268 9668 8332 10492
rect 9680 9668 9744 10492
rect 11092 9668 11156 10492
rect 12504 9668 12568 10492
rect 13916 9668 13980 10492
rect 15328 9668 15392 10492
rect 16740 9668 16804 10492
rect 18152 9668 18216 10492
rect 19564 9668 19628 10492
rect 20976 9668 21040 10492
rect 22388 9668 22452 10492
rect 23800 9668 23864 10492
rect -22796 8548 -22732 9372
rect -21384 8548 -21320 9372
rect -19972 8548 -19908 9372
rect -18560 8548 -18496 9372
rect -17148 8548 -17084 9372
rect -15736 8548 -15672 9372
rect -14324 8548 -14260 9372
rect -12912 8548 -12848 9372
rect -11500 8548 -11436 9372
rect -10088 8548 -10024 9372
rect -8676 8548 -8612 9372
rect -7264 8548 -7200 9372
rect -5852 8548 -5788 9372
rect -4440 8548 -4376 9372
rect -3028 8548 -2964 9372
rect -1616 8548 -1552 9372
rect -204 8548 -140 9372
rect 1208 8548 1272 9372
rect 2620 8548 2684 9372
rect 4032 8548 4096 9372
rect 5444 8548 5508 9372
rect 6856 8548 6920 9372
rect 8268 8548 8332 9372
rect 9680 8548 9744 9372
rect 11092 8548 11156 9372
rect 12504 8548 12568 9372
rect 13916 8548 13980 9372
rect 15328 8548 15392 9372
rect 16740 8548 16804 9372
rect 18152 8548 18216 9372
rect 19564 8548 19628 9372
rect 20976 8548 21040 9372
rect 22388 8548 22452 9372
rect 23800 8548 23864 9372
rect -22796 7428 -22732 8252
rect -21384 7428 -21320 8252
rect -19972 7428 -19908 8252
rect -18560 7428 -18496 8252
rect -17148 7428 -17084 8252
rect -15736 7428 -15672 8252
rect -14324 7428 -14260 8252
rect -12912 7428 -12848 8252
rect -11500 7428 -11436 8252
rect -10088 7428 -10024 8252
rect -8676 7428 -8612 8252
rect -7264 7428 -7200 8252
rect -5852 7428 -5788 8252
rect -4440 7428 -4376 8252
rect -3028 7428 -2964 8252
rect -1616 7428 -1552 8252
rect -204 7428 -140 8252
rect 1208 7428 1272 8252
rect 2620 7428 2684 8252
rect 4032 7428 4096 8252
rect 5444 7428 5508 8252
rect 6856 7428 6920 8252
rect 8268 7428 8332 8252
rect 9680 7428 9744 8252
rect 11092 7428 11156 8252
rect 12504 7428 12568 8252
rect 13916 7428 13980 8252
rect 15328 7428 15392 8252
rect 16740 7428 16804 8252
rect 18152 7428 18216 8252
rect 19564 7428 19628 8252
rect 20976 7428 21040 8252
rect 22388 7428 22452 8252
rect 23800 7428 23864 8252
rect -22796 6308 -22732 7132
rect -21384 6308 -21320 7132
rect -19972 6308 -19908 7132
rect -18560 6308 -18496 7132
rect -17148 6308 -17084 7132
rect -15736 6308 -15672 7132
rect -14324 6308 -14260 7132
rect -12912 6308 -12848 7132
rect -11500 6308 -11436 7132
rect -10088 6308 -10024 7132
rect -8676 6308 -8612 7132
rect -7264 6308 -7200 7132
rect -5852 6308 -5788 7132
rect -4440 6308 -4376 7132
rect -3028 6308 -2964 7132
rect -1616 6308 -1552 7132
rect -204 6308 -140 7132
rect 1208 6308 1272 7132
rect 2620 6308 2684 7132
rect 4032 6308 4096 7132
rect 5444 6308 5508 7132
rect 6856 6308 6920 7132
rect 8268 6308 8332 7132
rect 9680 6308 9744 7132
rect 11092 6308 11156 7132
rect 12504 6308 12568 7132
rect 13916 6308 13980 7132
rect 15328 6308 15392 7132
rect 16740 6308 16804 7132
rect 18152 6308 18216 7132
rect 19564 6308 19628 7132
rect 20976 6308 21040 7132
rect 22388 6308 22452 7132
rect 23800 6308 23864 7132
rect -22796 5188 -22732 6012
rect -21384 5188 -21320 6012
rect -19972 5188 -19908 6012
rect -18560 5188 -18496 6012
rect -17148 5188 -17084 6012
rect -15736 5188 -15672 6012
rect -14324 5188 -14260 6012
rect -12912 5188 -12848 6012
rect -11500 5188 -11436 6012
rect -10088 5188 -10024 6012
rect -8676 5188 -8612 6012
rect -7264 5188 -7200 6012
rect -5852 5188 -5788 6012
rect -4440 5188 -4376 6012
rect -3028 5188 -2964 6012
rect -1616 5188 -1552 6012
rect -204 5188 -140 6012
rect 1208 5188 1272 6012
rect 2620 5188 2684 6012
rect 4032 5188 4096 6012
rect 5444 5188 5508 6012
rect 6856 5188 6920 6012
rect 8268 5188 8332 6012
rect 9680 5188 9744 6012
rect 11092 5188 11156 6012
rect 12504 5188 12568 6012
rect 13916 5188 13980 6012
rect 15328 5188 15392 6012
rect 16740 5188 16804 6012
rect 18152 5188 18216 6012
rect 19564 5188 19628 6012
rect 20976 5188 21040 6012
rect 22388 5188 22452 6012
rect 23800 5188 23864 6012
rect -22796 4068 -22732 4892
rect -21384 4068 -21320 4892
rect -19972 4068 -19908 4892
rect -18560 4068 -18496 4892
rect -17148 4068 -17084 4892
rect -15736 4068 -15672 4892
rect -14324 4068 -14260 4892
rect -12912 4068 -12848 4892
rect -11500 4068 -11436 4892
rect -10088 4068 -10024 4892
rect -8676 4068 -8612 4892
rect -7264 4068 -7200 4892
rect -5852 4068 -5788 4892
rect -4440 4068 -4376 4892
rect -3028 4068 -2964 4892
rect -1616 4068 -1552 4892
rect -204 4068 -140 4892
rect 1208 4068 1272 4892
rect 2620 4068 2684 4892
rect 4032 4068 4096 4892
rect 5444 4068 5508 4892
rect 6856 4068 6920 4892
rect 8268 4068 8332 4892
rect 9680 4068 9744 4892
rect 11092 4068 11156 4892
rect 12504 4068 12568 4892
rect 13916 4068 13980 4892
rect 15328 4068 15392 4892
rect 16740 4068 16804 4892
rect 18152 4068 18216 4892
rect 19564 4068 19628 4892
rect 20976 4068 21040 4892
rect 22388 4068 22452 4892
rect 23800 4068 23864 4892
rect -22796 2948 -22732 3772
rect -21384 2948 -21320 3772
rect -19972 2948 -19908 3772
rect -18560 2948 -18496 3772
rect -17148 2948 -17084 3772
rect -15736 2948 -15672 3772
rect -14324 2948 -14260 3772
rect -12912 2948 -12848 3772
rect -11500 2948 -11436 3772
rect -10088 2948 -10024 3772
rect -8676 2948 -8612 3772
rect -7264 2948 -7200 3772
rect -5852 2948 -5788 3772
rect -4440 2948 -4376 3772
rect -3028 2948 -2964 3772
rect -1616 2948 -1552 3772
rect -204 2948 -140 3772
rect 1208 2948 1272 3772
rect 2620 2948 2684 3772
rect 4032 2948 4096 3772
rect 5444 2948 5508 3772
rect 6856 2948 6920 3772
rect 8268 2948 8332 3772
rect 9680 2948 9744 3772
rect 11092 2948 11156 3772
rect 12504 2948 12568 3772
rect 13916 2948 13980 3772
rect 15328 2948 15392 3772
rect 16740 2948 16804 3772
rect 18152 2948 18216 3772
rect 19564 2948 19628 3772
rect 20976 2948 21040 3772
rect 22388 2948 22452 3772
rect 23800 2948 23864 3772
rect -22796 1828 -22732 2652
rect -21384 1828 -21320 2652
rect -19972 1828 -19908 2652
rect -18560 1828 -18496 2652
rect -17148 1828 -17084 2652
rect -15736 1828 -15672 2652
rect -14324 1828 -14260 2652
rect -12912 1828 -12848 2652
rect -11500 1828 -11436 2652
rect -10088 1828 -10024 2652
rect -8676 1828 -8612 2652
rect -7264 1828 -7200 2652
rect -5852 1828 -5788 2652
rect -4440 1828 -4376 2652
rect -3028 1828 -2964 2652
rect -1616 1828 -1552 2652
rect -204 1828 -140 2652
rect 1208 1828 1272 2652
rect 2620 1828 2684 2652
rect 4032 1828 4096 2652
rect 5444 1828 5508 2652
rect 6856 1828 6920 2652
rect 8268 1828 8332 2652
rect 9680 1828 9744 2652
rect 11092 1828 11156 2652
rect 12504 1828 12568 2652
rect 13916 1828 13980 2652
rect 15328 1828 15392 2652
rect 16740 1828 16804 2652
rect 18152 1828 18216 2652
rect 19564 1828 19628 2652
rect 20976 1828 21040 2652
rect 22388 1828 22452 2652
rect 23800 1828 23864 2652
rect -22796 708 -22732 1532
rect -21384 708 -21320 1532
rect -19972 708 -19908 1532
rect -18560 708 -18496 1532
rect -17148 708 -17084 1532
rect -15736 708 -15672 1532
rect -14324 708 -14260 1532
rect -12912 708 -12848 1532
rect -11500 708 -11436 1532
rect -10088 708 -10024 1532
rect -8676 708 -8612 1532
rect -7264 708 -7200 1532
rect -5852 708 -5788 1532
rect -4440 708 -4376 1532
rect -3028 708 -2964 1532
rect -1616 708 -1552 1532
rect -204 708 -140 1532
rect 1208 708 1272 1532
rect 2620 708 2684 1532
rect 4032 708 4096 1532
rect 5444 708 5508 1532
rect 6856 708 6920 1532
rect 8268 708 8332 1532
rect 9680 708 9744 1532
rect 11092 708 11156 1532
rect 12504 708 12568 1532
rect 13916 708 13980 1532
rect 15328 708 15392 1532
rect 16740 708 16804 1532
rect 18152 708 18216 1532
rect 19564 708 19628 1532
rect 20976 708 21040 1532
rect 22388 708 22452 1532
rect 23800 708 23864 1532
rect -22796 -412 -22732 412
rect -21384 -412 -21320 412
rect -19972 -412 -19908 412
rect -18560 -412 -18496 412
rect -17148 -412 -17084 412
rect -15736 -412 -15672 412
rect -14324 -412 -14260 412
rect -12912 -412 -12848 412
rect -11500 -412 -11436 412
rect -10088 -412 -10024 412
rect -8676 -412 -8612 412
rect -7264 -412 -7200 412
rect -5852 -412 -5788 412
rect -4440 -412 -4376 412
rect -3028 -412 -2964 412
rect -1616 -412 -1552 412
rect -204 -412 -140 412
rect 1208 -412 1272 412
rect 2620 -412 2684 412
rect 4032 -412 4096 412
rect 5444 -412 5508 412
rect 6856 -412 6920 412
rect 8268 -412 8332 412
rect 9680 -412 9744 412
rect 11092 -412 11156 412
rect 12504 -412 12568 412
rect 13916 -412 13980 412
rect 15328 -412 15392 412
rect 16740 -412 16804 412
rect 18152 -412 18216 412
rect 19564 -412 19628 412
rect 20976 -412 21040 412
rect 22388 -412 22452 412
rect 23800 -412 23864 412
rect -22796 -1532 -22732 -708
rect -21384 -1532 -21320 -708
rect -19972 -1532 -19908 -708
rect -18560 -1532 -18496 -708
rect -17148 -1532 -17084 -708
rect -15736 -1532 -15672 -708
rect -14324 -1532 -14260 -708
rect -12912 -1532 -12848 -708
rect -11500 -1532 -11436 -708
rect -10088 -1532 -10024 -708
rect -8676 -1532 -8612 -708
rect -7264 -1532 -7200 -708
rect -5852 -1532 -5788 -708
rect -4440 -1532 -4376 -708
rect -3028 -1532 -2964 -708
rect -1616 -1532 -1552 -708
rect -204 -1532 -140 -708
rect 1208 -1532 1272 -708
rect 2620 -1532 2684 -708
rect 4032 -1532 4096 -708
rect 5444 -1532 5508 -708
rect 6856 -1532 6920 -708
rect 8268 -1532 8332 -708
rect 9680 -1532 9744 -708
rect 11092 -1532 11156 -708
rect 12504 -1532 12568 -708
rect 13916 -1532 13980 -708
rect 15328 -1532 15392 -708
rect 16740 -1532 16804 -708
rect 18152 -1532 18216 -708
rect 19564 -1532 19628 -708
rect 20976 -1532 21040 -708
rect 22388 -1532 22452 -708
rect 23800 -1532 23864 -708
rect -22796 -2652 -22732 -1828
rect -21384 -2652 -21320 -1828
rect -19972 -2652 -19908 -1828
rect -18560 -2652 -18496 -1828
rect -17148 -2652 -17084 -1828
rect -15736 -2652 -15672 -1828
rect -14324 -2652 -14260 -1828
rect -12912 -2652 -12848 -1828
rect -11500 -2652 -11436 -1828
rect -10088 -2652 -10024 -1828
rect -8676 -2652 -8612 -1828
rect -7264 -2652 -7200 -1828
rect -5852 -2652 -5788 -1828
rect -4440 -2652 -4376 -1828
rect -3028 -2652 -2964 -1828
rect -1616 -2652 -1552 -1828
rect -204 -2652 -140 -1828
rect 1208 -2652 1272 -1828
rect 2620 -2652 2684 -1828
rect 4032 -2652 4096 -1828
rect 5444 -2652 5508 -1828
rect 6856 -2652 6920 -1828
rect 8268 -2652 8332 -1828
rect 9680 -2652 9744 -1828
rect 11092 -2652 11156 -1828
rect 12504 -2652 12568 -1828
rect 13916 -2652 13980 -1828
rect 15328 -2652 15392 -1828
rect 16740 -2652 16804 -1828
rect 18152 -2652 18216 -1828
rect 19564 -2652 19628 -1828
rect 20976 -2652 21040 -1828
rect 22388 -2652 22452 -1828
rect 23800 -2652 23864 -1828
rect -22796 -3772 -22732 -2948
rect -21384 -3772 -21320 -2948
rect -19972 -3772 -19908 -2948
rect -18560 -3772 -18496 -2948
rect -17148 -3772 -17084 -2948
rect -15736 -3772 -15672 -2948
rect -14324 -3772 -14260 -2948
rect -12912 -3772 -12848 -2948
rect -11500 -3772 -11436 -2948
rect -10088 -3772 -10024 -2948
rect -8676 -3772 -8612 -2948
rect -7264 -3772 -7200 -2948
rect -5852 -3772 -5788 -2948
rect -4440 -3772 -4376 -2948
rect -3028 -3772 -2964 -2948
rect -1616 -3772 -1552 -2948
rect -204 -3772 -140 -2948
rect 1208 -3772 1272 -2948
rect 2620 -3772 2684 -2948
rect 4032 -3772 4096 -2948
rect 5444 -3772 5508 -2948
rect 6856 -3772 6920 -2948
rect 8268 -3772 8332 -2948
rect 9680 -3772 9744 -2948
rect 11092 -3772 11156 -2948
rect 12504 -3772 12568 -2948
rect 13916 -3772 13980 -2948
rect 15328 -3772 15392 -2948
rect 16740 -3772 16804 -2948
rect 18152 -3772 18216 -2948
rect 19564 -3772 19628 -2948
rect 20976 -3772 21040 -2948
rect 22388 -3772 22452 -2948
rect 23800 -3772 23864 -2948
rect -22796 -4892 -22732 -4068
rect -21384 -4892 -21320 -4068
rect -19972 -4892 -19908 -4068
rect -18560 -4892 -18496 -4068
rect -17148 -4892 -17084 -4068
rect -15736 -4892 -15672 -4068
rect -14324 -4892 -14260 -4068
rect -12912 -4892 -12848 -4068
rect -11500 -4892 -11436 -4068
rect -10088 -4892 -10024 -4068
rect -8676 -4892 -8612 -4068
rect -7264 -4892 -7200 -4068
rect -5852 -4892 -5788 -4068
rect -4440 -4892 -4376 -4068
rect -3028 -4892 -2964 -4068
rect -1616 -4892 -1552 -4068
rect -204 -4892 -140 -4068
rect 1208 -4892 1272 -4068
rect 2620 -4892 2684 -4068
rect 4032 -4892 4096 -4068
rect 5444 -4892 5508 -4068
rect 6856 -4892 6920 -4068
rect 8268 -4892 8332 -4068
rect 9680 -4892 9744 -4068
rect 11092 -4892 11156 -4068
rect 12504 -4892 12568 -4068
rect 13916 -4892 13980 -4068
rect 15328 -4892 15392 -4068
rect 16740 -4892 16804 -4068
rect 18152 -4892 18216 -4068
rect 19564 -4892 19628 -4068
rect 20976 -4892 21040 -4068
rect 22388 -4892 22452 -4068
rect 23800 -4892 23864 -4068
rect -22796 -6012 -22732 -5188
rect -21384 -6012 -21320 -5188
rect -19972 -6012 -19908 -5188
rect -18560 -6012 -18496 -5188
rect -17148 -6012 -17084 -5188
rect -15736 -6012 -15672 -5188
rect -14324 -6012 -14260 -5188
rect -12912 -6012 -12848 -5188
rect -11500 -6012 -11436 -5188
rect -10088 -6012 -10024 -5188
rect -8676 -6012 -8612 -5188
rect -7264 -6012 -7200 -5188
rect -5852 -6012 -5788 -5188
rect -4440 -6012 -4376 -5188
rect -3028 -6012 -2964 -5188
rect -1616 -6012 -1552 -5188
rect -204 -6012 -140 -5188
rect 1208 -6012 1272 -5188
rect 2620 -6012 2684 -5188
rect 4032 -6012 4096 -5188
rect 5444 -6012 5508 -5188
rect 6856 -6012 6920 -5188
rect 8268 -6012 8332 -5188
rect 9680 -6012 9744 -5188
rect 11092 -6012 11156 -5188
rect 12504 -6012 12568 -5188
rect 13916 -6012 13980 -5188
rect 15328 -6012 15392 -5188
rect 16740 -6012 16804 -5188
rect 18152 -6012 18216 -5188
rect 19564 -6012 19628 -5188
rect 20976 -6012 21040 -5188
rect 22388 -6012 22452 -5188
rect 23800 -6012 23864 -5188
rect -22796 -7132 -22732 -6308
rect -21384 -7132 -21320 -6308
rect -19972 -7132 -19908 -6308
rect -18560 -7132 -18496 -6308
rect -17148 -7132 -17084 -6308
rect -15736 -7132 -15672 -6308
rect -14324 -7132 -14260 -6308
rect -12912 -7132 -12848 -6308
rect -11500 -7132 -11436 -6308
rect -10088 -7132 -10024 -6308
rect -8676 -7132 -8612 -6308
rect -7264 -7132 -7200 -6308
rect -5852 -7132 -5788 -6308
rect -4440 -7132 -4376 -6308
rect -3028 -7132 -2964 -6308
rect -1616 -7132 -1552 -6308
rect -204 -7132 -140 -6308
rect 1208 -7132 1272 -6308
rect 2620 -7132 2684 -6308
rect 4032 -7132 4096 -6308
rect 5444 -7132 5508 -6308
rect 6856 -7132 6920 -6308
rect 8268 -7132 8332 -6308
rect 9680 -7132 9744 -6308
rect 11092 -7132 11156 -6308
rect 12504 -7132 12568 -6308
rect 13916 -7132 13980 -6308
rect 15328 -7132 15392 -6308
rect 16740 -7132 16804 -6308
rect 18152 -7132 18216 -6308
rect 19564 -7132 19628 -6308
rect 20976 -7132 21040 -6308
rect 22388 -7132 22452 -6308
rect 23800 -7132 23864 -6308
rect -22796 -8252 -22732 -7428
rect -21384 -8252 -21320 -7428
rect -19972 -8252 -19908 -7428
rect -18560 -8252 -18496 -7428
rect -17148 -8252 -17084 -7428
rect -15736 -8252 -15672 -7428
rect -14324 -8252 -14260 -7428
rect -12912 -8252 -12848 -7428
rect -11500 -8252 -11436 -7428
rect -10088 -8252 -10024 -7428
rect -8676 -8252 -8612 -7428
rect -7264 -8252 -7200 -7428
rect -5852 -8252 -5788 -7428
rect -4440 -8252 -4376 -7428
rect -3028 -8252 -2964 -7428
rect -1616 -8252 -1552 -7428
rect -204 -8252 -140 -7428
rect 1208 -8252 1272 -7428
rect 2620 -8252 2684 -7428
rect 4032 -8252 4096 -7428
rect 5444 -8252 5508 -7428
rect 6856 -8252 6920 -7428
rect 8268 -8252 8332 -7428
rect 9680 -8252 9744 -7428
rect 11092 -8252 11156 -7428
rect 12504 -8252 12568 -7428
rect 13916 -8252 13980 -7428
rect 15328 -8252 15392 -7428
rect 16740 -8252 16804 -7428
rect 18152 -8252 18216 -7428
rect 19564 -8252 19628 -7428
rect 20976 -8252 21040 -7428
rect 22388 -8252 22452 -7428
rect 23800 -8252 23864 -7428
rect -22796 -9372 -22732 -8548
rect -21384 -9372 -21320 -8548
rect -19972 -9372 -19908 -8548
rect -18560 -9372 -18496 -8548
rect -17148 -9372 -17084 -8548
rect -15736 -9372 -15672 -8548
rect -14324 -9372 -14260 -8548
rect -12912 -9372 -12848 -8548
rect -11500 -9372 -11436 -8548
rect -10088 -9372 -10024 -8548
rect -8676 -9372 -8612 -8548
rect -7264 -9372 -7200 -8548
rect -5852 -9372 -5788 -8548
rect -4440 -9372 -4376 -8548
rect -3028 -9372 -2964 -8548
rect -1616 -9372 -1552 -8548
rect -204 -9372 -140 -8548
rect 1208 -9372 1272 -8548
rect 2620 -9372 2684 -8548
rect 4032 -9372 4096 -8548
rect 5444 -9372 5508 -8548
rect 6856 -9372 6920 -8548
rect 8268 -9372 8332 -8548
rect 9680 -9372 9744 -8548
rect 11092 -9372 11156 -8548
rect 12504 -9372 12568 -8548
rect 13916 -9372 13980 -8548
rect 15328 -9372 15392 -8548
rect 16740 -9372 16804 -8548
rect 18152 -9372 18216 -8548
rect 19564 -9372 19628 -8548
rect 20976 -9372 21040 -8548
rect 22388 -9372 22452 -8548
rect 23800 -9372 23864 -8548
rect -22796 -10492 -22732 -9668
rect -21384 -10492 -21320 -9668
rect -19972 -10492 -19908 -9668
rect -18560 -10492 -18496 -9668
rect -17148 -10492 -17084 -9668
rect -15736 -10492 -15672 -9668
rect -14324 -10492 -14260 -9668
rect -12912 -10492 -12848 -9668
rect -11500 -10492 -11436 -9668
rect -10088 -10492 -10024 -9668
rect -8676 -10492 -8612 -9668
rect -7264 -10492 -7200 -9668
rect -5852 -10492 -5788 -9668
rect -4440 -10492 -4376 -9668
rect -3028 -10492 -2964 -9668
rect -1616 -10492 -1552 -9668
rect -204 -10492 -140 -9668
rect 1208 -10492 1272 -9668
rect 2620 -10492 2684 -9668
rect 4032 -10492 4096 -9668
rect 5444 -10492 5508 -9668
rect 6856 -10492 6920 -9668
rect 8268 -10492 8332 -9668
rect 9680 -10492 9744 -9668
rect 11092 -10492 11156 -9668
rect 12504 -10492 12568 -9668
rect 13916 -10492 13980 -9668
rect 15328 -10492 15392 -9668
rect 16740 -10492 16804 -9668
rect 18152 -10492 18216 -9668
rect 19564 -10492 19628 -9668
rect 20976 -10492 21040 -9668
rect 22388 -10492 22452 -9668
rect 23800 -10492 23864 -9668
rect -22796 -11612 -22732 -10788
rect -21384 -11612 -21320 -10788
rect -19972 -11612 -19908 -10788
rect -18560 -11612 -18496 -10788
rect -17148 -11612 -17084 -10788
rect -15736 -11612 -15672 -10788
rect -14324 -11612 -14260 -10788
rect -12912 -11612 -12848 -10788
rect -11500 -11612 -11436 -10788
rect -10088 -11612 -10024 -10788
rect -8676 -11612 -8612 -10788
rect -7264 -11612 -7200 -10788
rect -5852 -11612 -5788 -10788
rect -4440 -11612 -4376 -10788
rect -3028 -11612 -2964 -10788
rect -1616 -11612 -1552 -10788
rect -204 -11612 -140 -10788
rect 1208 -11612 1272 -10788
rect 2620 -11612 2684 -10788
rect 4032 -11612 4096 -10788
rect 5444 -11612 5508 -10788
rect 6856 -11612 6920 -10788
rect 8268 -11612 8332 -10788
rect 9680 -11612 9744 -10788
rect 11092 -11612 11156 -10788
rect 12504 -11612 12568 -10788
rect 13916 -11612 13980 -10788
rect 15328 -11612 15392 -10788
rect 16740 -11612 16804 -10788
rect 18152 -11612 18216 -10788
rect 19564 -11612 19628 -10788
rect 20976 -11612 21040 -10788
rect 22388 -11612 22452 -10788
rect 23800 -11612 23864 -10788
rect -22796 -12732 -22732 -11908
rect -21384 -12732 -21320 -11908
rect -19972 -12732 -19908 -11908
rect -18560 -12732 -18496 -11908
rect -17148 -12732 -17084 -11908
rect -15736 -12732 -15672 -11908
rect -14324 -12732 -14260 -11908
rect -12912 -12732 -12848 -11908
rect -11500 -12732 -11436 -11908
rect -10088 -12732 -10024 -11908
rect -8676 -12732 -8612 -11908
rect -7264 -12732 -7200 -11908
rect -5852 -12732 -5788 -11908
rect -4440 -12732 -4376 -11908
rect -3028 -12732 -2964 -11908
rect -1616 -12732 -1552 -11908
rect -204 -12732 -140 -11908
rect 1208 -12732 1272 -11908
rect 2620 -12732 2684 -11908
rect 4032 -12732 4096 -11908
rect 5444 -12732 5508 -11908
rect 6856 -12732 6920 -11908
rect 8268 -12732 8332 -11908
rect 9680 -12732 9744 -11908
rect 11092 -12732 11156 -11908
rect 12504 -12732 12568 -11908
rect 13916 -12732 13980 -11908
rect 15328 -12732 15392 -11908
rect 16740 -12732 16804 -11908
rect 18152 -12732 18216 -11908
rect 19564 -12732 19628 -11908
rect 20976 -12732 21040 -11908
rect 22388 -12732 22452 -11908
rect 23800 -12732 23864 -11908
rect -22796 -13852 -22732 -13028
rect -21384 -13852 -21320 -13028
rect -19972 -13852 -19908 -13028
rect -18560 -13852 -18496 -13028
rect -17148 -13852 -17084 -13028
rect -15736 -13852 -15672 -13028
rect -14324 -13852 -14260 -13028
rect -12912 -13852 -12848 -13028
rect -11500 -13852 -11436 -13028
rect -10088 -13852 -10024 -13028
rect -8676 -13852 -8612 -13028
rect -7264 -13852 -7200 -13028
rect -5852 -13852 -5788 -13028
rect -4440 -13852 -4376 -13028
rect -3028 -13852 -2964 -13028
rect -1616 -13852 -1552 -13028
rect -204 -13852 -140 -13028
rect 1208 -13852 1272 -13028
rect 2620 -13852 2684 -13028
rect 4032 -13852 4096 -13028
rect 5444 -13852 5508 -13028
rect 6856 -13852 6920 -13028
rect 8268 -13852 8332 -13028
rect 9680 -13852 9744 -13028
rect 11092 -13852 11156 -13028
rect 12504 -13852 12568 -13028
rect 13916 -13852 13980 -13028
rect 15328 -13852 15392 -13028
rect 16740 -13852 16804 -13028
rect 18152 -13852 18216 -13028
rect 19564 -13852 19628 -13028
rect 20976 -13852 21040 -13028
rect 22388 -13852 22452 -13028
rect 23800 -13852 23864 -13028
rect -22796 -14972 -22732 -14148
rect -21384 -14972 -21320 -14148
rect -19972 -14972 -19908 -14148
rect -18560 -14972 -18496 -14148
rect -17148 -14972 -17084 -14148
rect -15736 -14972 -15672 -14148
rect -14324 -14972 -14260 -14148
rect -12912 -14972 -12848 -14148
rect -11500 -14972 -11436 -14148
rect -10088 -14972 -10024 -14148
rect -8676 -14972 -8612 -14148
rect -7264 -14972 -7200 -14148
rect -5852 -14972 -5788 -14148
rect -4440 -14972 -4376 -14148
rect -3028 -14972 -2964 -14148
rect -1616 -14972 -1552 -14148
rect -204 -14972 -140 -14148
rect 1208 -14972 1272 -14148
rect 2620 -14972 2684 -14148
rect 4032 -14972 4096 -14148
rect 5444 -14972 5508 -14148
rect 6856 -14972 6920 -14148
rect 8268 -14972 8332 -14148
rect 9680 -14972 9744 -14148
rect 11092 -14972 11156 -14148
rect 12504 -14972 12568 -14148
rect 13916 -14972 13980 -14148
rect 15328 -14972 15392 -14148
rect 16740 -14972 16804 -14148
rect 18152 -14972 18216 -14148
rect 19564 -14972 19628 -14148
rect 20976 -14972 21040 -14148
rect 22388 -14972 22452 -14148
rect 23800 -14972 23864 -14148
rect -22796 -16092 -22732 -15268
rect -21384 -16092 -21320 -15268
rect -19972 -16092 -19908 -15268
rect -18560 -16092 -18496 -15268
rect -17148 -16092 -17084 -15268
rect -15736 -16092 -15672 -15268
rect -14324 -16092 -14260 -15268
rect -12912 -16092 -12848 -15268
rect -11500 -16092 -11436 -15268
rect -10088 -16092 -10024 -15268
rect -8676 -16092 -8612 -15268
rect -7264 -16092 -7200 -15268
rect -5852 -16092 -5788 -15268
rect -4440 -16092 -4376 -15268
rect -3028 -16092 -2964 -15268
rect -1616 -16092 -1552 -15268
rect -204 -16092 -140 -15268
rect 1208 -16092 1272 -15268
rect 2620 -16092 2684 -15268
rect 4032 -16092 4096 -15268
rect 5444 -16092 5508 -15268
rect 6856 -16092 6920 -15268
rect 8268 -16092 8332 -15268
rect 9680 -16092 9744 -15268
rect 11092 -16092 11156 -15268
rect 12504 -16092 12568 -15268
rect 13916 -16092 13980 -15268
rect 15328 -16092 15392 -15268
rect 16740 -16092 16804 -15268
rect 18152 -16092 18216 -15268
rect 19564 -16092 19628 -15268
rect 20976 -16092 21040 -15268
rect 22388 -16092 22452 -15268
rect 23800 -16092 23864 -15268
rect -22796 -17212 -22732 -16388
rect -21384 -17212 -21320 -16388
rect -19972 -17212 -19908 -16388
rect -18560 -17212 -18496 -16388
rect -17148 -17212 -17084 -16388
rect -15736 -17212 -15672 -16388
rect -14324 -17212 -14260 -16388
rect -12912 -17212 -12848 -16388
rect -11500 -17212 -11436 -16388
rect -10088 -17212 -10024 -16388
rect -8676 -17212 -8612 -16388
rect -7264 -17212 -7200 -16388
rect -5852 -17212 -5788 -16388
rect -4440 -17212 -4376 -16388
rect -3028 -17212 -2964 -16388
rect -1616 -17212 -1552 -16388
rect -204 -17212 -140 -16388
rect 1208 -17212 1272 -16388
rect 2620 -17212 2684 -16388
rect 4032 -17212 4096 -16388
rect 5444 -17212 5508 -16388
rect 6856 -17212 6920 -16388
rect 8268 -17212 8332 -16388
rect 9680 -17212 9744 -16388
rect 11092 -17212 11156 -16388
rect 12504 -17212 12568 -16388
rect 13916 -17212 13980 -16388
rect 15328 -17212 15392 -16388
rect 16740 -17212 16804 -16388
rect 18152 -17212 18216 -16388
rect 19564 -17212 19628 -16388
rect 20976 -17212 21040 -16388
rect 22388 -17212 22452 -16388
rect 23800 -17212 23864 -16388
rect -22796 -18332 -22732 -17508
rect -21384 -18332 -21320 -17508
rect -19972 -18332 -19908 -17508
rect -18560 -18332 -18496 -17508
rect -17148 -18332 -17084 -17508
rect -15736 -18332 -15672 -17508
rect -14324 -18332 -14260 -17508
rect -12912 -18332 -12848 -17508
rect -11500 -18332 -11436 -17508
rect -10088 -18332 -10024 -17508
rect -8676 -18332 -8612 -17508
rect -7264 -18332 -7200 -17508
rect -5852 -18332 -5788 -17508
rect -4440 -18332 -4376 -17508
rect -3028 -18332 -2964 -17508
rect -1616 -18332 -1552 -17508
rect -204 -18332 -140 -17508
rect 1208 -18332 1272 -17508
rect 2620 -18332 2684 -17508
rect 4032 -18332 4096 -17508
rect 5444 -18332 5508 -17508
rect 6856 -18332 6920 -17508
rect 8268 -18332 8332 -17508
rect 9680 -18332 9744 -17508
rect 11092 -18332 11156 -17508
rect 12504 -18332 12568 -17508
rect 13916 -18332 13980 -17508
rect 15328 -18332 15392 -17508
rect 16740 -18332 16804 -17508
rect 18152 -18332 18216 -17508
rect 19564 -18332 19628 -17508
rect 20976 -18332 21040 -17508
rect 22388 -18332 22452 -17508
rect 23800 -18332 23864 -17508
<< mimcap >>
rect -23844 18280 -23044 18320
rect -23844 17560 -23804 18280
rect -23084 17560 -23044 18280
rect -23844 17520 -23044 17560
rect -22432 18280 -21632 18320
rect -22432 17560 -22392 18280
rect -21672 17560 -21632 18280
rect -22432 17520 -21632 17560
rect -21020 18280 -20220 18320
rect -21020 17560 -20980 18280
rect -20260 17560 -20220 18280
rect -21020 17520 -20220 17560
rect -19608 18280 -18808 18320
rect -19608 17560 -19568 18280
rect -18848 17560 -18808 18280
rect -19608 17520 -18808 17560
rect -18196 18280 -17396 18320
rect -18196 17560 -18156 18280
rect -17436 17560 -17396 18280
rect -18196 17520 -17396 17560
rect -16784 18280 -15984 18320
rect -16784 17560 -16744 18280
rect -16024 17560 -15984 18280
rect -16784 17520 -15984 17560
rect -15372 18280 -14572 18320
rect -15372 17560 -15332 18280
rect -14612 17560 -14572 18280
rect -15372 17520 -14572 17560
rect -13960 18280 -13160 18320
rect -13960 17560 -13920 18280
rect -13200 17560 -13160 18280
rect -13960 17520 -13160 17560
rect -12548 18280 -11748 18320
rect -12548 17560 -12508 18280
rect -11788 17560 -11748 18280
rect -12548 17520 -11748 17560
rect -11136 18280 -10336 18320
rect -11136 17560 -11096 18280
rect -10376 17560 -10336 18280
rect -11136 17520 -10336 17560
rect -9724 18280 -8924 18320
rect -9724 17560 -9684 18280
rect -8964 17560 -8924 18280
rect -9724 17520 -8924 17560
rect -8312 18280 -7512 18320
rect -8312 17560 -8272 18280
rect -7552 17560 -7512 18280
rect -8312 17520 -7512 17560
rect -6900 18280 -6100 18320
rect -6900 17560 -6860 18280
rect -6140 17560 -6100 18280
rect -6900 17520 -6100 17560
rect -5488 18280 -4688 18320
rect -5488 17560 -5448 18280
rect -4728 17560 -4688 18280
rect -5488 17520 -4688 17560
rect -4076 18280 -3276 18320
rect -4076 17560 -4036 18280
rect -3316 17560 -3276 18280
rect -4076 17520 -3276 17560
rect -2664 18280 -1864 18320
rect -2664 17560 -2624 18280
rect -1904 17560 -1864 18280
rect -2664 17520 -1864 17560
rect -1252 18280 -452 18320
rect -1252 17560 -1212 18280
rect -492 17560 -452 18280
rect -1252 17520 -452 17560
rect 160 18280 960 18320
rect 160 17560 200 18280
rect 920 17560 960 18280
rect 160 17520 960 17560
rect 1572 18280 2372 18320
rect 1572 17560 1612 18280
rect 2332 17560 2372 18280
rect 1572 17520 2372 17560
rect 2984 18280 3784 18320
rect 2984 17560 3024 18280
rect 3744 17560 3784 18280
rect 2984 17520 3784 17560
rect 4396 18280 5196 18320
rect 4396 17560 4436 18280
rect 5156 17560 5196 18280
rect 4396 17520 5196 17560
rect 5808 18280 6608 18320
rect 5808 17560 5848 18280
rect 6568 17560 6608 18280
rect 5808 17520 6608 17560
rect 7220 18280 8020 18320
rect 7220 17560 7260 18280
rect 7980 17560 8020 18280
rect 7220 17520 8020 17560
rect 8632 18280 9432 18320
rect 8632 17560 8672 18280
rect 9392 17560 9432 18280
rect 8632 17520 9432 17560
rect 10044 18280 10844 18320
rect 10044 17560 10084 18280
rect 10804 17560 10844 18280
rect 10044 17520 10844 17560
rect 11456 18280 12256 18320
rect 11456 17560 11496 18280
rect 12216 17560 12256 18280
rect 11456 17520 12256 17560
rect 12868 18280 13668 18320
rect 12868 17560 12908 18280
rect 13628 17560 13668 18280
rect 12868 17520 13668 17560
rect 14280 18280 15080 18320
rect 14280 17560 14320 18280
rect 15040 17560 15080 18280
rect 14280 17520 15080 17560
rect 15692 18280 16492 18320
rect 15692 17560 15732 18280
rect 16452 17560 16492 18280
rect 15692 17520 16492 17560
rect 17104 18280 17904 18320
rect 17104 17560 17144 18280
rect 17864 17560 17904 18280
rect 17104 17520 17904 17560
rect 18516 18280 19316 18320
rect 18516 17560 18556 18280
rect 19276 17560 19316 18280
rect 18516 17520 19316 17560
rect 19928 18280 20728 18320
rect 19928 17560 19968 18280
rect 20688 17560 20728 18280
rect 19928 17520 20728 17560
rect 21340 18280 22140 18320
rect 21340 17560 21380 18280
rect 22100 17560 22140 18280
rect 21340 17520 22140 17560
rect 22752 18280 23552 18320
rect 22752 17560 22792 18280
rect 23512 17560 23552 18280
rect 22752 17520 23552 17560
rect -23844 17160 -23044 17200
rect -23844 16440 -23804 17160
rect -23084 16440 -23044 17160
rect -23844 16400 -23044 16440
rect -22432 17160 -21632 17200
rect -22432 16440 -22392 17160
rect -21672 16440 -21632 17160
rect -22432 16400 -21632 16440
rect -21020 17160 -20220 17200
rect -21020 16440 -20980 17160
rect -20260 16440 -20220 17160
rect -21020 16400 -20220 16440
rect -19608 17160 -18808 17200
rect -19608 16440 -19568 17160
rect -18848 16440 -18808 17160
rect -19608 16400 -18808 16440
rect -18196 17160 -17396 17200
rect -18196 16440 -18156 17160
rect -17436 16440 -17396 17160
rect -18196 16400 -17396 16440
rect -16784 17160 -15984 17200
rect -16784 16440 -16744 17160
rect -16024 16440 -15984 17160
rect -16784 16400 -15984 16440
rect -15372 17160 -14572 17200
rect -15372 16440 -15332 17160
rect -14612 16440 -14572 17160
rect -15372 16400 -14572 16440
rect -13960 17160 -13160 17200
rect -13960 16440 -13920 17160
rect -13200 16440 -13160 17160
rect -13960 16400 -13160 16440
rect -12548 17160 -11748 17200
rect -12548 16440 -12508 17160
rect -11788 16440 -11748 17160
rect -12548 16400 -11748 16440
rect -11136 17160 -10336 17200
rect -11136 16440 -11096 17160
rect -10376 16440 -10336 17160
rect -11136 16400 -10336 16440
rect -9724 17160 -8924 17200
rect -9724 16440 -9684 17160
rect -8964 16440 -8924 17160
rect -9724 16400 -8924 16440
rect -8312 17160 -7512 17200
rect -8312 16440 -8272 17160
rect -7552 16440 -7512 17160
rect -8312 16400 -7512 16440
rect -6900 17160 -6100 17200
rect -6900 16440 -6860 17160
rect -6140 16440 -6100 17160
rect -6900 16400 -6100 16440
rect -5488 17160 -4688 17200
rect -5488 16440 -5448 17160
rect -4728 16440 -4688 17160
rect -5488 16400 -4688 16440
rect -4076 17160 -3276 17200
rect -4076 16440 -4036 17160
rect -3316 16440 -3276 17160
rect -4076 16400 -3276 16440
rect -2664 17160 -1864 17200
rect -2664 16440 -2624 17160
rect -1904 16440 -1864 17160
rect -2664 16400 -1864 16440
rect -1252 17160 -452 17200
rect -1252 16440 -1212 17160
rect -492 16440 -452 17160
rect -1252 16400 -452 16440
rect 160 17160 960 17200
rect 160 16440 200 17160
rect 920 16440 960 17160
rect 160 16400 960 16440
rect 1572 17160 2372 17200
rect 1572 16440 1612 17160
rect 2332 16440 2372 17160
rect 1572 16400 2372 16440
rect 2984 17160 3784 17200
rect 2984 16440 3024 17160
rect 3744 16440 3784 17160
rect 2984 16400 3784 16440
rect 4396 17160 5196 17200
rect 4396 16440 4436 17160
rect 5156 16440 5196 17160
rect 4396 16400 5196 16440
rect 5808 17160 6608 17200
rect 5808 16440 5848 17160
rect 6568 16440 6608 17160
rect 5808 16400 6608 16440
rect 7220 17160 8020 17200
rect 7220 16440 7260 17160
rect 7980 16440 8020 17160
rect 7220 16400 8020 16440
rect 8632 17160 9432 17200
rect 8632 16440 8672 17160
rect 9392 16440 9432 17160
rect 8632 16400 9432 16440
rect 10044 17160 10844 17200
rect 10044 16440 10084 17160
rect 10804 16440 10844 17160
rect 10044 16400 10844 16440
rect 11456 17160 12256 17200
rect 11456 16440 11496 17160
rect 12216 16440 12256 17160
rect 11456 16400 12256 16440
rect 12868 17160 13668 17200
rect 12868 16440 12908 17160
rect 13628 16440 13668 17160
rect 12868 16400 13668 16440
rect 14280 17160 15080 17200
rect 14280 16440 14320 17160
rect 15040 16440 15080 17160
rect 14280 16400 15080 16440
rect 15692 17160 16492 17200
rect 15692 16440 15732 17160
rect 16452 16440 16492 17160
rect 15692 16400 16492 16440
rect 17104 17160 17904 17200
rect 17104 16440 17144 17160
rect 17864 16440 17904 17160
rect 17104 16400 17904 16440
rect 18516 17160 19316 17200
rect 18516 16440 18556 17160
rect 19276 16440 19316 17160
rect 18516 16400 19316 16440
rect 19928 17160 20728 17200
rect 19928 16440 19968 17160
rect 20688 16440 20728 17160
rect 19928 16400 20728 16440
rect 21340 17160 22140 17200
rect 21340 16440 21380 17160
rect 22100 16440 22140 17160
rect 21340 16400 22140 16440
rect 22752 17160 23552 17200
rect 22752 16440 22792 17160
rect 23512 16440 23552 17160
rect 22752 16400 23552 16440
rect -23844 16040 -23044 16080
rect -23844 15320 -23804 16040
rect -23084 15320 -23044 16040
rect -23844 15280 -23044 15320
rect -22432 16040 -21632 16080
rect -22432 15320 -22392 16040
rect -21672 15320 -21632 16040
rect -22432 15280 -21632 15320
rect -21020 16040 -20220 16080
rect -21020 15320 -20980 16040
rect -20260 15320 -20220 16040
rect -21020 15280 -20220 15320
rect -19608 16040 -18808 16080
rect -19608 15320 -19568 16040
rect -18848 15320 -18808 16040
rect -19608 15280 -18808 15320
rect -18196 16040 -17396 16080
rect -18196 15320 -18156 16040
rect -17436 15320 -17396 16040
rect -18196 15280 -17396 15320
rect -16784 16040 -15984 16080
rect -16784 15320 -16744 16040
rect -16024 15320 -15984 16040
rect -16784 15280 -15984 15320
rect -15372 16040 -14572 16080
rect -15372 15320 -15332 16040
rect -14612 15320 -14572 16040
rect -15372 15280 -14572 15320
rect -13960 16040 -13160 16080
rect -13960 15320 -13920 16040
rect -13200 15320 -13160 16040
rect -13960 15280 -13160 15320
rect -12548 16040 -11748 16080
rect -12548 15320 -12508 16040
rect -11788 15320 -11748 16040
rect -12548 15280 -11748 15320
rect -11136 16040 -10336 16080
rect -11136 15320 -11096 16040
rect -10376 15320 -10336 16040
rect -11136 15280 -10336 15320
rect -9724 16040 -8924 16080
rect -9724 15320 -9684 16040
rect -8964 15320 -8924 16040
rect -9724 15280 -8924 15320
rect -8312 16040 -7512 16080
rect -8312 15320 -8272 16040
rect -7552 15320 -7512 16040
rect -8312 15280 -7512 15320
rect -6900 16040 -6100 16080
rect -6900 15320 -6860 16040
rect -6140 15320 -6100 16040
rect -6900 15280 -6100 15320
rect -5488 16040 -4688 16080
rect -5488 15320 -5448 16040
rect -4728 15320 -4688 16040
rect -5488 15280 -4688 15320
rect -4076 16040 -3276 16080
rect -4076 15320 -4036 16040
rect -3316 15320 -3276 16040
rect -4076 15280 -3276 15320
rect -2664 16040 -1864 16080
rect -2664 15320 -2624 16040
rect -1904 15320 -1864 16040
rect -2664 15280 -1864 15320
rect -1252 16040 -452 16080
rect -1252 15320 -1212 16040
rect -492 15320 -452 16040
rect -1252 15280 -452 15320
rect 160 16040 960 16080
rect 160 15320 200 16040
rect 920 15320 960 16040
rect 160 15280 960 15320
rect 1572 16040 2372 16080
rect 1572 15320 1612 16040
rect 2332 15320 2372 16040
rect 1572 15280 2372 15320
rect 2984 16040 3784 16080
rect 2984 15320 3024 16040
rect 3744 15320 3784 16040
rect 2984 15280 3784 15320
rect 4396 16040 5196 16080
rect 4396 15320 4436 16040
rect 5156 15320 5196 16040
rect 4396 15280 5196 15320
rect 5808 16040 6608 16080
rect 5808 15320 5848 16040
rect 6568 15320 6608 16040
rect 5808 15280 6608 15320
rect 7220 16040 8020 16080
rect 7220 15320 7260 16040
rect 7980 15320 8020 16040
rect 7220 15280 8020 15320
rect 8632 16040 9432 16080
rect 8632 15320 8672 16040
rect 9392 15320 9432 16040
rect 8632 15280 9432 15320
rect 10044 16040 10844 16080
rect 10044 15320 10084 16040
rect 10804 15320 10844 16040
rect 10044 15280 10844 15320
rect 11456 16040 12256 16080
rect 11456 15320 11496 16040
rect 12216 15320 12256 16040
rect 11456 15280 12256 15320
rect 12868 16040 13668 16080
rect 12868 15320 12908 16040
rect 13628 15320 13668 16040
rect 12868 15280 13668 15320
rect 14280 16040 15080 16080
rect 14280 15320 14320 16040
rect 15040 15320 15080 16040
rect 14280 15280 15080 15320
rect 15692 16040 16492 16080
rect 15692 15320 15732 16040
rect 16452 15320 16492 16040
rect 15692 15280 16492 15320
rect 17104 16040 17904 16080
rect 17104 15320 17144 16040
rect 17864 15320 17904 16040
rect 17104 15280 17904 15320
rect 18516 16040 19316 16080
rect 18516 15320 18556 16040
rect 19276 15320 19316 16040
rect 18516 15280 19316 15320
rect 19928 16040 20728 16080
rect 19928 15320 19968 16040
rect 20688 15320 20728 16040
rect 19928 15280 20728 15320
rect 21340 16040 22140 16080
rect 21340 15320 21380 16040
rect 22100 15320 22140 16040
rect 21340 15280 22140 15320
rect 22752 16040 23552 16080
rect 22752 15320 22792 16040
rect 23512 15320 23552 16040
rect 22752 15280 23552 15320
rect -23844 14920 -23044 14960
rect -23844 14200 -23804 14920
rect -23084 14200 -23044 14920
rect -23844 14160 -23044 14200
rect -22432 14920 -21632 14960
rect -22432 14200 -22392 14920
rect -21672 14200 -21632 14920
rect -22432 14160 -21632 14200
rect -21020 14920 -20220 14960
rect -21020 14200 -20980 14920
rect -20260 14200 -20220 14920
rect -21020 14160 -20220 14200
rect -19608 14920 -18808 14960
rect -19608 14200 -19568 14920
rect -18848 14200 -18808 14920
rect -19608 14160 -18808 14200
rect -18196 14920 -17396 14960
rect -18196 14200 -18156 14920
rect -17436 14200 -17396 14920
rect -18196 14160 -17396 14200
rect -16784 14920 -15984 14960
rect -16784 14200 -16744 14920
rect -16024 14200 -15984 14920
rect -16784 14160 -15984 14200
rect -15372 14920 -14572 14960
rect -15372 14200 -15332 14920
rect -14612 14200 -14572 14920
rect -15372 14160 -14572 14200
rect -13960 14920 -13160 14960
rect -13960 14200 -13920 14920
rect -13200 14200 -13160 14920
rect -13960 14160 -13160 14200
rect -12548 14920 -11748 14960
rect -12548 14200 -12508 14920
rect -11788 14200 -11748 14920
rect -12548 14160 -11748 14200
rect -11136 14920 -10336 14960
rect -11136 14200 -11096 14920
rect -10376 14200 -10336 14920
rect -11136 14160 -10336 14200
rect -9724 14920 -8924 14960
rect -9724 14200 -9684 14920
rect -8964 14200 -8924 14920
rect -9724 14160 -8924 14200
rect -8312 14920 -7512 14960
rect -8312 14200 -8272 14920
rect -7552 14200 -7512 14920
rect -8312 14160 -7512 14200
rect -6900 14920 -6100 14960
rect -6900 14200 -6860 14920
rect -6140 14200 -6100 14920
rect -6900 14160 -6100 14200
rect -5488 14920 -4688 14960
rect -5488 14200 -5448 14920
rect -4728 14200 -4688 14920
rect -5488 14160 -4688 14200
rect -4076 14920 -3276 14960
rect -4076 14200 -4036 14920
rect -3316 14200 -3276 14920
rect -4076 14160 -3276 14200
rect -2664 14920 -1864 14960
rect -2664 14200 -2624 14920
rect -1904 14200 -1864 14920
rect -2664 14160 -1864 14200
rect -1252 14920 -452 14960
rect -1252 14200 -1212 14920
rect -492 14200 -452 14920
rect -1252 14160 -452 14200
rect 160 14920 960 14960
rect 160 14200 200 14920
rect 920 14200 960 14920
rect 160 14160 960 14200
rect 1572 14920 2372 14960
rect 1572 14200 1612 14920
rect 2332 14200 2372 14920
rect 1572 14160 2372 14200
rect 2984 14920 3784 14960
rect 2984 14200 3024 14920
rect 3744 14200 3784 14920
rect 2984 14160 3784 14200
rect 4396 14920 5196 14960
rect 4396 14200 4436 14920
rect 5156 14200 5196 14920
rect 4396 14160 5196 14200
rect 5808 14920 6608 14960
rect 5808 14200 5848 14920
rect 6568 14200 6608 14920
rect 5808 14160 6608 14200
rect 7220 14920 8020 14960
rect 7220 14200 7260 14920
rect 7980 14200 8020 14920
rect 7220 14160 8020 14200
rect 8632 14920 9432 14960
rect 8632 14200 8672 14920
rect 9392 14200 9432 14920
rect 8632 14160 9432 14200
rect 10044 14920 10844 14960
rect 10044 14200 10084 14920
rect 10804 14200 10844 14920
rect 10044 14160 10844 14200
rect 11456 14920 12256 14960
rect 11456 14200 11496 14920
rect 12216 14200 12256 14920
rect 11456 14160 12256 14200
rect 12868 14920 13668 14960
rect 12868 14200 12908 14920
rect 13628 14200 13668 14920
rect 12868 14160 13668 14200
rect 14280 14920 15080 14960
rect 14280 14200 14320 14920
rect 15040 14200 15080 14920
rect 14280 14160 15080 14200
rect 15692 14920 16492 14960
rect 15692 14200 15732 14920
rect 16452 14200 16492 14920
rect 15692 14160 16492 14200
rect 17104 14920 17904 14960
rect 17104 14200 17144 14920
rect 17864 14200 17904 14920
rect 17104 14160 17904 14200
rect 18516 14920 19316 14960
rect 18516 14200 18556 14920
rect 19276 14200 19316 14920
rect 18516 14160 19316 14200
rect 19928 14920 20728 14960
rect 19928 14200 19968 14920
rect 20688 14200 20728 14920
rect 19928 14160 20728 14200
rect 21340 14920 22140 14960
rect 21340 14200 21380 14920
rect 22100 14200 22140 14920
rect 21340 14160 22140 14200
rect 22752 14920 23552 14960
rect 22752 14200 22792 14920
rect 23512 14200 23552 14920
rect 22752 14160 23552 14200
rect -23844 13800 -23044 13840
rect -23844 13080 -23804 13800
rect -23084 13080 -23044 13800
rect -23844 13040 -23044 13080
rect -22432 13800 -21632 13840
rect -22432 13080 -22392 13800
rect -21672 13080 -21632 13800
rect -22432 13040 -21632 13080
rect -21020 13800 -20220 13840
rect -21020 13080 -20980 13800
rect -20260 13080 -20220 13800
rect -21020 13040 -20220 13080
rect -19608 13800 -18808 13840
rect -19608 13080 -19568 13800
rect -18848 13080 -18808 13800
rect -19608 13040 -18808 13080
rect -18196 13800 -17396 13840
rect -18196 13080 -18156 13800
rect -17436 13080 -17396 13800
rect -18196 13040 -17396 13080
rect -16784 13800 -15984 13840
rect -16784 13080 -16744 13800
rect -16024 13080 -15984 13800
rect -16784 13040 -15984 13080
rect -15372 13800 -14572 13840
rect -15372 13080 -15332 13800
rect -14612 13080 -14572 13800
rect -15372 13040 -14572 13080
rect -13960 13800 -13160 13840
rect -13960 13080 -13920 13800
rect -13200 13080 -13160 13800
rect -13960 13040 -13160 13080
rect -12548 13800 -11748 13840
rect -12548 13080 -12508 13800
rect -11788 13080 -11748 13800
rect -12548 13040 -11748 13080
rect -11136 13800 -10336 13840
rect -11136 13080 -11096 13800
rect -10376 13080 -10336 13800
rect -11136 13040 -10336 13080
rect -9724 13800 -8924 13840
rect -9724 13080 -9684 13800
rect -8964 13080 -8924 13800
rect -9724 13040 -8924 13080
rect -8312 13800 -7512 13840
rect -8312 13080 -8272 13800
rect -7552 13080 -7512 13800
rect -8312 13040 -7512 13080
rect -6900 13800 -6100 13840
rect -6900 13080 -6860 13800
rect -6140 13080 -6100 13800
rect -6900 13040 -6100 13080
rect -5488 13800 -4688 13840
rect -5488 13080 -5448 13800
rect -4728 13080 -4688 13800
rect -5488 13040 -4688 13080
rect -4076 13800 -3276 13840
rect -4076 13080 -4036 13800
rect -3316 13080 -3276 13800
rect -4076 13040 -3276 13080
rect -2664 13800 -1864 13840
rect -2664 13080 -2624 13800
rect -1904 13080 -1864 13800
rect -2664 13040 -1864 13080
rect -1252 13800 -452 13840
rect -1252 13080 -1212 13800
rect -492 13080 -452 13800
rect -1252 13040 -452 13080
rect 160 13800 960 13840
rect 160 13080 200 13800
rect 920 13080 960 13800
rect 160 13040 960 13080
rect 1572 13800 2372 13840
rect 1572 13080 1612 13800
rect 2332 13080 2372 13800
rect 1572 13040 2372 13080
rect 2984 13800 3784 13840
rect 2984 13080 3024 13800
rect 3744 13080 3784 13800
rect 2984 13040 3784 13080
rect 4396 13800 5196 13840
rect 4396 13080 4436 13800
rect 5156 13080 5196 13800
rect 4396 13040 5196 13080
rect 5808 13800 6608 13840
rect 5808 13080 5848 13800
rect 6568 13080 6608 13800
rect 5808 13040 6608 13080
rect 7220 13800 8020 13840
rect 7220 13080 7260 13800
rect 7980 13080 8020 13800
rect 7220 13040 8020 13080
rect 8632 13800 9432 13840
rect 8632 13080 8672 13800
rect 9392 13080 9432 13800
rect 8632 13040 9432 13080
rect 10044 13800 10844 13840
rect 10044 13080 10084 13800
rect 10804 13080 10844 13800
rect 10044 13040 10844 13080
rect 11456 13800 12256 13840
rect 11456 13080 11496 13800
rect 12216 13080 12256 13800
rect 11456 13040 12256 13080
rect 12868 13800 13668 13840
rect 12868 13080 12908 13800
rect 13628 13080 13668 13800
rect 12868 13040 13668 13080
rect 14280 13800 15080 13840
rect 14280 13080 14320 13800
rect 15040 13080 15080 13800
rect 14280 13040 15080 13080
rect 15692 13800 16492 13840
rect 15692 13080 15732 13800
rect 16452 13080 16492 13800
rect 15692 13040 16492 13080
rect 17104 13800 17904 13840
rect 17104 13080 17144 13800
rect 17864 13080 17904 13800
rect 17104 13040 17904 13080
rect 18516 13800 19316 13840
rect 18516 13080 18556 13800
rect 19276 13080 19316 13800
rect 18516 13040 19316 13080
rect 19928 13800 20728 13840
rect 19928 13080 19968 13800
rect 20688 13080 20728 13800
rect 19928 13040 20728 13080
rect 21340 13800 22140 13840
rect 21340 13080 21380 13800
rect 22100 13080 22140 13800
rect 21340 13040 22140 13080
rect 22752 13800 23552 13840
rect 22752 13080 22792 13800
rect 23512 13080 23552 13800
rect 22752 13040 23552 13080
rect -23844 12680 -23044 12720
rect -23844 11960 -23804 12680
rect -23084 11960 -23044 12680
rect -23844 11920 -23044 11960
rect -22432 12680 -21632 12720
rect -22432 11960 -22392 12680
rect -21672 11960 -21632 12680
rect -22432 11920 -21632 11960
rect -21020 12680 -20220 12720
rect -21020 11960 -20980 12680
rect -20260 11960 -20220 12680
rect -21020 11920 -20220 11960
rect -19608 12680 -18808 12720
rect -19608 11960 -19568 12680
rect -18848 11960 -18808 12680
rect -19608 11920 -18808 11960
rect -18196 12680 -17396 12720
rect -18196 11960 -18156 12680
rect -17436 11960 -17396 12680
rect -18196 11920 -17396 11960
rect -16784 12680 -15984 12720
rect -16784 11960 -16744 12680
rect -16024 11960 -15984 12680
rect -16784 11920 -15984 11960
rect -15372 12680 -14572 12720
rect -15372 11960 -15332 12680
rect -14612 11960 -14572 12680
rect -15372 11920 -14572 11960
rect -13960 12680 -13160 12720
rect -13960 11960 -13920 12680
rect -13200 11960 -13160 12680
rect -13960 11920 -13160 11960
rect -12548 12680 -11748 12720
rect -12548 11960 -12508 12680
rect -11788 11960 -11748 12680
rect -12548 11920 -11748 11960
rect -11136 12680 -10336 12720
rect -11136 11960 -11096 12680
rect -10376 11960 -10336 12680
rect -11136 11920 -10336 11960
rect -9724 12680 -8924 12720
rect -9724 11960 -9684 12680
rect -8964 11960 -8924 12680
rect -9724 11920 -8924 11960
rect -8312 12680 -7512 12720
rect -8312 11960 -8272 12680
rect -7552 11960 -7512 12680
rect -8312 11920 -7512 11960
rect -6900 12680 -6100 12720
rect -6900 11960 -6860 12680
rect -6140 11960 -6100 12680
rect -6900 11920 -6100 11960
rect -5488 12680 -4688 12720
rect -5488 11960 -5448 12680
rect -4728 11960 -4688 12680
rect -5488 11920 -4688 11960
rect -4076 12680 -3276 12720
rect -4076 11960 -4036 12680
rect -3316 11960 -3276 12680
rect -4076 11920 -3276 11960
rect -2664 12680 -1864 12720
rect -2664 11960 -2624 12680
rect -1904 11960 -1864 12680
rect -2664 11920 -1864 11960
rect -1252 12680 -452 12720
rect -1252 11960 -1212 12680
rect -492 11960 -452 12680
rect -1252 11920 -452 11960
rect 160 12680 960 12720
rect 160 11960 200 12680
rect 920 11960 960 12680
rect 160 11920 960 11960
rect 1572 12680 2372 12720
rect 1572 11960 1612 12680
rect 2332 11960 2372 12680
rect 1572 11920 2372 11960
rect 2984 12680 3784 12720
rect 2984 11960 3024 12680
rect 3744 11960 3784 12680
rect 2984 11920 3784 11960
rect 4396 12680 5196 12720
rect 4396 11960 4436 12680
rect 5156 11960 5196 12680
rect 4396 11920 5196 11960
rect 5808 12680 6608 12720
rect 5808 11960 5848 12680
rect 6568 11960 6608 12680
rect 5808 11920 6608 11960
rect 7220 12680 8020 12720
rect 7220 11960 7260 12680
rect 7980 11960 8020 12680
rect 7220 11920 8020 11960
rect 8632 12680 9432 12720
rect 8632 11960 8672 12680
rect 9392 11960 9432 12680
rect 8632 11920 9432 11960
rect 10044 12680 10844 12720
rect 10044 11960 10084 12680
rect 10804 11960 10844 12680
rect 10044 11920 10844 11960
rect 11456 12680 12256 12720
rect 11456 11960 11496 12680
rect 12216 11960 12256 12680
rect 11456 11920 12256 11960
rect 12868 12680 13668 12720
rect 12868 11960 12908 12680
rect 13628 11960 13668 12680
rect 12868 11920 13668 11960
rect 14280 12680 15080 12720
rect 14280 11960 14320 12680
rect 15040 11960 15080 12680
rect 14280 11920 15080 11960
rect 15692 12680 16492 12720
rect 15692 11960 15732 12680
rect 16452 11960 16492 12680
rect 15692 11920 16492 11960
rect 17104 12680 17904 12720
rect 17104 11960 17144 12680
rect 17864 11960 17904 12680
rect 17104 11920 17904 11960
rect 18516 12680 19316 12720
rect 18516 11960 18556 12680
rect 19276 11960 19316 12680
rect 18516 11920 19316 11960
rect 19928 12680 20728 12720
rect 19928 11960 19968 12680
rect 20688 11960 20728 12680
rect 19928 11920 20728 11960
rect 21340 12680 22140 12720
rect 21340 11960 21380 12680
rect 22100 11960 22140 12680
rect 21340 11920 22140 11960
rect 22752 12680 23552 12720
rect 22752 11960 22792 12680
rect 23512 11960 23552 12680
rect 22752 11920 23552 11960
rect -23844 11560 -23044 11600
rect -23844 10840 -23804 11560
rect -23084 10840 -23044 11560
rect -23844 10800 -23044 10840
rect -22432 11560 -21632 11600
rect -22432 10840 -22392 11560
rect -21672 10840 -21632 11560
rect -22432 10800 -21632 10840
rect -21020 11560 -20220 11600
rect -21020 10840 -20980 11560
rect -20260 10840 -20220 11560
rect -21020 10800 -20220 10840
rect -19608 11560 -18808 11600
rect -19608 10840 -19568 11560
rect -18848 10840 -18808 11560
rect -19608 10800 -18808 10840
rect -18196 11560 -17396 11600
rect -18196 10840 -18156 11560
rect -17436 10840 -17396 11560
rect -18196 10800 -17396 10840
rect -16784 11560 -15984 11600
rect -16784 10840 -16744 11560
rect -16024 10840 -15984 11560
rect -16784 10800 -15984 10840
rect -15372 11560 -14572 11600
rect -15372 10840 -15332 11560
rect -14612 10840 -14572 11560
rect -15372 10800 -14572 10840
rect -13960 11560 -13160 11600
rect -13960 10840 -13920 11560
rect -13200 10840 -13160 11560
rect -13960 10800 -13160 10840
rect -12548 11560 -11748 11600
rect -12548 10840 -12508 11560
rect -11788 10840 -11748 11560
rect -12548 10800 -11748 10840
rect -11136 11560 -10336 11600
rect -11136 10840 -11096 11560
rect -10376 10840 -10336 11560
rect -11136 10800 -10336 10840
rect -9724 11560 -8924 11600
rect -9724 10840 -9684 11560
rect -8964 10840 -8924 11560
rect -9724 10800 -8924 10840
rect -8312 11560 -7512 11600
rect -8312 10840 -8272 11560
rect -7552 10840 -7512 11560
rect -8312 10800 -7512 10840
rect -6900 11560 -6100 11600
rect -6900 10840 -6860 11560
rect -6140 10840 -6100 11560
rect -6900 10800 -6100 10840
rect -5488 11560 -4688 11600
rect -5488 10840 -5448 11560
rect -4728 10840 -4688 11560
rect -5488 10800 -4688 10840
rect -4076 11560 -3276 11600
rect -4076 10840 -4036 11560
rect -3316 10840 -3276 11560
rect -4076 10800 -3276 10840
rect -2664 11560 -1864 11600
rect -2664 10840 -2624 11560
rect -1904 10840 -1864 11560
rect -2664 10800 -1864 10840
rect -1252 11560 -452 11600
rect -1252 10840 -1212 11560
rect -492 10840 -452 11560
rect -1252 10800 -452 10840
rect 160 11560 960 11600
rect 160 10840 200 11560
rect 920 10840 960 11560
rect 160 10800 960 10840
rect 1572 11560 2372 11600
rect 1572 10840 1612 11560
rect 2332 10840 2372 11560
rect 1572 10800 2372 10840
rect 2984 11560 3784 11600
rect 2984 10840 3024 11560
rect 3744 10840 3784 11560
rect 2984 10800 3784 10840
rect 4396 11560 5196 11600
rect 4396 10840 4436 11560
rect 5156 10840 5196 11560
rect 4396 10800 5196 10840
rect 5808 11560 6608 11600
rect 5808 10840 5848 11560
rect 6568 10840 6608 11560
rect 5808 10800 6608 10840
rect 7220 11560 8020 11600
rect 7220 10840 7260 11560
rect 7980 10840 8020 11560
rect 7220 10800 8020 10840
rect 8632 11560 9432 11600
rect 8632 10840 8672 11560
rect 9392 10840 9432 11560
rect 8632 10800 9432 10840
rect 10044 11560 10844 11600
rect 10044 10840 10084 11560
rect 10804 10840 10844 11560
rect 10044 10800 10844 10840
rect 11456 11560 12256 11600
rect 11456 10840 11496 11560
rect 12216 10840 12256 11560
rect 11456 10800 12256 10840
rect 12868 11560 13668 11600
rect 12868 10840 12908 11560
rect 13628 10840 13668 11560
rect 12868 10800 13668 10840
rect 14280 11560 15080 11600
rect 14280 10840 14320 11560
rect 15040 10840 15080 11560
rect 14280 10800 15080 10840
rect 15692 11560 16492 11600
rect 15692 10840 15732 11560
rect 16452 10840 16492 11560
rect 15692 10800 16492 10840
rect 17104 11560 17904 11600
rect 17104 10840 17144 11560
rect 17864 10840 17904 11560
rect 17104 10800 17904 10840
rect 18516 11560 19316 11600
rect 18516 10840 18556 11560
rect 19276 10840 19316 11560
rect 18516 10800 19316 10840
rect 19928 11560 20728 11600
rect 19928 10840 19968 11560
rect 20688 10840 20728 11560
rect 19928 10800 20728 10840
rect 21340 11560 22140 11600
rect 21340 10840 21380 11560
rect 22100 10840 22140 11560
rect 21340 10800 22140 10840
rect 22752 11560 23552 11600
rect 22752 10840 22792 11560
rect 23512 10840 23552 11560
rect 22752 10800 23552 10840
rect -23844 10440 -23044 10480
rect -23844 9720 -23804 10440
rect -23084 9720 -23044 10440
rect -23844 9680 -23044 9720
rect -22432 10440 -21632 10480
rect -22432 9720 -22392 10440
rect -21672 9720 -21632 10440
rect -22432 9680 -21632 9720
rect -21020 10440 -20220 10480
rect -21020 9720 -20980 10440
rect -20260 9720 -20220 10440
rect -21020 9680 -20220 9720
rect -19608 10440 -18808 10480
rect -19608 9720 -19568 10440
rect -18848 9720 -18808 10440
rect -19608 9680 -18808 9720
rect -18196 10440 -17396 10480
rect -18196 9720 -18156 10440
rect -17436 9720 -17396 10440
rect -18196 9680 -17396 9720
rect -16784 10440 -15984 10480
rect -16784 9720 -16744 10440
rect -16024 9720 -15984 10440
rect -16784 9680 -15984 9720
rect -15372 10440 -14572 10480
rect -15372 9720 -15332 10440
rect -14612 9720 -14572 10440
rect -15372 9680 -14572 9720
rect -13960 10440 -13160 10480
rect -13960 9720 -13920 10440
rect -13200 9720 -13160 10440
rect -13960 9680 -13160 9720
rect -12548 10440 -11748 10480
rect -12548 9720 -12508 10440
rect -11788 9720 -11748 10440
rect -12548 9680 -11748 9720
rect -11136 10440 -10336 10480
rect -11136 9720 -11096 10440
rect -10376 9720 -10336 10440
rect -11136 9680 -10336 9720
rect -9724 10440 -8924 10480
rect -9724 9720 -9684 10440
rect -8964 9720 -8924 10440
rect -9724 9680 -8924 9720
rect -8312 10440 -7512 10480
rect -8312 9720 -8272 10440
rect -7552 9720 -7512 10440
rect -8312 9680 -7512 9720
rect -6900 10440 -6100 10480
rect -6900 9720 -6860 10440
rect -6140 9720 -6100 10440
rect -6900 9680 -6100 9720
rect -5488 10440 -4688 10480
rect -5488 9720 -5448 10440
rect -4728 9720 -4688 10440
rect -5488 9680 -4688 9720
rect -4076 10440 -3276 10480
rect -4076 9720 -4036 10440
rect -3316 9720 -3276 10440
rect -4076 9680 -3276 9720
rect -2664 10440 -1864 10480
rect -2664 9720 -2624 10440
rect -1904 9720 -1864 10440
rect -2664 9680 -1864 9720
rect -1252 10440 -452 10480
rect -1252 9720 -1212 10440
rect -492 9720 -452 10440
rect -1252 9680 -452 9720
rect 160 10440 960 10480
rect 160 9720 200 10440
rect 920 9720 960 10440
rect 160 9680 960 9720
rect 1572 10440 2372 10480
rect 1572 9720 1612 10440
rect 2332 9720 2372 10440
rect 1572 9680 2372 9720
rect 2984 10440 3784 10480
rect 2984 9720 3024 10440
rect 3744 9720 3784 10440
rect 2984 9680 3784 9720
rect 4396 10440 5196 10480
rect 4396 9720 4436 10440
rect 5156 9720 5196 10440
rect 4396 9680 5196 9720
rect 5808 10440 6608 10480
rect 5808 9720 5848 10440
rect 6568 9720 6608 10440
rect 5808 9680 6608 9720
rect 7220 10440 8020 10480
rect 7220 9720 7260 10440
rect 7980 9720 8020 10440
rect 7220 9680 8020 9720
rect 8632 10440 9432 10480
rect 8632 9720 8672 10440
rect 9392 9720 9432 10440
rect 8632 9680 9432 9720
rect 10044 10440 10844 10480
rect 10044 9720 10084 10440
rect 10804 9720 10844 10440
rect 10044 9680 10844 9720
rect 11456 10440 12256 10480
rect 11456 9720 11496 10440
rect 12216 9720 12256 10440
rect 11456 9680 12256 9720
rect 12868 10440 13668 10480
rect 12868 9720 12908 10440
rect 13628 9720 13668 10440
rect 12868 9680 13668 9720
rect 14280 10440 15080 10480
rect 14280 9720 14320 10440
rect 15040 9720 15080 10440
rect 14280 9680 15080 9720
rect 15692 10440 16492 10480
rect 15692 9720 15732 10440
rect 16452 9720 16492 10440
rect 15692 9680 16492 9720
rect 17104 10440 17904 10480
rect 17104 9720 17144 10440
rect 17864 9720 17904 10440
rect 17104 9680 17904 9720
rect 18516 10440 19316 10480
rect 18516 9720 18556 10440
rect 19276 9720 19316 10440
rect 18516 9680 19316 9720
rect 19928 10440 20728 10480
rect 19928 9720 19968 10440
rect 20688 9720 20728 10440
rect 19928 9680 20728 9720
rect 21340 10440 22140 10480
rect 21340 9720 21380 10440
rect 22100 9720 22140 10440
rect 21340 9680 22140 9720
rect 22752 10440 23552 10480
rect 22752 9720 22792 10440
rect 23512 9720 23552 10440
rect 22752 9680 23552 9720
rect -23844 9320 -23044 9360
rect -23844 8600 -23804 9320
rect -23084 8600 -23044 9320
rect -23844 8560 -23044 8600
rect -22432 9320 -21632 9360
rect -22432 8600 -22392 9320
rect -21672 8600 -21632 9320
rect -22432 8560 -21632 8600
rect -21020 9320 -20220 9360
rect -21020 8600 -20980 9320
rect -20260 8600 -20220 9320
rect -21020 8560 -20220 8600
rect -19608 9320 -18808 9360
rect -19608 8600 -19568 9320
rect -18848 8600 -18808 9320
rect -19608 8560 -18808 8600
rect -18196 9320 -17396 9360
rect -18196 8600 -18156 9320
rect -17436 8600 -17396 9320
rect -18196 8560 -17396 8600
rect -16784 9320 -15984 9360
rect -16784 8600 -16744 9320
rect -16024 8600 -15984 9320
rect -16784 8560 -15984 8600
rect -15372 9320 -14572 9360
rect -15372 8600 -15332 9320
rect -14612 8600 -14572 9320
rect -15372 8560 -14572 8600
rect -13960 9320 -13160 9360
rect -13960 8600 -13920 9320
rect -13200 8600 -13160 9320
rect -13960 8560 -13160 8600
rect -12548 9320 -11748 9360
rect -12548 8600 -12508 9320
rect -11788 8600 -11748 9320
rect -12548 8560 -11748 8600
rect -11136 9320 -10336 9360
rect -11136 8600 -11096 9320
rect -10376 8600 -10336 9320
rect -11136 8560 -10336 8600
rect -9724 9320 -8924 9360
rect -9724 8600 -9684 9320
rect -8964 8600 -8924 9320
rect -9724 8560 -8924 8600
rect -8312 9320 -7512 9360
rect -8312 8600 -8272 9320
rect -7552 8600 -7512 9320
rect -8312 8560 -7512 8600
rect -6900 9320 -6100 9360
rect -6900 8600 -6860 9320
rect -6140 8600 -6100 9320
rect -6900 8560 -6100 8600
rect -5488 9320 -4688 9360
rect -5488 8600 -5448 9320
rect -4728 8600 -4688 9320
rect -5488 8560 -4688 8600
rect -4076 9320 -3276 9360
rect -4076 8600 -4036 9320
rect -3316 8600 -3276 9320
rect -4076 8560 -3276 8600
rect -2664 9320 -1864 9360
rect -2664 8600 -2624 9320
rect -1904 8600 -1864 9320
rect -2664 8560 -1864 8600
rect -1252 9320 -452 9360
rect -1252 8600 -1212 9320
rect -492 8600 -452 9320
rect -1252 8560 -452 8600
rect 160 9320 960 9360
rect 160 8600 200 9320
rect 920 8600 960 9320
rect 160 8560 960 8600
rect 1572 9320 2372 9360
rect 1572 8600 1612 9320
rect 2332 8600 2372 9320
rect 1572 8560 2372 8600
rect 2984 9320 3784 9360
rect 2984 8600 3024 9320
rect 3744 8600 3784 9320
rect 2984 8560 3784 8600
rect 4396 9320 5196 9360
rect 4396 8600 4436 9320
rect 5156 8600 5196 9320
rect 4396 8560 5196 8600
rect 5808 9320 6608 9360
rect 5808 8600 5848 9320
rect 6568 8600 6608 9320
rect 5808 8560 6608 8600
rect 7220 9320 8020 9360
rect 7220 8600 7260 9320
rect 7980 8600 8020 9320
rect 7220 8560 8020 8600
rect 8632 9320 9432 9360
rect 8632 8600 8672 9320
rect 9392 8600 9432 9320
rect 8632 8560 9432 8600
rect 10044 9320 10844 9360
rect 10044 8600 10084 9320
rect 10804 8600 10844 9320
rect 10044 8560 10844 8600
rect 11456 9320 12256 9360
rect 11456 8600 11496 9320
rect 12216 8600 12256 9320
rect 11456 8560 12256 8600
rect 12868 9320 13668 9360
rect 12868 8600 12908 9320
rect 13628 8600 13668 9320
rect 12868 8560 13668 8600
rect 14280 9320 15080 9360
rect 14280 8600 14320 9320
rect 15040 8600 15080 9320
rect 14280 8560 15080 8600
rect 15692 9320 16492 9360
rect 15692 8600 15732 9320
rect 16452 8600 16492 9320
rect 15692 8560 16492 8600
rect 17104 9320 17904 9360
rect 17104 8600 17144 9320
rect 17864 8600 17904 9320
rect 17104 8560 17904 8600
rect 18516 9320 19316 9360
rect 18516 8600 18556 9320
rect 19276 8600 19316 9320
rect 18516 8560 19316 8600
rect 19928 9320 20728 9360
rect 19928 8600 19968 9320
rect 20688 8600 20728 9320
rect 19928 8560 20728 8600
rect 21340 9320 22140 9360
rect 21340 8600 21380 9320
rect 22100 8600 22140 9320
rect 21340 8560 22140 8600
rect 22752 9320 23552 9360
rect 22752 8600 22792 9320
rect 23512 8600 23552 9320
rect 22752 8560 23552 8600
rect -23844 8200 -23044 8240
rect -23844 7480 -23804 8200
rect -23084 7480 -23044 8200
rect -23844 7440 -23044 7480
rect -22432 8200 -21632 8240
rect -22432 7480 -22392 8200
rect -21672 7480 -21632 8200
rect -22432 7440 -21632 7480
rect -21020 8200 -20220 8240
rect -21020 7480 -20980 8200
rect -20260 7480 -20220 8200
rect -21020 7440 -20220 7480
rect -19608 8200 -18808 8240
rect -19608 7480 -19568 8200
rect -18848 7480 -18808 8200
rect -19608 7440 -18808 7480
rect -18196 8200 -17396 8240
rect -18196 7480 -18156 8200
rect -17436 7480 -17396 8200
rect -18196 7440 -17396 7480
rect -16784 8200 -15984 8240
rect -16784 7480 -16744 8200
rect -16024 7480 -15984 8200
rect -16784 7440 -15984 7480
rect -15372 8200 -14572 8240
rect -15372 7480 -15332 8200
rect -14612 7480 -14572 8200
rect -15372 7440 -14572 7480
rect -13960 8200 -13160 8240
rect -13960 7480 -13920 8200
rect -13200 7480 -13160 8200
rect -13960 7440 -13160 7480
rect -12548 8200 -11748 8240
rect -12548 7480 -12508 8200
rect -11788 7480 -11748 8200
rect -12548 7440 -11748 7480
rect -11136 8200 -10336 8240
rect -11136 7480 -11096 8200
rect -10376 7480 -10336 8200
rect -11136 7440 -10336 7480
rect -9724 8200 -8924 8240
rect -9724 7480 -9684 8200
rect -8964 7480 -8924 8200
rect -9724 7440 -8924 7480
rect -8312 8200 -7512 8240
rect -8312 7480 -8272 8200
rect -7552 7480 -7512 8200
rect -8312 7440 -7512 7480
rect -6900 8200 -6100 8240
rect -6900 7480 -6860 8200
rect -6140 7480 -6100 8200
rect -6900 7440 -6100 7480
rect -5488 8200 -4688 8240
rect -5488 7480 -5448 8200
rect -4728 7480 -4688 8200
rect -5488 7440 -4688 7480
rect -4076 8200 -3276 8240
rect -4076 7480 -4036 8200
rect -3316 7480 -3276 8200
rect -4076 7440 -3276 7480
rect -2664 8200 -1864 8240
rect -2664 7480 -2624 8200
rect -1904 7480 -1864 8200
rect -2664 7440 -1864 7480
rect -1252 8200 -452 8240
rect -1252 7480 -1212 8200
rect -492 7480 -452 8200
rect -1252 7440 -452 7480
rect 160 8200 960 8240
rect 160 7480 200 8200
rect 920 7480 960 8200
rect 160 7440 960 7480
rect 1572 8200 2372 8240
rect 1572 7480 1612 8200
rect 2332 7480 2372 8200
rect 1572 7440 2372 7480
rect 2984 8200 3784 8240
rect 2984 7480 3024 8200
rect 3744 7480 3784 8200
rect 2984 7440 3784 7480
rect 4396 8200 5196 8240
rect 4396 7480 4436 8200
rect 5156 7480 5196 8200
rect 4396 7440 5196 7480
rect 5808 8200 6608 8240
rect 5808 7480 5848 8200
rect 6568 7480 6608 8200
rect 5808 7440 6608 7480
rect 7220 8200 8020 8240
rect 7220 7480 7260 8200
rect 7980 7480 8020 8200
rect 7220 7440 8020 7480
rect 8632 8200 9432 8240
rect 8632 7480 8672 8200
rect 9392 7480 9432 8200
rect 8632 7440 9432 7480
rect 10044 8200 10844 8240
rect 10044 7480 10084 8200
rect 10804 7480 10844 8200
rect 10044 7440 10844 7480
rect 11456 8200 12256 8240
rect 11456 7480 11496 8200
rect 12216 7480 12256 8200
rect 11456 7440 12256 7480
rect 12868 8200 13668 8240
rect 12868 7480 12908 8200
rect 13628 7480 13668 8200
rect 12868 7440 13668 7480
rect 14280 8200 15080 8240
rect 14280 7480 14320 8200
rect 15040 7480 15080 8200
rect 14280 7440 15080 7480
rect 15692 8200 16492 8240
rect 15692 7480 15732 8200
rect 16452 7480 16492 8200
rect 15692 7440 16492 7480
rect 17104 8200 17904 8240
rect 17104 7480 17144 8200
rect 17864 7480 17904 8200
rect 17104 7440 17904 7480
rect 18516 8200 19316 8240
rect 18516 7480 18556 8200
rect 19276 7480 19316 8200
rect 18516 7440 19316 7480
rect 19928 8200 20728 8240
rect 19928 7480 19968 8200
rect 20688 7480 20728 8200
rect 19928 7440 20728 7480
rect 21340 8200 22140 8240
rect 21340 7480 21380 8200
rect 22100 7480 22140 8200
rect 21340 7440 22140 7480
rect 22752 8200 23552 8240
rect 22752 7480 22792 8200
rect 23512 7480 23552 8200
rect 22752 7440 23552 7480
rect -23844 7080 -23044 7120
rect -23844 6360 -23804 7080
rect -23084 6360 -23044 7080
rect -23844 6320 -23044 6360
rect -22432 7080 -21632 7120
rect -22432 6360 -22392 7080
rect -21672 6360 -21632 7080
rect -22432 6320 -21632 6360
rect -21020 7080 -20220 7120
rect -21020 6360 -20980 7080
rect -20260 6360 -20220 7080
rect -21020 6320 -20220 6360
rect -19608 7080 -18808 7120
rect -19608 6360 -19568 7080
rect -18848 6360 -18808 7080
rect -19608 6320 -18808 6360
rect -18196 7080 -17396 7120
rect -18196 6360 -18156 7080
rect -17436 6360 -17396 7080
rect -18196 6320 -17396 6360
rect -16784 7080 -15984 7120
rect -16784 6360 -16744 7080
rect -16024 6360 -15984 7080
rect -16784 6320 -15984 6360
rect -15372 7080 -14572 7120
rect -15372 6360 -15332 7080
rect -14612 6360 -14572 7080
rect -15372 6320 -14572 6360
rect -13960 7080 -13160 7120
rect -13960 6360 -13920 7080
rect -13200 6360 -13160 7080
rect -13960 6320 -13160 6360
rect -12548 7080 -11748 7120
rect -12548 6360 -12508 7080
rect -11788 6360 -11748 7080
rect -12548 6320 -11748 6360
rect -11136 7080 -10336 7120
rect -11136 6360 -11096 7080
rect -10376 6360 -10336 7080
rect -11136 6320 -10336 6360
rect -9724 7080 -8924 7120
rect -9724 6360 -9684 7080
rect -8964 6360 -8924 7080
rect -9724 6320 -8924 6360
rect -8312 7080 -7512 7120
rect -8312 6360 -8272 7080
rect -7552 6360 -7512 7080
rect -8312 6320 -7512 6360
rect -6900 7080 -6100 7120
rect -6900 6360 -6860 7080
rect -6140 6360 -6100 7080
rect -6900 6320 -6100 6360
rect -5488 7080 -4688 7120
rect -5488 6360 -5448 7080
rect -4728 6360 -4688 7080
rect -5488 6320 -4688 6360
rect -4076 7080 -3276 7120
rect -4076 6360 -4036 7080
rect -3316 6360 -3276 7080
rect -4076 6320 -3276 6360
rect -2664 7080 -1864 7120
rect -2664 6360 -2624 7080
rect -1904 6360 -1864 7080
rect -2664 6320 -1864 6360
rect -1252 7080 -452 7120
rect -1252 6360 -1212 7080
rect -492 6360 -452 7080
rect -1252 6320 -452 6360
rect 160 7080 960 7120
rect 160 6360 200 7080
rect 920 6360 960 7080
rect 160 6320 960 6360
rect 1572 7080 2372 7120
rect 1572 6360 1612 7080
rect 2332 6360 2372 7080
rect 1572 6320 2372 6360
rect 2984 7080 3784 7120
rect 2984 6360 3024 7080
rect 3744 6360 3784 7080
rect 2984 6320 3784 6360
rect 4396 7080 5196 7120
rect 4396 6360 4436 7080
rect 5156 6360 5196 7080
rect 4396 6320 5196 6360
rect 5808 7080 6608 7120
rect 5808 6360 5848 7080
rect 6568 6360 6608 7080
rect 5808 6320 6608 6360
rect 7220 7080 8020 7120
rect 7220 6360 7260 7080
rect 7980 6360 8020 7080
rect 7220 6320 8020 6360
rect 8632 7080 9432 7120
rect 8632 6360 8672 7080
rect 9392 6360 9432 7080
rect 8632 6320 9432 6360
rect 10044 7080 10844 7120
rect 10044 6360 10084 7080
rect 10804 6360 10844 7080
rect 10044 6320 10844 6360
rect 11456 7080 12256 7120
rect 11456 6360 11496 7080
rect 12216 6360 12256 7080
rect 11456 6320 12256 6360
rect 12868 7080 13668 7120
rect 12868 6360 12908 7080
rect 13628 6360 13668 7080
rect 12868 6320 13668 6360
rect 14280 7080 15080 7120
rect 14280 6360 14320 7080
rect 15040 6360 15080 7080
rect 14280 6320 15080 6360
rect 15692 7080 16492 7120
rect 15692 6360 15732 7080
rect 16452 6360 16492 7080
rect 15692 6320 16492 6360
rect 17104 7080 17904 7120
rect 17104 6360 17144 7080
rect 17864 6360 17904 7080
rect 17104 6320 17904 6360
rect 18516 7080 19316 7120
rect 18516 6360 18556 7080
rect 19276 6360 19316 7080
rect 18516 6320 19316 6360
rect 19928 7080 20728 7120
rect 19928 6360 19968 7080
rect 20688 6360 20728 7080
rect 19928 6320 20728 6360
rect 21340 7080 22140 7120
rect 21340 6360 21380 7080
rect 22100 6360 22140 7080
rect 21340 6320 22140 6360
rect 22752 7080 23552 7120
rect 22752 6360 22792 7080
rect 23512 6360 23552 7080
rect 22752 6320 23552 6360
rect -23844 5960 -23044 6000
rect -23844 5240 -23804 5960
rect -23084 5240 -23044 5960
rect -23844 5200 -23044 5240
rect -22432 5960 -21632 6000
rect -22432 5240 -22392 5960
rect -21672 5240 -21632 5960
rect -22432 5200 -21632 5240
rect -21020 5960 -20220 6000
rect -21020 5240 -20980 5960
rect -20260 5240 -20220 5960
rect -21020 5200 -20220 5240
rect -19608 5960 -18808 6000
rect -19608 5240 -19568 5960
rect -18848 5240 -18808 5960
rect -19608 5200 -18808 5240
rect -18196 5960 -17396 6000
rect -18196 5240 -18156 5960
rect -17436 5240 -17396 5960
rect -18196 5200 -17396 5240
rect -16784 5960 -15984 6000
rect -16784 5240 -16744 5960
rect -16024 5240 -15984 5960
rect -16784 5200 -15984 5240
rect -15372 5960 -14572 6000
rect -15372 5240 -15332 5960
rect -14612 5240 -14572 5960
rect -15372 5200 -14572 5240
rect -13960 5960 -13160 6000
rect -13960 5240 -13920 5960
rect -13200 5240 -13160 5960
rect -13960 5200 -13160 5240
rect -12548 5960 -11748 6000
rect -12548 5240 -12508 5960
rect -11788 5240 -11748 5960
rect -12548 5200 -11748 5240
rect -11136 5960 -10336 6000
rect -11136 5240 -11096 5960
rect -10376 5240 -10336 5960
rect -11136 5200 -10336 5240
rect -9724 5960 -8924 6000
rect -9724 5240 -9684 5960
rect -8964 5240 -8924 5960
rect -9724 5200 -8924 5240
rect -8312 5960 -7512 6000
rect -8312 5240 -8272 5960
rect -7552 5240 -7512 5960
rect -8312 5200 -7512 5240
rect -6900 5960 -6100 6000
rect -6900 5240 -6860 5960
rect -6140 5240 -6100 5960
rect -6900 5200 -6100 5240
rect -5488 5960 -4688 6000
rect -5488 5240 -5448 5960
rect -4728 5240 -4688 5960
rect -5488 5200 -4688 5240
rect -4076 5960 -3276 6000
rect -4076 5240 -4036 5960
rect -3316 5240 -3276 5960
rect -4076 5200 -3276 5240
rect -2664 5960 -1864 6000
rect -2664 5240 -2624 5960
rect -1904 5240 -1864 5960
rect -2664 5200 -1864 5240
rect -1252 5960 -452 6000
rect -1252 5240 -1212 5960
rect -492 5240 -452 5960
rect -1252 5200 -452 5240
rect 160 5960 960 6000
rect 160 5240 200 5960
rect 920 5240 960 5960
rect 160 5200 960 5240
rect 1572 5960 2372 6000
rect 1572 5240 1612 5960
rect 2332 5240 2372 5960
rect 1572 5200 2372 5240
rect 2984 5960 3784 6000
rect 2984 5240 3024 5960
rect 3744 5240 3784 5960
rect 2984 5200 3784 5240
rect 4396 5960 5196 6000
rect 4396 5240 4436 5960
rect 5156 5240 5196 5960
rect 4396 5200 5196 5240
rect 5808 5960 6608 6000
rect 5808 5240 5848 5960
rect 6568 5240 6608 5960
rect 5808 5200 6608 5240
rect 7220 5960 8020 6000
rect 7220 5240 7260 5960
rect 7980 5240 8020 5960
rect 7220 5200 8020 5240
rect 8632 5960 9432 6000
rect 8632 5240 8672 5960
rect 9392 5240 9432 5960
rect 8632 5200 9432 5240
rect 10044 5960 10844 6000
rect 10044 5240 10084 5960
rect 10804 5240 10844 5960
rect 10044 5200 10844 5240
rect 11456 5960 12256 6000
rect 11456 5240 11496 5960
rect 12216 5240 12256 5960
rect 11456 5200 12256 5240
rect 12868 5960 13668 6000
rect 12868 5240 12908 5960
rect 13628 5240 13668 5960
rect 12868 5200 13668 5240
rect 14280 5960 15080 6000
rect 14280 5240 14320 5960
rect 15040 5240 15080 5960
rect 14280 5200 15080 5240
rect 15692 5960 16492 6000
rect 15692 5240 15732 5960
rect 16452 5240 16492 5960
rect 15692 5200 16492 5240
rect 17104 5960 17904 6000
rect 17104 5240 17144 5960
rect 17864 5240 17904 5960
rect 17104 5200 17904 5240
rect 18516 5960 19316 6000
rect 18516 5240 18556 5960
rect 19276 5240 19316 5960
rect 18516 5200 19316 5240
rect 19928 5960 20728 6000
rect 19928 5240 19968 5960
rect 20688 5240 20728 5960
rect 19928 5200 20728 5240
rect 21340 5960 22140 6000
rect 21340 5240 21380 5960
rect 22100 5240 22140 5960
rect 21340 5200 22140 5240
rect 22752 5960 23552 6000
rect 22752 5240 22792 5960
rect 23512 5240 23552 5960
rect 22752 5200 23552 5240
rect -23844 4840 -23044 4880
rect -23844 4120 -23804 4840
rect -23084 4120 -23044 4840
rect -23844 4080 -23044 4120
rect -22432 4840 -21632 4880
rect -22432 4120 -22392 4840
rect -21672 4120 -21632 4840
rect -22432 4080 -21632 4120
rect -21020 4840 -20220 4880
rect -21020 4120 -20980 4840
rect -20260 4120 -20220 4840
rect -21020 4080 -20220 4120
rect -19608 4840 -18808 4880
rect -19608 4120 -19568 4840
rect -18848 4120 -18808 4840
rect -19608 4080 -18808 4120
rect -18196 4840 -17396 4880
rect -18196 4120 -18156 4840
rect -17436 4120 -17396 4840
rect -18196 4080 -17396 4120
rect -16784 4840 -15984 4880
rect -16784 4120 -16744 4840
rect -16024 4120 -15984 4840
rect -16784 4080 -15984 4120
rect -15372 4840 -14572 4880
rect -15372 4120 -15332 4840
rect -14612 4120 -14572 4840
rect -15372 4080 -14572 4120
rect -13960 4840 -13160 4880
rect -13960 4120 -13920 4840
rect -13200 4120 -13160 4840
rect -13960 4080 -13160 4120
rect -12548 4840 -11748 4880
rect -12548 4120 -12508 4840
rect -11788 4120 -11748 4840
rect -12548 4080 -11748 4120
rect -11136 4840 -10336 4880
rect -11136 4120 -11096 4840
rect -10376 4120 -10336 4840
rect -11136 4080 -10336 4120
rect -9724 4840 -8924 4880
rect -9724 4120 -9684 4840
rect -8964 4120 -8924 4840
rect -9724 4080 -8924 4120
rect -8312 4840 -7512 4880
rect -8312 4120 -8272 4840
rect -7552 4120 -7512 4840
rect -8312 4080 -7512 4120
rect -6900 4840 -6100 4880
rect -6900 4120 -6860 4840
rect -6140 4120 -6100 4840
rect -6900 4080 -6100 4120
rect -5488 4840 -4688 4880
rect -5488 4120 -5448 4840
rect -4728 4120 -4688 4840
rect -5488 4080 -4688 4120
rect -4076 4840 -3276 4880
rect -4076 4120 -4036 4840
rect -3316 4120 -3276 4840
rect -4076 4080 -3276 4120
rect -2664 4840 -1864 4880
rect -2664 4120 -2624 4840
rect -1904 4120 -1864 4840
rect -2664 4080 -1864 4120
rect -1252 4840 -452 4880
rect -1252 4120 -1212 4840
rect -492 4120 -452 4840
rect -1252 4080 -452 4120
rect 160 4840 960 4880
rect 160 4120 200 4840
rect 920 4120 960 4840
rect 160 4080 960 4120
rect 1572 4840 2372 4880
rect 1572 4120 1612 4840
rect 2332 4120 2372 4840
rect 1572 4080 2372 4120
rect 2984 4840 3784 4880
rect 2984 4120 3024 4840
rect 3744 4120 3784 4840
rect 2984 4080 3784 4120
rect 4396 4840 5196 4880
rect 4396 4120 4436 4840
rect 5156 4120 5196 4840
rect 4396 4080 5196 4120
rect 5808 4840 6608 4880
rect 5808 4120 5848 4840
rect 6568 4120 6608 4840
rect 5808 4080 6608 4120
rect 7220 4840 8020 4880
rect 7220 4120 7260 4840
rect 7980 4120 8020 4840
rect 7220 4080 8020 4120
rect 8632 4840 9432 4880
rect 8632 4120 8672 4840
rect 9392 4120 9432 4840
rect 8632 4080 9432 4120
rect 10044 4840 10844 4880
rect 10044 4120 10084 4840
rect 10804 4120 10844 4840
rect 10044 4080 10844 4120
rect 11456 4840 12256 4880
rect 11456 4120 11496 4840
rect 12216 4120 12256 4840
rect 11456 4080 12256 4120
rect 12868 4840 13668 4880
rect 12868 4120 12908 4840
rect 13628 4120 13668 4840
rect 12868 4080 13668 4120
rect 14280 4840 15080 4880
rect 14280 4120 14320 4840
rect 15040 4120 15080 4840
rect 14280 4080 15080 4120
rect 15692 4840 16492 4880
rect 15692 4120 15732 4840
rect 16452 4120 16492 4840
rect 15692 4080 16492 4120
rect 17104 4840 17904 4880
rect 17104 4120 17144 4840
rect 17864 4120 17904 4840
rect 17104 4080 17904 4120
rect 18516 4840 19316 4880
rect 18516 4120 18556 4840
rect 19276 4120 19316 4840
rect 18516 4080 19316 4120
rect 19928 4840 20728 4880
rect 19928 4120 19968 4840
rect 20688 4120 20728 4840
rect 19928 4080 20728 4120
rect 21340 4840 22140 4880
rect 21340 4120 21380 4840
rect 22100 4120 22140 4840
rect 21340 4080 22140 4120
rect 22752 4840 23552 4880
rect 22752 4120 22792 4840
rect 23512 4120 23552 4840
rect 22752 4080 23552 4120
rect -23844 3720 -23044 3760
rect -23844 3000 -23804 3720
rect -23084 3000 -23044 3720
rect -23844 2960 -23044 3000
rect -22432 3720 -21632 3760
rect -22432 3000 -22392 3720
rect -21672 3000 -21632 3720
rect -22432 2960 -21632 3000
rect -21020 3720 -20220 3760
rect -21020 3000 -20980 3720
rect -20260 3000 -20220 3720
rect -21020 2960 -20220 3000
rect -19608 3720 -18808 3760
rect -19608 3000 -19568 3720
rect -18848 3000 -18808 3720
rect -19608 2960 -18808 3000
rect -18196 3720 -17396 3760
rect -18196 3000 -18156 3720
rect -17436 3000 -17396 3720
rect -18196 2960 -17396 3000
rect -16784 3720 -15984 3760
rect -16784 3000 -16744 3720
rect -16024 3000 -15984 3720
rect -16784 2960 -15984 3000
rect -15372 3720 -14572 3760
rect -15372 3000 -15332 3720
rect -14612 3000 -14572 3720
rect -15372 2960 -14572 3000
rect -13960 3720 -13160 3760
rect -13960 3000 -13920 3720
rect -13200 3000 -13160 3720
rect -13960 2960 -13160 3000
rect -12548 3720 -11748 3760
rect -12548 3000 -12508 3720
rect -11788 3000 -11748 3720
rect -12548 2960 -11748 3000
rect -11136 3720 -10336 3760
rect -11136 3000 -11096 3720
rect -10376 3000 -10336 3720
rect -11136 2960 -10336 3000
rect -9724 3720 -8924 3760
rect -9724 3000 -9684 3720
rect -8964 3000 -8924 3720
rect -9724 2960 -8924 3000
rect -8312 3720 -7512 3760
rect -8312 3000 -8272 3720
rect -7552 3000 -7512 3720
rect -8312 2960 -7512 3000
rect -6900 3720 -6100 3760
rect -6900 3000 -6860 3720
rect -6140 3000 -6100 3720
rect -6900 2960 -6100 3000
rect -5488 3720 -4688 3760
rect -5488 3000 -5448 3720
rect -4728 3000 -4688 3720
rect -5488 2960 -4688 3000
rect -4076 3720 -3276 3760
rect -4076 3000 -4036 3720
rect -3316 3000 -3276 3720
rect -4076 2960 -3276 3000
rect -2664 3720 -1864 3760
rect -2664 3000 -2624 3720
rect -1904 3000 -1864 3720
rect -2664 2960 -1864 3000
rect -1252 3720 -452 3760
rect -1252 3000 -1212 3720
rect -492 3000 -452 3720
rect -1252 2960 -452 3000
rect 160 3720 960 3760
rect 160 3000 200 3720
rect 920 3000 960 3720
rect 160 2960 960 3000
rect 1572 3720 2372 3760
rect 1572 3000 1612 3720
rect 2332 3000 2372 3720
rect 1572 2960 2372 3000
rect 2984 3720 3784 3760
rect 2984 3000 3024 3720
rect 3744 3000 3784 3720
rect 2984 2960 3784 3000
rect 4396 3720 5196 3760
rect 4396 3000 4436 3720
rect 5156 3000 5196 3720
rect 4396 2960 5196 3000
rect 5808 3720 6608 3760
rect 5808 3000 5848 3720
rect 6568 3000 6608 3720
rect 5808 2960 6608 3000
rect 7220 3720 8020 3760
rect 7220 3000 7260 3720
rect 7980 3000 8020 3720
rect 7220 2960 8020 3000
rect 8632 3720 9432 3760
rect 8632 3000 8672 3720
rect 9392 3000 9432 3720
rect 8632 2960 9432 3000
rect 10044 3720 10844 3760
rect 10044 3000 10084 3720
rect 10804 3000 10844 3720
rect 10044 2960 10844 3000
rect 11456 3720 12256 3760
rect 11456 3000 11496 3720
rect 12216 3000 12256 3720
rect 11456 2960 12256 3000
rect 12868 3720 13668 3760
rect 12868 3000 12908 3720
rect 13628 3000 13668 3720
rect 12868 2960 13668 3000
rect 14280 3720 15080 3760
rect 14280 3000 14320 3720
rect 15040 3000 15080 3720
rect 14280 2960 15080 3000
rect 15692 3720 16492 3760
rect 15692 3000 15732 3720
rect 16452 3000 16492 3720
rect 15692 2960 16492 3000
rect 17104 3720 17904 3760
rect 17104 3000 17144 3720
rect 17864 3000 17904 3720
rect 17104 2960 17904 3000
rect 18516 3720 19316 3760
rect 18516 3000 18556 3720
rect 19276 3000 19316 3720
rect 18516 2960 19316 3000
rect 19928 3720 20728 3760
rect 19928 3000 19968 3720
rect 20688 3000 20728 3720
rect 19928 2960 20728 3000
rect 21340 3720 22140 3760
rect 21340 3000 21380 3720
rect 22100 3000 22140 3720
rect 21340 2960 22140 3000
rect 22752 3720 23552 3760
rect 22752 3000 22792 3720
rect 23512 3000 23552 3720
rect 22752 2960 23552 3000
rect -23844 2600 -23044 2640
rect -23844 1880 -23804 2600
rect -23084 1880 -23044 2600
rect -23844 1840 -23044 1880
rect -22432 2600 -21632 2640
rect -22432 1880 -22392 2600
rect -21672 1880 -21632 2600
rect -22432 1840 -21632 1880
rect -21020 2600 -20220 2640
rect -21020 1880 -20980 2600
rect -20260 1880 -20220 2600
rect -21020 1840 -20220 1880
rect -19608 2600 -18808 2640
rect -19608 1880 -19568 2600
rect -18848 1880 -18808 2600
rect -19608 1840 -18808 1880
rect -18196 2600 -17396 2640
rect -18196 1880 -18156 2600
rect -17436 1880 -17396 2600
rect -18196 1840 -17396 1880
rect -16784 2600 -15984 2640
rect -16784 1880 -16744 2600
rect -16024 1880 -15984 2600
rect -16784 1840 -15984 1880
rect -15372 2600 -14572 2640
rect -15372 1880 -15332 2600
rect -14612 1880 -14572 2600
rect -15372 1840 -14572 1880
rect -13960 2600 -13160 2640
rect -13960 1880 -13920 2600
rect -13200 1880 -13160 2600
rect -13960 1840 -13160 1880
rect -12548 2600 -11748 2640
rect -12548 1880 -12508 2600
rect -11788 1880 -11748 2600
rect -12548 1840 -11748 1880
rect -11136 2600 -10336 2640
rect -11136 1880 -11096 2600
rect -10376 1880 -10336 2600
rect -11136 1840 -10336 1880
rect -9724 2600 -8924 2640
rect -9724 1880 -9684 2600
rect -8964 1880 -8924 2600
rect -9724 1840 -8924 1880
rect -8312 2600 -7512 2640
rect -8312 1880 -8272 2600
rect -7552 1880 -7512 2600
rect -8312 1840 -7512 1880
rect -6900 2600 -6100 2640
rect -6900 1880 -6860 2600
rect -6140 1880 -6100 2600
rect -6900 1840 -6100 1880
rect -5488 2600 -4688 2640
rect -5488 1880 -5448 2600
rect -4728 1880 -4688 2600
rect -5488 1840 -4688 1880
rect -4076 2600 -3276 2640
rect -4076 1880 -4036 2600
rect -3316 1880 -3276 2600
rect -4076 1840 -3276 1880
rect -2664 2600 -1864 2640
rect -2664 1880 -2624 2600
rect -1904 1880 -1864 2600
rect -2664 1840 -1864 1880
rect -1252 2600 -452 2640
rect -1252 1880 -1212 2600
rect -492 1880 -452 2600
rect -1252 1840 -452 1880
rect 160 2600 960 2640
rect 160 1880 200 2600
rect 920 1880 960 2600
rect 160 1840 960 1880
rect 1572 2600 2372 2640
rect 1572 1880 1612 2600
rect 2332 1880 2372 2600
rect 1572 1840 2372 1880
rect 2984 2600 3784 2640
rect 2984 1880 3024 2600
rect 3744 1880 3784 2600
rect 2984 1840 3784 1880
rect 4396 2600 5196 2640
rect 4396 1880 4436 2600
rect 5156 1880 5196 2600
rect 4396 1840 5196 1880
rect 5808 2600 6608 2640
rect 5808 1880 5848 2600
rect 6568 1880 6608 2600
rect 5808 1840 6608 1880
rect 7220 2600 8020 2640
rect 7220 1880 7260 2600
rect 7980 1880 8020 2600
rect 7220 1840 8020 1880
rect 8632 2600 9432 2640
rect 8632 1880 8672 2600
rect 9392 1880 9432 2600
rect 8632 1840 9432 1880
rect 10044 2600 10844 2640
rect 10044 1880 10084 2600
rect 10804 1880 10844 2600
rect 10044 1840 10844 1880
rect 11456 2600 12256 2640
rect 11456 1880 11496 2600
rect 12216 1880 12256 2600
rect 11456 1840 12256 1880
rect 12868 2600 13668 2640
rect 12868 1880 12908 2600
rect 13628 1880 13668 2600
rect 12868 1840 13668 1880
rect 14280 2600 15080 2640
rect 14280 1880 14320 2600
rect 15040 1880 15080 2600
rect 14280 1840 15080 1880
rect 15692 2600 16492 2640
rect 15692 1880 15732 2600
rect 16452 1880 16492 2600
rect 15692 1840 16492 1880
rect 17104 2600 17904 2640
rect 17104 1880 17144 2600
rect 17864 1880 17904 2600
rect 17104 1840 17904 1880
rect 18516 2600 19316 2640
rect 18516 1880 18556 2600
rect 19276 1880 19316 2600
rect 18516 1840 19316 1880
rect 19928 2600 20728 2640
rect 19928 1880 19968 2600
rect 20688 1880 20728 2600
rect 19928 1840 20728 1880
rect 21340 2600 22140 2640
rect 21340 1880 21380 2600
rect 22100 1880 22140 2600
rect 21340 1840 22140 1880
rect 22752 2600 23552 2640
rect 22752 1880 22792 2600
rect 23512 1880 23552 2600
rect 22752 1840 23552 1880
rect -23844 1480 -23044 1520
rect -23844 760 -23804 1480
rect -23084 760 -23044 1480
rect -23844 720 -23044 760
rect -22432 1480 -21632 1520
rect -22432 760 -22392 1480
rect -21672 760 -21632 1480
rect -22432 720 -21632 760
rect -21020 1480 -20220 1520
rect -21020 760 -20980 1480
rect -20260 760 -20220 1480
rect -21020 720 -20220 760
rect -19608 1480 -18808 1520
rect -19608 760 -19568 1480
rect -18848 760 -18808 1480
rect -19608 720 -18808 760
rect -18196 1480 -17396 1520
rect -18196 760 -18156 1480
rect -17436 760 -17396 1480
rect -18196 720 -17396 760
rect -16784 1480 -15984 1520
rect -16784 760 -16744 1480
rect -16024 760 -15984 1480
rect -16784 720 -15984 760
rect -15372 1480 -14572 1520
rect -15372 760 -15332 1480
rect -14612 760 -14572 1480
rect -15372 720 -14572 760
rect -13960 1480 -13160 1520
rect -13960 760 -13920 1480
rect -13200 760 -13160 1480
rect -13960 720 -13160 760
rect -12548 1480 -11748 1520
rect -12548 760 -12508 1480
rect -11788 760 -11748 1480
rect -12548 720 -11748 760
rect -11136 1480 -10336 1520
rect -11136 760 -11096 1480
rect -10376 760 -10336 1480
rect -11136 720 -10336 760
rect -9724 1480 -8924 1520
rect -9724 760 -9684 1480
rect -8964 760 -8924 1480
rect -9724 720 -8924 760
rect -8312 1480 -7512 1520
rect -8312 760 -8272 1480
rect -7552 760 -7512 1480
rect -8312 720 -7512 760
rect -6900 1480 -6100 1520
rect -6900 760 -6860 1480
rect -6140 760 -6100 1480
rect -6900 720 -6100 760
rect -5488 1480 -4688 1520
rect -5488 760 -5448 1480
rect -4728 760 -4688 1480
rect -5488 720 -4688 760
rect -4076 1480 -3276 1520
rect -4076 760 -4036 1480
rect -3316 760 -3276 1480
rect -4076 720 -3276 760
rect -2664 1480 -1864 1520
rect -2664 760 -2624 1480
rect -1904 760 -1864 1480
rect -2664 720 -1864 760
rect -1252 1480 -452 1520
rect -1252 760 -1212 1480
rect -492 760 -452 1480
rect -1252 720 -452 760
rect 160 1480 960 1520
rect 160 760 200 1480
rect 920 760 960 1480
rect 160 720 960 760
rect 1572 1480 2372 1520
rect 1572 760 1612 1480
rect 2332 760 2372 1480
rect 1572 720 2372 760
rect 2984 1480 3784 1520
rect 2984 760 3024 1480
rect 3744 760 3784 1480
rect 2984 720 3784 760
rect 4396 1480 5196 1520
rect 4396 760 4436 1480
rect 5156 760 5196 1480
rect 4396 720 5196 760
rect 5808 1480 6608 1520
rect 5808 760 5848 1480
rect 6568 760 6608 1480
rect 5808 720 6608 760
rect 7220 1480 8020 1520
rect 7220 760 7260 1480
rect 7980 760 8020 1480
rect 7220 720 8020 760
rect 8632 1480 9432 1520
rect 8632 760 8672 1480
rect 9392 760 9432 1480
rect 8632 720 9432 760
rect 10044 1480 10844 1520
rect 10044 760 10084 1480
rect 10804 760 10844 1480
rect 10044 720 10844 760
rect 11456 1480 12256 1520
rect 11456 760 11496 1480
rect 12216 760 12256 1480
rect 11456 720 12256 760
rect 12868 1480 13668 1520
rect 12868 760 12908 1480
rect 13628 760 13668 1480
rect 12868 720 13668 760
rect 14280 1480 15080 1520
rect 14280 760 14320 1480
rect 15040 760 15080 1480
rect 14280 720 15080 760
rect 15692 1480 16492 1520
rect 15692 760 15732 1480
rect 16452 760 16492 1480
rect 15692 720 16492 760
rect 17104 1480 17904 1520
rect 17104 760 17144 1480
rect 17864 760 17904 1480
rect 17104 720 17904 760
rect 18516 1480 19316 1520
rect 18516 760 18556 1480
rect 19276 760 19316 1480
rect 18516 720 19316 760
rect 19928 1480 20728 1520
rect 19928 760 19968 1480
rect 20688 760 20728 1480
rect 19928 720 20728 760
rect 21340 1480 22140 1520
rect 21340 760 21380 1480
rect 22100 760 22140 1480
rect 21340 720 22140 760
rect 22752 1480 23552 1520
rect 22752 760 22792 1480
rect 23512 760 23552 1480
rect 22752 720 23552 760
rect -23844 360 -23044 400
rect -23844 -360 -23804 360
rect -23084 -360 -23044 360
rect -23844 -400 -23044 -360
rect -22432 360 -21632 400
rect -22432 -360 -22392 360
rect -21672 -360 -21632 360
rect -22432 -400 -21632 -360
rect -21020 360 -20220 400
rect -21020 -360 -20980 360
rect -20260 -360 -20220 360
rect -21020 -400 -20220 -360
rect -19608 360 -18808 400
rect -19608 -360 -19568 360
rect -18848 -360 -18808 360
rect -19608 -400 -18808 -360
rect -18196 360 -17396 400
rect -18196 -360 -18156 360
rect -17436 -360 -17396 360
rect -18196 -400 -17396 -360
rect -16784 360 -15984 400
rect -16784 -360 -16744 360
rect -16024 -360 -15984 360
rect -16784 -400 -15984 -360
rect -15372 360 -14572 400
rect -15372 -360 -15332 360
rect -14612 -360 -14572 360
rect -15372 -400 -14572 -360
rect -13960 360 -13160 400
rect -13960 -360 -13920 360
rect -13200 -360 -13160 360
rect -13960 -400 -13160 -360
rect -12548 360 -11748 400
rect -12548 -360 -12508 360
rect -11788 -360 -11748 360
rect -12548 -400 -11748 -360
rect -11136 360 -10336 400
rect -11136 -360 -11096 360
rect -10376 -360 -10336 360
rect -11136 -400 -10336 -360
rect -9724 360 -8924 400
rect -9724 -360 -9684 360
rect -8964 -360 -8924 360
rect -9724 -400 -8924 -360
rect -8312 360 -7512 400
rect -8312 -360 -8272 360
rect -7552 -360 -7512 360
rect -8312 -400 -7512 -360
rect -6900 360 -6100 400
rect -6900 -360 -6860 360
rect -6140 -360 -6100 360
rect -6900 -400 -6100 -360
rect -5488 360 -4688 400
rect -5488 -360 -5448 360
rect -4728 -360 -4688 360
rect -5488 -400 -4688 -360
rect -4076 360 -3276 400
rect -4076 -360 -4036 360
rect -3316 -360 -3276 360
rect -4076 -400 -3276 -360
rect -2664 360 -1864 400
rect -2664 -360 -2624 360
rect -1904 -360 -1864 360
rect -2664 -400 -1864 -360
rect -1252 360 -452 400
rect -1252 -360 -1212 360
rect -492 -360 -452 360
rect -1252 -400 -452 -360
rect 160 360 960 400
rect 160 -360 200 360
rect 920 -360 960 360
rect 160 -400 960 -360
rect 1572 360 2372 400
rect 1572 -360 1612 360
rect 2332 -360 2372 360
rect 1572 -400 2372 -360
rect 2984 360 3784 400
rect 2984 -360 3024 360
rect 3744 -360 3784 360
rect 2984 -400 3784 -360
rect 4396 360 5196 400
rect 4396 -360 4436 360
rect 5156 -360 5196 360
rect 4396 -400 5196 -360
rect 5808 360 6608 400
rect 5808 -360 5848 360
rect 6568 -360 6608 360
rect 5808 -400 6608 -360
rect 7220 360 8020 400
rect 7220 -360 7260 360
rect 7980 -360 8020 360
rect 7220 -400 8020 -360
rect 8632 360 9432 400
rect 8632 -360 8672 360
rect 9392 -360 9432 360
rect 8632 -400 9432 -360
rect 10044 360 10844 400
rect 10044 -360 10084 360
rect 10804 -360 10844 360
rect 10044 -400 10844 -360
rect 11456 360 12256 400
rect 11456 -360 11496 360
rect 12216 -360 12256 360
rect 11456 -400 12256 -360
rect 12868 360 13668 400
rect 12868 -360 12908 360
rect 13628 -360 13668 360
rect 12868 -400 13668 -360
rect 14280 360 15080 400
rect 14280 -360 14320 360
rect 15040 -360 15080 360
rect 14280 -400 15080 -360
rect 15692 360 16492 400
rect 15692 -360 15732 360
rect 16452 -360 16492 360
rect 15692 -400 16492 -360
rect 17104 360 17904 400
rect 17104 -360 17144 360
rect 17864 -360 17904 360
rect 17104 -400 17904 -360
rect 18516 360 19316 400
rect 18516 -360 18556 360
rect 19276 -360 19316 360
rect 18516 -400 19316 -360
rect 19928 360 20728 400
rect 19928 -360 19968 360
rect 20688 -360 20728 360
rect 19928 -400 20728 -360
rect 21340 360 22140 400
rect 21340 -360 21380 360
rect 22100 -360 22140 360
rect 21340 -400 22140 -360
rect 22752 360 23552 400
rect 22752 -360 22792 360
rect 23512 -360 23552 360
rect 22752 -400 23552 -360
rect -23844 -760 -23044 -720
rect -23844 -1480 -23804 -760
rect -23084 -1480 -23044 -760
rect -23844 -1520 -23044 -1480
rect -22432 -760 -21632 -720
rect -22432 -1480 -22392 -760
rect -21672 -1480 -21632 -760
rect -22432 -1520 -21632 -1480
rect -21020 -760 -20220 -720
rect -21020 -1480 -20980 -760
rect -20260 -1480 -20220 -760
rect -21020 -1520 -20220 -1480
rect -19608 -760 -18808 -720
rect -19608 -1480 -19568 -760
rect -18848 -1480 -18808 -760
rect -19608 -1520 -18808 -1480
rect -18196 -760 -17396 -720
rect -18196 -1480 -18156 -760
rect -17436 -1480 -17396 -760
rect -18196 -1520 -17396 -1480
rect -16784 -760 -15984 -720
rect -16784 -1480 -16744 -760
rect -16024 -1480 -15984 -760
rect -16784 -1520 -15984 -1480
rect -15372 -760 -14572 -720
rect -15372 -1480 -15332 -760
rect -14612 -1480 -14572 -760
rect -15372 -1520 -14572 -1480
rect -13960 -760 -13160 -720
rect -13960 -1480 -13920 -760
rect -13200 -1480 -13160 -760
rect -13960 -1520 -13160 -1480
rect -12548 -760 -11748 -720
rect -12548 -1480 -12508 -760
rect -11788 -1480 -11748 -760
rect -12548 -1520 -11748 -1480
rect -11136 -760 -10336 -720
rect -11136 -1480 -11096 -760
rect -10376 -1480 -10336 -760
rect -11136 -1520 -10336 -1480
rect -9724 -760 -8924 -720
rect -9724 -1480 -9684 -760
rect -8964 -1480 -8924 -760
rect -9724 -1520 -8924 -1480
rect -8312 -760 -7512 -720
rect -8312 -1480 -8272 -760
rect -7552 -1480 -7512 -760
rect -8312 -1520 -7512 -1480
rect -6900 -760 -6100 -720
rect -6900 -1480 -6860 -760
rect -6140 -1480 -6100 -760
rect -6900 -1520 -6100 -1480
rect -5488 -760 -4688 -720
rect -5488 -1480 -5448 -760
rect -4728 -1480 -4688 -760
rect -5488 -1520 -4688 -1480
rect -4076 -760 -3276 -720
rect -4076 -1480 -4036 -760
rect -3316 -1480 -3276 -760
rect -4076 -1520 -3276 -1480
rect -2664 -760 -1864 -720
rect -2664 -1480 -2624 -760
rect -1904 -1480 -1864 -760
rect -2664 -1520 -1864 -1480
rect -1252 -760 -452 -720
rect -1252 -1480 -1212 -760
rect -492 -1480 -452 -760
rect -1252 -1520 -452 -1480
rect 160 -760 960 -720
rect 160 -1480 200 -760
rect 920 -1480 960 -760
rect 160 -1520 960 -1480
rect 1572 -760 2372 -720
rect 1572 -1480 1612 -760
rect 2332 -1480 2372 -760
rect 1572 -1520 2372 -1480
rect 2984 -760 3784 -720
rect 2984 -1480 3024 -760
rect 3744 -1480 3784 -760
rect 2984 -1520 3784 -1480
rect 4396 -760 5196 -720
rect 4396 -1480 4436 -760
rect 5156 -1480 5196 -760
rect 4396 -1520 5196 -1480
rect 5808 -760 6608 -720
rect 5808 -1480 5848 -760
rect 6568 -1480 6608 -760
rect 5808 -1520 6608 -1480
rect 7220 -760 8020 -720
rect 7220 -1480 7260 -760
rect 7980 -1480 8020 -760
rect 7220 -1520 8020 -1480
rect 8632 -760 9432 -720
rect 8632 -1480 8672 -760
rect 9392 -1480 9432 -760
rect 8632 -1520 9432 -1480
rect 10044 -760 10844 -720
rect 10044 -1480 10084 -760
rect 10804 -1480 10844 -760
rect 10044 -1520 10844 -1480
rect 11456 -760 12256 -720
rect 11456 -1480 11496 -760
rect 12216 -1480 12256 -760
rect 11456 -1520 12256 -1480
rect 12868 -760 13668 -720
rect 12868 -1480 12908 -760
rect 13628 -1480 13668 -760
rect 12868 -1520 13668 -1480
rect 14280 -760 15080 -720
rect 14280 -1480 14320 -760
rect 15040 -1480 15080 -760
rect 14280 -1520 15080 -1480
rect 15692 -760 16492 -720
rect 15692 -1480 15732 -760
rect 16452 -1480 16492 -760
rect 15692 -1520 16492 -1480
rect 17104 -760 17904 -720
rect 17104 -1480 17144 -760
rect 17864 -1480 17904 -760
rect 17104 -1520 17904 -1480
rect 18516 -760 19316 -720
rect 18516 -1480 18556 -760
rect 19276 -1480 19316 -760
rect 18516 -1520 19316 -1480
rect 19928 -760 20728 -720
rect 19928 -1480 19968 -760
rect 20688 -1480 20728 -760
rect 19928 -1520 20728 -1480
rect 21340 -760 22140 -720
rect 21340 -1480 21380 -760
rect 22100 -1480 22140 -760
rect 21340 -1520 22140 -1480
rect 22752 -760 23552 -720
rect 22752 -1480 22792 -760
rect 23512 -1480 23552 -760
rect 22752 -1520 23552 -1480
rect -23844 -1880 -23044 -1840
rect -23844 -2600 -23804 -1880
rect -23084 -2600 -23044 -1880
rect -23844 -2640 -23044 -2600
rect -22432 -1880 -21632 -1840
rect -22432 -2600 -22392 -1880
rect -21672 -2600 -21632 -1880
rect -22432 -2640 -21632 -2600
rect -21020 -1880 -20220 -1840
rect -21020 -2600 -20980 -1880
rect -20260 -2600 -20220 -1880
rect -21020 -2640 -20220 -2600
rect -19608 -1880 -18808 -1840
rect -19608 -2600 -19568 -1880
rect -18848 -2600 -18808 -1880
rect -19608 -2640 -18808 -2600
rect -18196 -1880 -17396 -1840
rect -18196 -2600 -18156 -1880
rect -17436 -2600 -17396 -1880
rect -18196 -2640 -17396 -2600
rect -16784 -1880 -15984 -1840
rect -16784 -2600 -16744 -1880
rect -16024 -2600 -15984 -1880
rect -16784 -2640 -15984 -2600
rect -15372 -1880 -14572 -1840
rect -15372 -2600 -15332 -1880
rect -14612 -2600 -14572 -1880
rect -15372 -2640 -14572 -2600
rect -13960 -1880 -13160 -1840
rect -13960 -2600 -13920 -1880
rect -13200 -2600 -13160 -1880
rect -13960 -2640 -13160 -2600
rect -12548 -1880 -11748 -1840
rect -12548 -2600 -12508 -1880
rect -11788 -2600 -11748 -1880
rect -12548 -2640 -11748 -2600
rect -11136 -1880 -10336 -1840
rect -11136 -2600 -11096 -1880
rect -10376 -2600 -10336 -1880
rect -11136 -2640 -10336 -2600
rect -9724 -1880 -8924 -1840
rect -9724 -2600 -9684 -1880
rect -8964 -2600 -8924 -1880
rect -9724 -2640 -8924 -2600
rect -8312 -1880 -7512 -1840
rect -8312 -2600 -8272 -1880
rect -7552 -2600 -7512 -1880
rect -8312 -2640 -7512 -2600
rect -6900 -1880 -6100 -1840
rect -6900 -2600 -6860 -1880
rect -6140 -2600 -6100 -1880
rect -6900 -2640 -6100 -2600
rect -5488 -1880 -4688 -1840
rect -5488 -2600 -5448 -1880
rect -4728 -2600 -4688 -1880
rect -5488 -2640 -4688 -2600
rect -4076 -1880 -3276 -1840
rect -4076 -2600 -4036 -1880
rect -3316 -2600 -3276 -1880
rect -4076 -2640 -3276 -2600
rect -2664 -1880 -1864 -1840
rect -2664 -2600 -2624 -1880
rect -1904 -2600 -1864 -1880
rect -2664 -2640 -1864 -2600
rect -1252 -1880 -452 -1840
rect -1252 -2600 -1212 -1880
rect -492 -2600 -452 -1880
rect -1252 -2640 -452 -2600
rect 160 -1880 960 -1840
rect 160 -2600 200 -1880
rect 920 -2600 960 -1880
rect 160 -2640 960 -2600
rect 1572 -1880 2372 -1840
rect 1572 -2600 1612 -1880
rect 2332 -2600 2372 -1880
rect 1572 -2640 2372 -2600
rect 2984 -1880 3784 -1840
rect 2984 -2600 3024 -1880
rect 3744 -2600 3784 -1880
rect 2984 -2640 3784 -2600
rect 4396 -1880 5196 -1840
rect 4396 -2600 4436 -1880
rect 5156 -2600 5196 -1880
rect 4396 -2640 5196 -2600
rect 5808 -1880 6608 -1840
rect 5808 -2600 5848 -1880
rect 6568 -2600 6608 -1880
rect 5808 -2640 6608 -2600
rect 7220 -1880 8020 -1840
rect 7220 -2600 7260 -1880
rect 7980 -2600 8020 -1880
rect 7220 -2640 8020 -2600
rect 8632 -1880 9432 -1840
rect 8632 -2600 8672 -1880
rect 9392 -2600 9432 -1880
rect 8632 -2640 9432 -2600
rect 10044 -1880 10844 -1840
rect 10044 -2600 10084 -1880
rect 10804 -2600 10844 -1880
rect 10044 -2640 10844 -2600
rect 11456 -1880 12256 -1840
rect 11456 -2600 11496 -1880
rect 12216 -2600 12256 -1880
rect 11456 -2640 12256 -2600
rect 12868 -1880 13668 -1840
rect 12868 -2600 12908 -1880
rect 13628 -2600 13668 -1880
rect 12868 -2640 13668 -2600
rect 14280 -1880 15080 -1840
rect 14280 -2600 14320 -1880
rect 15040 -2600 15080 -1880
rect 14280 -2640 15080 -2600
rect 15692 -1880 16492 -1840
rect 15692 -2600 15732 -1880
rect 16452 -2600 16492 -1880
rect 15692 -2640 16492 -2600
rect 17104 -1880 17904 -1840
rect 17104 -2600 17144 -1880
rect 17864 -2600 17904 -1880
rect 17104 -2640 17904 -2600
rect 18516 -1880 19316 -1840
rect 18516 -2600 18556 -1880
rect 19276 -2600 19316 -1880
rect 18516 -2640 19316 -2600
rect 19928 -1880 20728 -1840
rect 19928 -2600 19968 -1880
rect 20688 -2600 20728 -1880
rect 19928 -2640 20728 -2600
rect 21340 -1880 22140 -1840
rect 21340 -2600 21380 -1880
rect 22100 -2600 22140 -1880
rect 21340 -2640 22140 -2600
rect 22752 -1880 23552 -1840
rect 22752 -2600 22792 -1880
rect 23512 -2600 23552 -1880
rect 22752 -2640 23552 -2600
rect -23844 -3000 -23044 -2960
rect -23844 -3720 -23804 -3000
rect -23084 -3720 -23044 -3000
rect -23844 -3760 -23044 -3720
rect -22432 -3000 -21632 -2960
rect -22432 -3720 -22392 -3000
rect -21672 -3720 -21632 -3000
rect -22432 -3760 -21632 -3720
rect -21020 -3000 -20220 -2960
rect -21020 -3720 -20980 -3000
rect -20260 -3720 -20220 -3000
rect -21020 -3760 -20220 -3720
rect -19608 -3000 -18808 -2960
rect -19608 -3720 -19568 -3000
rect -18848 -3720 -18808 -3000
rect -19608 -3760 -18808 -3720
rect -18196 -3000 -17396 -2960
rect -18196 -3720 -18156 -3000
rect -17436 -3720 -17396 -3000
rect -18196 -3760 -17396 -3720
rect -16784 -3000 -15984 -2960
rect -16784 -3720 -16744 -3000
rect -16024 -3720 -15984 -3000
rect -16784 -3760 -15984 -3720
rect -15372 -3000 -14572 -2960
rect -15372 -3720 -15332 -3000
rect -14612 -3720 -14572 -3000
rect -15372 -3760 -14572 -3720
rect -13960 -3000 -13160 -2960
rect -13960 -3720 -13920 -3000
rect -13200 -3720 -13160 -3000
rect -13960 -3760 -13160 -3720
rect -12548 -3000 -11748 -2960
rect -12548 -3720 -12508 -3000
rect -11788 -3720 -11748 -3000
rect -12548 -3760 -11748 -3720
rect -11136 -3000 -10336 -2960
rect -11136 -3720 -11096 -3000
rect -10376 -3720 -10336 -3000
rect -11136 -3760 -10336 -3720
rect -9724 -3000 -8924 -2960
rect -9724 -3720 -9684 -3000
rect -8964 -3720 -8924 -3000
rect -9724 -3760 -8924 -3720
rect -8312 -3000 -7512 -2960
rect -8312 -3720 -8272 -3000
rect -7552 -3720 -7512 -3000
rect -8312 -3760 -7512 -3720
rect -6900 -3000 -6100 -2960
rect -6900 -3720 -6860 -3000
rect -6140 -3720 -6100 -3000
rect -6900 -3760 -6100 -3720
rect -5488 -3000 -4688 -2960
rect -5488 -3720 -5448 -3000
rect -4728 -3720 -4688 -3000
rect -5488 -3760 -4688 -3720
rect -4076 -3000 -3276 -2960
rect -4076 -3720 -4036 -3000
rect -3316 -3720 -3276 -3000
rect -4076 -3760 -3276 -3720
rect -2664 -3000 -1864 -2960
rect -2664 -3720 -2624 -3000
rect -1904 -3720 -1864 -3000
rect -2664 -3760 -1864 -3720
rect -1252 -3000 -452 -2960
rect -1252 -3720 -1212 -3000
rect -492 -3720 -452 -3000
rect -1252 -3760 -452 -3720
rect 160 -3000 960 -2960
rect 160 -3720 200 -3000
rect 920 -3720 960 -3000
rect 160 -3760 960 -3720
rect 1572 -3000 2372 -2960
rect 1572 -3720 1612 -3000
rect 2332 -3720 2372 -3000
rect 1572 -3760 2372 -3720
rect 2984 -3000 3784 -2960
rect 2984 -3720 3024 -3000
rect 3744 -3720 3784 -3000
rect 2984 -3760 3784 -3720
rect 4396 -3000 5196 -2960
rect 4396 -3720 4436 -3000
rect 5156 -3720 5196 -3000
rect 4396 -3760 5196 -3720
rect 5808 -3000 6608 -2960
rect 5808 -3720 5848 -3000
rect 6568 -3720 6608 -3000
rect 5808 -3760 6608 -3720
rect 7220 -3000 8020 -2960
rect 7220 -3720 7260 -3000
rect 7980 -3720 8020 -3000
rect 7220 -3760 8020 -3720
rect 8632 -3000 9432 -2960
rect 8632 -3720 8672 -3000
rect 9392 -3720 9432 -3000
rect 8632 -3760 9432 -3720
rect 10044 -3000 10844 -2960
rect 10044 -3720 10084 -3000
rect 10804 -3720 10844 -3000
rect 10044 -3760 10844 -3720
rect 11456 -3000 12256 -2960
rect 11456 -3720 11496 -3000
rect 12216 -3720 12256 -3000
rect 11456 -3760 12256 -3720
rect 12868 -3000 13668 -2960
rect 12868 -3720 12908 -3000
rect 13628 -3720 13668 -3000
rect 12868 -3760 13668 -3720
rect 14280 -3000 15080 -2960
rect 14280 -3720 14320 -3000
rect 15040 -3720 15080 -3000
rect 14280 -3760 15080 -3720
rect 15692 -3000 16492 -2960
rect 15692 -3720 15732 -3000
rect 16452 -3720 16492 -3000
rect 15692 -3760 16492 -3720
rect 17104 -3000 17904 -2960
rect 17104 -3720 17144 -3000
rect 17864 -3720 17904 -3000
rect 17104 -3760 17904 -3720
rect 18516 -3000 19316 -2960
rect 18516 -3720 18556 -3000
rect 19276 -3720 19316 -3000
rect 18516 -3760 19316 -3720
rect 19928 -3000 20728 -2960
rect 19928 -3720 19968 -3000
rect 20688 -3720 20728 -3000
rect 19928 -3760 20728 -3720
rect 21340 -3000 22140 -2960
rect 21340 -3720 21380 -3000
rect 22100 -3720 22140 -3000
rect 21340 -3760 22140 -3720
rect 22752 -3000 23552 -2960
rect 22752 -3720 22792 -3000
rect 23512 -3720 23552 -3000
rect 22752 -3760 23552 -3720
rect -23844 -4120 -23044 -4080
rect -23844 -4840 -23804 -4120
rect -23084 -4840 -23044 -4120
rect -23844 -4880 -23044 -4840
rect -22432 -4120 -21632 -4080
rect -22432 -4840 -22392 -4120
rect -21672 -4840 -21632 -4120
rect -22432 -4880 -21632 -4840
rect -21020 -4120 -20220 -4080
rect -21020 -4840 -20980 -4120
rect -20260 -4840 -20220 -4120
rect -21020 -4880 -20220 -4840
rect -19608 -4120 -18808 -4080
rect -19608 -4840 -19568 -4120
rect -18848 -4840 -18808 -4120
rect -19608 -4880 -18808 -4840
rect -18196 -4120 -17396 -4080
rect -18196 -4840 -18156 -4120
rect -17436 -4840 -17396 -4120
rect -18196 -4880 -17396 -4840
rect -16784 -4120 -15984 -4080
rect -16784 -4840 -16744 -4120
rect -16024 -4840 -15984 -4120
rect -16784 -4880 -15984 -4840
rect -15372 -4120 -14572 -4080
rect -15372 -4840 -15332 -4120
rect -14612 -4840 -14572 -4120
rect -15372 -4880 -14572 -4840
rect -13960 -4120 -13160 -4080
rect -13960 -4840 -13920 -4120
rect -13200 -4840 -13160 -4120
rect -13960 -4880 -13160 -4840
rect -12548 -4120 -11748 -4080
rect -12548 -4840 -12508 -4120
rect -11788 -4840 -11748 -4120
rect -12548 -4880 -11748 -4840
rect -11136 -4120 -10336 -4080
rect -11136 -4840 -11096 -4120
rect -10376 -4840 -10336 -4120
rect -11136 -4880 -10336 -4840
rect -9724 -4120 -8924 -4080
rect -9724 -4840 -9684 -4120
rect -8964 -4840 -8924 -4120
rect -9724 -4880 -8924 -4840
rect -8312 -4120 -7512 -4080
rect -8312 -4840 -8272 -4120
rect -7552 -4840 -7512 -4120
rect -8312 -4880 -7512 -4840
rect -6900 -4120 -6100 -4080
rect -6900 -4840 -6860 -4120
rect -6140 -4840 -6100 -4120
rect -6900 -4880 -6100 -4840
rect -5488 -4120 -4688 -4080
rect -5488 -4840 -5448 -4120
rect -4728 -4840 -4688 -4120
rect -5488 -4880 -4688 -4840
rect -4076 -4120 -3276 -4080
rect -4076 -4840 -4036 -4120
rect -3316 -4840 -3276 -4120
rect -4076 -4880 -3276 -4840
rect -2664 -4120 -1864 -4080
rect -2664 -4840 -2624 -4120
rect -1904 -4840 -1864 -4120
rect -2664 -4880 -1864 -4840
rect -1252 -4120 -452 -4080
rect -1252 -4840 -1212 -4120
rect -492 -4840 -452 -4120
rect -1252 -4880 -452 -4840
rect 160 -4120 960 -4080
rect 160 -4840 200 -4120
rect 920 -4840 960 -4120
rect 160 -4880 960 -4840
rect 1572 -4120 2372 -4080
rect 1572 -4840 1612 -4120
rect 2332 -4840 2372 -4120
rect 1572 -4880 2372 -4840
rect 2984 -4120 3784 -4080
rect 2984 -4840 3024 -4120
rect 3744 -4840 3784 -4120
rect 2984 -4880 3784 -4840
rect 4396 -4120 5196 -4080
rect 4396 -4840 4436 -4120
rect 5156 -4840 5196 -4120
rect 4396 -4880 5196 -4840
rect 5808 -4120 6608 -4080
rect 5808 -4840 5848 -4120
rect 6568 -4840 6608 -4120
rect 5808 -4880 6608 -4840
rect 7220 -4120 8020 -4080
rect 7220 -4840 7260 -4120
rect 7980 -4840 8020 -4120
rect 7220 -4880 8020 -4840
rect 8632 -4120 9432 -4080
rect 8632 -4840 8672 -4120
rect 9392 -4840 9432 -4120
rect 8632 -4880 9432 -4840
rect 10044 -4120 10844 -4080
rect 10044 -4840 10084 -4120
rect 10804 -4840 10844 -4120
rect 10044 -4880 10844 -4840
rect 11456 -4120 12256 -4080
rect 11456 -4840 11496 -4120
rect 12216 -4840 12256 -4120
rect 11456 -4880 12256 -4840
rect 12868 -4120 13668 -4080
rect 12868 -4840 12908 -4120
rect 13628 -4840 13668 -4120
rect 12868 -4880 13668 -4840
rect 14280 -4120 15080 -4080
rect 14280 -4840 14320 -4120
rect 15040 -4840 15080 -4120
rect 14280 -4880 15080 -4840
rect 15692 -4120 16492 -4080
rect 15692 -4840 15732 -4120
rect 16452 -4840 16492 -4120
rect 15692 -4880 16492 -4840
rect 17104 -4120 17904 -4080
rect 17104 -4840 17144 -4120
rect 17864 -4840 17904 -4120
rect 17104 -4880 17904 -4840
rect 18516 -4120 19316 -4080
rect 18516 -4840 18556 -4120
rect 19276 -4840 19316 -4120
rect 18516 -4880 19316 -4840
rect 19928 -4120 20728 -4080
rect 19928 -4840 19968 -4120
rect 20688 -4840 20728 -4120
rect 19928 -4880 20728 -4840
rect 21340 -4120 22140 -4080
rect 21340 -4840 21380 -4120
rect 22100 -4840 22140 -4120
rect 21340 -4880 22140 -4840
rect 22752 -4120 23552 -4080
rect 22752 -4840 22792 -4120
rect 23512 -4840 23552 -4120
rect 22752 -4880 23552 -4840
rect -23844 -5240 -23044 -5200
rect -23844 -5960 -23804 -5240
rect -23084 -5960 -23044 -5240
rect -23844 -6000 -23044 -5960
rect -22432 -5240 -21632 -5200
rect -22432 -5960 -22392 -5240
rect -21672 -5960 -21632 -5240
rect -22432 -6000 -21632 -5960
rect -21020 -5240 -20220 -5200
rect -21020 -5960 -20980 -5240
rect -20260 -5960 -20220 -5240
rect -21020 -6000 -20220 -5960
rect -19608 -5240 -18808 -5200
rect -19608 -5960 -19568 -5240
rect -18848 -5960 -18808 -5240
rect -19608 -6000 -18808 -5960
rect -18196 -5240 -17396 -5200
rect -18196 -5960 -18156 -5240
rect -17436 -5960 -17396 -5240
rect -18196 -6000 -17396 -5960
rect -16784 -5240 -15984 -5200
rect -16784 -5960 -16744 -5240
rect -16024 -5960 -15984 -5240
rect -16784 -6000 -15984 -5960
rect -15372 -5240 -14572 -5200
rect -15372 -5960 -15332 -5240
rect -14612 -5960 -14572 -5240
rect -15372 -6000 -14572 -5960
rect -13960 -5240 -13160 -5200
rect -13960 -5960 -13920 -5240
rect -13200 -5960 -13160 -5240
rect -13960 -6000 -13160 -5960
rect -12548 -5240 -11748 -5200
rect -12548 -5960 -12508 -5240
rect -11788 -5960 -11748 -5240
rect -12548 -6000 -11748 -5960
rect -11136 -5240 -10336 -5200
rect -11136 -5960 -11096 -5240
rect -10376 -5960 -10336 -5240
rect -11136 -6000 -10336 -5960
rect -9724 -5240 -8924 -5200
rect -9724 -5960 -9684 -5240
rect -8964 -5960 -8924 -5240
rect -9724 -6000 -8924 -5960
rect -8312 -5240 -7512 -5200
rect -8312 -5960 -8272 -5240
rect -7552 -5960 -7512 -5240
rect -8312 -6000 -7512 -5960
rect -6900 -5240 -6100 -5200
rect -6900 -5960 -6860 -5240
rect -6140 -5960 -6100 -5240
rect -6900 -6000 -6100 -5960
rect -5488 -5240 -4688 -5200
rect -5488 -5960 -5448 -5240
rect -4728 -5960 -4688 -5240
rect -5488 -6000 -4688 -5960
rect -4076 -5240 -3276 -5200
rect -4076 -5960 -4036 -5240
rect -3316 -5960 -3276 -5240
rect -4076 -6000 -3276 -5960
rect -2664 -5240 -1864 -5200
rect -2664 -5960 -2624 -5240
rect -1904 -5960 -1864 -5240
rect -2664 -6000 -1864 -5960
rect -1252 -5240 -452 -5200
rect -1252 -5960 -1212 -5240
rect -492 -5960 -452 -5240
rect -1252 -6000 -452 -5960
rect 160 -5240 960 -5200
rect 160 -5960 200 -5240
rect 920 -5960 960 -5240
rect 160 -6000 960 -5960
rect 1572 -5240 2372 -5200
rect 1572 -5960 1612 -5240
rect 2332 -5960 2372 -5240
rect 1572 -6000 2372 -5960
rect 2984 -5240 3784 -5200
rect 2984 -5960 3024 -5240
rect 3744 -5960 3784 -5240
rect 2984 -6000 3784 -5960
rect 4396 -5240 5196 -5200
rect 4396 -5960 4436 -5240
rect 5156 -5960 5196 -5240
rect 4396 -6000 5196 -5960
rect 5808 -5240 6608 -5200
rect 5808 -5960 5848 -5240
rect 6568 -5960 6608 -5240
rect 5808 -6000 6608 -5960
rect 7220 -5240 8020 -5200
rect 7220 -5960 7260 -5240
rect 7980 -5960 8020 -5240
rect 7220 -6000 8020 -5960
rect 8632 -5240 9432 -5200
rect 8632 -5960 8672 -5240
rect 9392 -5960 9432 -5240
rect 8632 -6000 9432 -5960
rect 10044 -5240 10844 -5200
rect 10044 -5960 10084 -5240
rect 10804 -5960 10844 -5240
rect 10044 -6000 10844 -5960
rect 11456 -5240 12256 -5200
rect 11456 -5960 11496 -5240
rect 12216 -5960 12256 -5240
rect 11456 -6000 12256 -5960
rect 12868 -5240 13668 -5200
rect 12868 -5960 12908 -5240
rect 13628 -5960 13668 -5240
rect 12868 -6000 13668 -5960
rect 14280 -5240 15080 -5200
rect 14280 -5960 14320 -5240
rect 15040 -5960 15080 -5240
rect 14280 -6000 15080 -5960
rect 15692 -5240 16492 -5200
rect 15692 -5960 15732 -5240
rect 16452 -5960 16492 -5240
rect 15692 -6000 16492 -5960
rect 17104 -5240 17904 -5200
rect 17104 -5960 17144 -5240
rect 17864 -5960 17904 -5240
rect 17104 -6000 17904 -5960
rect 18516 -5240 19316 -5200
rect 18516 -5960 18556 -5240
rect 19276 -5960 19316 -5240
rect 18516 -6000 19316 -5960
rect 19928 -5240 20728 -5200
rect 19928 -5960 19968 -5240
rect 20688 -5960 20728 -5240
rect 19928 -6000 20728 -5960
rect 21340 -5240 22140 -5200
rect 21340 -5960 21380 -5240
rect 22100 -5960 22140 -5240
rect 21340 -6000 22140 -5960
rect 22752 -5240 23552 -5200
rect 22752 -5960 22792 -5240
rect 23512 -5960 23552 -5240
rect 22752 -6000 23552 -5960
rect -23844 -6360 -23044 -6320
rect -23844 -7080 -23804 -6360
rect -23084 -7080 -23044 -6360
rect -23844 -7120 -23044 -7080
rect -22432 -6360 -21632 -6320
rect -22432 -7080 -22392 -6360
rect -21672 -7080 -21632 -6360
rect -22432 -7120 -21632 -7080
rect -21020 -6360 -20220 -6320
rect -21020 -7080 -20980 -6360
rect -20260 -7080 -20220 -6360
rect -21020 -7120 -20220 -7080
rect -19608 -6360 -18808 -6320
rect -19608 -7080 -19568 -6360
rect -18848 -7080 -18808 -6360
rect -19608 -7120 -18808 -7080
rect -18196 -6360 -17396 -6320
rect -18196 -7080 -18156 -6360
rect -17436 -7080 -17396 -6360
rect -18196 -7120 -17396 -7080
rect -16784 -6360 -15984 -6320
rect -16784 -7080 -16744 -6360
rect -16024 -7080 -15984 -6360
rect -16784 -7120 -15984 -7080
rect -15372 -6360 -14572 -6320
rect -15372 -7080 -15332 -6360
rect -14612 -7080 -14572 -6360
rect -15372 -7120 -14572 -7080
rect -13960 -6360 -13160 -6320
rect -13960 -7080 -13920 -6360
rect -13200 -7080 -13160 -6360
rect -13960 -7120 -13160 -7080
rect -12548 -6360 -11748 -6320
rect -12548 -7080 -12508 -6360
rect -11788 -7080 -11748 -6360
rect -12548 -7120 -11748 -7080
rect -11136 -6360 -10336 -6320
rect -11136 -7080 -11096 -6360
rect -10376 -7080 -10336 -6360
rect -11136 -7120 -10336 -7080
rect -9724 -6360 -8924 -6320
rect -9724 -7080 -9684 -6360
rect -8964 -7080 -8924 -6360
rect -9724 -7120 -8924 -7080
rect -8312 -6360 -7512 -6320
rect -8312 -7080 -8272 -6360
rect -7552 -7080 -7512 -6360
rect -8312 -7120 -7512 -7080
rect -6900 -6360 -6100 -6320
rect -6900 -7080 -6860 -6360
rect -6140 -7080 -6100 -6360
rect -6900 -7120 -6100 -7080
rect -5488 -6360 -4688 -6320
rect -5488 -7080 -5448 -6360
rect -4728 -7080 -4688 -6360
rect -5488 -7120 -4688 -7080
rect -4076 -6360 -3276 -6320
rect -4076 -7080 -4036 -6360
rect -3316 -7080 -3276 -6360
rect -4076 -7120 -3276 -7080
rect -2664 -6360 -1864 -6320
rect -2664 -7080 -2624 -6360
rect -1904 -7080 -1864 -6360
rect -2664 -7120 -1864 -7080
rect -1252 -6360 -452 -6320
rect -1252 -7080 -1212 -6360
rect -492 -7080 -452 -6360
rect -1252 -7120 -452 -7080
rect 160 -6360 960 -6320
rect 160 -7080 200 -6360
rect 920 -7080 960 -6360
rect 160 -7120 960 -7080
rect 1572 -6360 2372 -6320
rect 1572 -7080 1612 -6360
rect 2332 -7080 2372 -6360
rect 1572 -7120 2372 -7080
rect 2984 -6360 3784 -6320
rect 2984 -7080 3024 -6360
rect 3744 -7080 3784 -6360
rect 2984 -7120 3784 -7080
rect 4396 -6360 5196 -6320
rect 4396 -7080 4436 -6360
rect 5156 -7080 5196 -6360
rect 4396 -7120 5196 -7080
rect 5808 -6360 6608 -6320
rect 5808 -7080 5848 -6360
rect 6568 -7080 6608 -6360
rect 5808 -7120 6608 -7080
rect 7220 -6360 8020 -6320
rect 7220 -7080 7260 -6360
rect 7980 -7080 8020 -6360
rect 7220 -7120 8020 -7080
rect 8632 -6360 9432 -6320
rect 8632 -7080 8672 -6360
rect 9392 -7080 9432 -6360
rect 8632 -7120 9432 -7080
rect 10044 -6360 10844 -6320
rect 10044 -7080 10084 -6360
rect 10804 -7080 10844 -6360
rect 10044 -7120 10844 -7080
rect 11456 -6360 12256 -6320
rect 11456 -7080 11496 -6360
rect 12216 -7080 12256 -6360
rect 11456 -7120 12256 -7080
rect 12868 -6360 13668 -6320
rect 12868 -7080 12908 -6360
rect 13628 -7080 13668 -6360
rect 12868 -7120 13668 -7080
rect 14280 -6360 15080 -6320
rect 14280 -7080 14320 -6360
rect 15040 -7080 15080 -6360
rect 14280 -7120 15080 -7080
rect 15692 -6360 16492 -6320
rect 15692 -7080 15732 -6360
rect 16452 -7080 16492 -6360
rect 15692 -7120 16492 -7080
rect 17104 -6360 17904 -6320
rect 17104 -7080 17144 -6360
rect 17864 -7080 17904 -6360
rect 17104 -7120 17904 -7080
rect 18516 -6360 19316 -6320
rect 18516 -7080 18556 -6360
rect 19276 -7080 19316 -6360
rect 18516 -7120 19316 -7080
rect 19928 -6360 20728 -6320
rect 19928 -7080 19968 -6360
rect 20688 -7080 20728 -6360
rect 19928 -7120 20728 -7080
rect 21340 -6360 22140 -6320
rect 21340 -7080 21380 -6360
rect 22100 -7080 22140 -6360
rect 21340 -7120 22140 -7080
rect 22752 -6360 23552 -6320
rect 22752 -7080 22792 -6360
rect 23512 -7080 23552 -6360
rect 22752 -7120 23552 -7080
rect -23844 -7480 -23044 -7440
rect -23844 -8200 -23804 -7480
rect -23084 -8200 -23044 -7480
rect -23844 -8240 -23044 -8200
rect -22432 -7480 -21632 -7440
rect -22432 -8200 -22392 -7480
rect -21672 -8200 -21632 -7480
rect -22432 -8240 -21632 -8200
rect -21020 -7480 -20220 -7440
rect -21020 -8200 -20980 -7480
rect -20260 -8200 -20220 -7480
rect -21020 -8240 -20220 -8200
rect -19608 -7480 -18808 -7440
rect -19608 -8200 -19568 -7480
rect -18848 -8200 -18808 -7480
rect -19608 -8240 -18808 -8200
rect -18196 -7480 -17396 -7440
rect -18196 -8200 -18156 -7480
rect -17436 -8200 -17396 -7480
rect -18196 -8240 -17396 -8200
rect -16784 -7480 -15984 -7440
rect -16784 -8200 -16744 -7480
rect -16024 -8200 -15984 -7480
rect -16784 -8240 -15984 -8200
rect -15372 -7480 -14572 -7440
rect -15372 -8200 -15332 -7480
rect -14612 -8200 -14572 -7480
rect -15372 -8240 -14572 -8200
rect -13960 -7480 -13160 -7440
rect -13960 -8200 -13920 -7480
rect -13200 -8200 -13160 -7480
rect -13960 -8240 -13160 -8200
rect -12548 -7480 -11748 -7440
rect -12548 -8200 -12508 -7480
rect -11788 -8200 -11748 -7480
rect -12548 -8240 -11748 -8200
rect -11136 -7480 -10336 -7440
rect -11136 -8200 -11096 -7480
rect -10376 -8200 -10336 -7480
rect -11136 -8240 -10336 -8200
rect -9724 -7480 -8924 -7440
rect -9724 -8200 -9684 -7480
rect -8964 -8200 -8924 -7480
rect -9724 -8240 -8924 -8200
rect -8312 -7480 -7512 -7440
rect -8312 -8200 -8272 -7480
rect -7552 -8200 -7512 -7480
rect -8312 -8240 -7512 -8200
rect -6900 -7480 -6100 -7440
rect -6900 -8200 -6860 -7480
rect -6140 -8200 -6100 -7480
rect -6900 -8240 -6100 -8200
rect -5488 -7480 -4688 -7440
rect -5488 -8200 -5448 -7480
rect -4728 -8200 -4688 -7480
rect -5488 -8240 -4688 -8200
rect -4076 -7480 -3276 -7440
rect -4076 -8200 -4036 -7480
rect -3316 -8200 -3276 -7480
rect -4076 -8240 -3276 -8200
rect -2664 -7480 -1864 -7440
rect -2664 -8200 -2624 -7480
rect -1904 -8200 -1864 -7480
rect -2664 -8240 -1864 -8200
rect -1252 -7480 -452 -7440
rect -1252 -8200 -1212 -7480
rect -492 -8200 -452 -7480
rect -1252 -8240 -452 -8200
rect 160 -7480 960 -7440
rect 160 -8200 200 -7480
rect 920 -8200 960 -7480
rect 160 -8240 960 -8200
rect 1572 -7480 2372 -7440
rect 1572 -8200 1612 -7480
rect 2332 -8200 2372 -7480
rect 1572 -8240 2372 -8200
rect 2984 -7480 3784 -7440
rect 2984 -8200 3024 -7480
rect 3744 -8200 3784 -7480
rect 2984 -8240 3784 -8200
rect 4396 -7480 5196 -7440
rect 4396 -8200 4436 -7480
rect 5156 -8200 5196 -7480
rect 4396 -8240 5196 -8200
rect 5808 -7480 6608 -7440
rect 5808 -8200 5848 -7480
rect 6568 -8200 6608 -7480
rect 5808 -8240 6608 -8200
rect 7220 -7480 8020 -7440
rect 7220 -8200 7260 -7480
rect 7980 -8200 8020 -7480
rect 7220 -8240 8020 -8200
rect 8632 -7480 9432 -7440
rect 8632 -8200 8672 -7480
rect 9392 -8200 9432 -7480
rect 8632 -8240 9432 -8200
rect 10044 -7480 10844 -7440
rect 10044 -8200 10084 -7480
rect 10804 -8200 10844 -7480
rect 10044 -8240 10844 -8200
rect 11456 -7480 12256 -7440
rect 11456 -8200 11496 -7480
rect 12216 -8200 12256 -7480
rect 11456 -8240 12256 -8200
rect 12868 -7480 13668 -7440
rect 12868 -8200 12908 -7480
rect 13628 -8200 13668 -7480
rect 12868 -8240 13668 -8200
rect 14280 -7480 15080 -7440
rect 14280 -8200 14320 -7480
rect 15040 -8200 15080 -7480
rect 14280 -8240 15080 -8200
rect 15692 -7480 16492 -7440
rect 15692 -8200 15732 -7480
rect 16452 -8200 16492 -7480
rect 15692 -8240 16492 -8200
rect 17104 -7480 17904 -7440
rect 17104 -8200 17144 -7480
rect 17864 -8200 17904 -7480
rect 17104 -8240 17904 -8200
rect 18516 -7480 19316 -7440
rect 18516 -8200 18556 -7480
rect 19276 -8200 19316 -7480
rect 18516 -8240 19316 -8200
rect 19928 -7480 20728 -7440
rect 19928 -8200 19968 -7480
rect 20688 -8200 20728 -7480
rect 19928 -8240 20728 -8200
rect 21340 -7480 22140 -7440
rect 21340 -8200 21380 -7480
rect 22100 -8200 22140 -7480
rect 21340 -8240 22140 -8200
rect 22752 -7480 23552 -7440
rect 22752 -8200 22792 -7480
rect 23512 -8200 23552 -7480
rect 22752 -8240 23552 -8200
rect -23844 -8600 -23044 -8560
rect -23844 -9320 -23804 -8600
rect -23084 -9320 -23044 -8600
rect -23844 -9360 -23044 -9320
rect -22432 -8600 -21632 -8560
rect -22432 -9320 -22392 -8600
rect -21672 -9320 -21632 -8600
rect -22432 -9360 -21632 -9320
rect -21020 -8600 -20220 -8560
rect -21020 -9320 -20980 -8600
rect -20260 -9320 -20220 -8600
rect -21020 -9360 -20220 -9320
rect -19608 -8600 -18808 -8560
rect -19608 -9320 -19568 -8600
rect -18848 -9320 -18808 -8600
rect -19608 -9360 -18808 -9320
rect -18196 -8600 -17396 -8560
rect -18196 -9320 -18156 -8600
rect -17436 -9320 -17396 -8600
rect -18196 -9360 -17396 -9320
rect -16784 -8600 -15984 -8560
rect -16784 -9320 -16744 -8600
rect -16024 -9320 -15984 -8600
rect -16784 -9360 -15984 -9320
rect -15372 -8600 -14572 -8560
rect -15372 -9320 -15332 -8600
rect -14612 -9320 -14572 -8600
rect -15372 -9360 -14572 -9320
rect -13960 -8600 -13160 -8560
rect -13960 -9320 -13920 -8600
rect -13200 -9320 -13160 -8600
rect -13960 -9360 -13160 -9320
rect -12548 -8600 -11748 -8560
rect -12548 -9320 -12508 -8600
rect -11788 -9320 -11748 -8600
rect -12548 -9360 -11748 -9320
rect -11136 -8600 -10336 -8560
rect -11136 -9320 -11096 -8600
rect -10376 -9320 -10336 -8600
rect -11136 -9360 -10336 -9320
rect -9724 -8600 -8924 -8560
rect -9724 -9320 -9684 -8600
rect -8964 -9320 -8924 -8600
rect -9724 -9360 -8924 -9320
rect -8312 -8600 -7512 -8560
rect -8312 -9320 -8272 -8600
rect -7552 -9320 -7512 -8600
rect -8312 -9360 -7512 -9320
rect -6900 -8600 -6100 -8560
rect -6900 -9320 -6860 -8600
rect -6140 -9320 -6100 -8600
rect -6900 -9360 -6100 -9320
rect -5488 -8600 -4688 -8560
rect -5488 -9320 -5448 -8600
rect -4728 -9320 -4688 -8600
rect -5488 -9360 -4688 -9320
rect -4076 -8600 -3276 -8560
rect -4076 -9320 -4036 -8600
rect -3316 -9320 -3276 -8600
rect -4076 -9360 -3276 -9320
rect -2664 -8600 -1864 -8560
rect -2664 -9320 -2624 -8600
rect -1904 -9320 -1864 -8600
rect -2664 -9360 -1864 -9320
rect -1252 -8600 -452 -8560
rect -1252 -9320 -1212 -8600
rect -492 -9320 -452 -8600
rect -1252 -9360 -452 -9320
rect 160 -8600 960 -8560
rect 160 -9320 200 -8600
rect 920 -9320 960 -8600
rect 160 -9360 960 -9320
rect 1572 -8600 2372 -8560
rect 1572 -9320 1612 -8600
rect 2332 -9320 2372 -8600
rect 1572 -9360 2372 -9320
rect 2984 -8600 3784 -8560
rect 2984 -9320 3024 -8600
rect 3744 -9320 3784 -8600
rect 2984 -9360 3784 -9320
rect 4396 -8600 5196 -8560
rect 4396 -9320 4436 -8600
rect 5156 -9320 5196 -8600
rect 4396 -9360 5196 -9320
rect 5808 -8600 6608 -8560
rect 5808 -9320 5848 -8600
rect 6568 -9320 6608 -8600
rect 5808 -9360 6608 -9320
rect 7220 -8600 8020 -8560
rect 7220 -9320 7260 -8600
rect 7980 -9320 8020 -8600
rect 7220 -9360 8020 -9320
rect 8632 -8600 9432 -8560
rect 8632 -9320 8672 -8600
rect 9392 -9320 9432 -8600
rect 8632 -9360 9432 -9320
rect 10044 -8600 10844 -8560
rect 10044 -9320 10084 -8600
rect 10804 -9320 10844 -8600
rect 10044 -9360 10844 -9320
rect 11456 -8600 12256 -8560
rect 11456 -9320 11496 -8600
rect 12216 -9320 12256 -8600
rect 11456 -9360 12256 -9320
rect 12868 -8600 13668 -8560
rect 12868 -9320 12908 -8600
rect 13628 -9320 13668 -8600
rect 12868 -9360 13668 -9320
rect 14280 -8600 15080 -8560
rect 14280 -9320 14320 -8600
rect 15040 -9320 15080 -8600
rect 14280 -9360 15080 -9320
rect 15692 -8600 16492 -8560
rect 15692 -9320 15732 -8600
rect 16452 -9320 16492 -8600
rect 15692 -9360 16492 -9320
rect 17104 -8600 17904 -8560
rect 17104 -9320 17144 -8600
rect 17864 -9320 17904 -8600
rect 17104 -9360 17904 -9320
rect 18516 -8600 19316 -8560
rect 18516 -9320 18556 -8600
rect 19276 -9320 19316 -8600
rect 18516 -9360 19316 -9320
rect 19928 -8600 20728 -8560
rect 19928 -9320 19968 -8600
rect 20688 -9320 20728 -8600
rect 19928 -9360 20728 -9320
rect 21340 -8600 22140 -8560
rect 21340 -9320 21380 -8600
rect 22100 -9320 22140 -8600
rect 21340 -9360 22140 -9320
rect 22752 -8600 23552 -8560
rect 22752 -9320 22792 -8600
rect 23512 -9320 23552 -8600
rect 22752 -9360 23552 -9320
rect -23844 -9720 -23044 -9680
rect -23844 -10440 -23804 -9720
rect -23084 -10440 -23044 -9720
rect -23844 -10480 -23044 -10440
rect -22432 -9720 -21632 -9680
rect -22432 -10440 -22392 -9720
rect -21672 -10440 -21632 -9720
rect -22432 -10480 -21632 -10440
rect -21020 -9720 -20220 -9680
rect -21020 -10440 -20980 -9720
rect -20260 -10440 -20220 -9720
rect -21020 -10480 -20220 -10440
rect -19608 -9720 -18808 -9680
rect -19608 -10440 -19568 -9720
rect -18848 -10440 -18808 -9720
rect -19608 -10480 -18808 -10440
rect -18196 -9720 -17396 -9680
rect -18196 -10440 -18156 -9720
rect -17436 -10440 -17396 -9720
rect -18196 -10480 -17396 -10440
rect -16784 -9720 -15984 -9680
rect -16784 -10440 -16744 -9720
rect -16024 -10440 -15984 -9720
rect -16784 -10480 -15984 -10440
rect -15372 -9720 -14572 -9680
rect -15372 -10440 -15332 -9720
rect -14612 -10440 -14572 -9720
rect -15372 -10480 -14572 -10440
rect -13960 -9720 -13160 -9680
rect -13960 -10440 -13920 -9720
rect -13200 -10440 -13160 -9720
rect -13960 -10480 -13160 -10440
rect -12548 -9720 -11748 -9680
rect -12548 -10440 -12508 -9720
rect -11788 -10440 -11748 -9720
rect -12548 -10480 -11748 -10440
rect -11136 -9720 -10336 -9680
rect -11136 -10440 -11096 -9720
rect -10376 -10440 -10336 -9720
rect -11136 -10480 -10336 -10440
rect -9724 -9720 -8924 -9680
rect -9724 -10440 -9684 -9720
rect -8964 -10440 -8924 -9720
rect -9724 -10480 -8924 -10440
rect -8312 -9720 -7512 -9680
rect -8312 -10440 -8272 -9720
rect -7552 -10440 -7512 -9720
rect -8312 -10480 -7512 -10440
rect -6900 -9720 -6100 -9680
rect -6900 -10440 -6860 -9720
rect -6140 -10440 -6100 -9720
rect -6900 -10480 -6100 -10440
rect -5488 -9720 -4688 -9680
rect -5488 -10440 -5448 -9720
rect -4728 -10440 -4688 -9720
rect -5488 -10480 -4688 -10440
rect -4076 -9720 -3276 -9680
rect -4076 -10440 -4036 -9720
rect -3316 -10440 -3276 -9720
rect -4076 -10480 -3276 -10440
rect -2664 -9720 -1864 -9680
rect -2664 -10440 -2624 -9720
rect -1904 -10440 -1864 -9720
rect -2664 -10480 -1864 -10440
rect -1252 -9720 -452 -9680
rect -1252 -10440 -1212 -9720
rect -492 -10440 -452 -9720
rect -1252 -10480 -452 -10440
rect 160 -9720 960 -9680
rect 160 -10440 200 -9720
rect 920 -10440 960 -9720
rect 160 -10480 960 -10440
rect 1572 -9720 2372 -9680
rect 1572 -10440 1612 -9720
rect 2332 -10440 2372 -9720
rect 1572 -10480 2372 -10440
rect 2984 -9720 3784 -9680
rect 2984 -10440 3024 -9720
rect 3744 -10440 3784 -9720
rect 2984 -10480 3784 -10440
rect 4396 -9720 5196 -9680
rect 4396 -10440 4436 -9720
rect 5156 -10440 5196 -9720
rect 4396 -10480 5196 -10440
rect 5808 -9720 6608 -9680
rect 5808 -10440 5848 -9720
rect 6568 -10440 6608 -9720
rect 5808 -10480 6608 -10440
rect 7220 -9720 8020 -9680
rect 7220 -10440 7260 -9720
rect 7980 -10440 8020 -9720
rect 7220 -10480 8020 -10440
rect 8632 -9720 9432 -9680
rect 8632 -10440 8672 -9720
rect 9392 -10440 9432 -9720
rect 8632 -10480 9432 -10440
rect 10044 -9720 10844 -9680
rect 10044 -10440 10084 -9720
rect 10804 -10440 10844 -9720
rect 10044 -10480 10844 -10440
rect 11456 -9720 12256 -9680
rect 11456 -10440 11496 -9720
rect 12216 -10440 12256 -9720
rect 11456 -10480 12256 -10440
rect 12868 -9720 13668 -9680
rect 12868 -10440 12908 -9720
rect 13628 -10440 13668 -9720
rect 12868 -10480 13668 -10440
rect 14280 -9720 15080 -9680
rect 14280 -10440 14320 -9720
rect 15040 -10440 15080 -9720
rect 14280 -10480 15080 -10440
rect 15692 -9720 16492 -9680
rect 15692 -10440 15732 -9720
rect 16452 -10440 16492 -9720
rect 15692 -10480 16492 -10440
rect 17104 -9720 17904 -9680
rect 17104 -10440 17144 -9720
rect 17864 -10440 17904 -9720
rect 17104 -10480 17904 -10440
rect 18516 -9720 19316 -9680
rect 18516 -10440 18556 -9720
rect 19276 -10440 19316 -9720
rect 18516 -10480 19316 -10440
rect 19928 -9720 20728 -9680
rect 19928 -10440 19968 -9720
rect 20688 -10440 20728 -9720
rect 19928 -10480 20728 -10440
rect 21340 -9720 22140 -9680
rect 21340 -10440 21380 -9720
rect 22100 -10440 22140 -9720
rect 21340 -10480 22140 -10440
rect 22752 -9720 23552 -9680
rect 22752 -10440 22792 -9720
rect 23512 -10440 23552 -9720
rect 22752 -10480 23552 -10440
rect -23844 -10840 -23044 -10800
rect -23844 -11560 -23804 -10840
rect -23084 -11560 -23044 -10840
rect -23844 -11600 -23044 -11560
rect -22432 -10840 -21632 -10800
rect -22432 -11560 -22392 -10840
rect -21672 -11560 -21632 -10840
rect -22432 -11600 -21632 -11560
rect -21020 -10840 -20220 -10800
rect -21020 -11560 -20980 -10840
rect -20260 -11560 -20220 -10840
rect -21020 -11600 -20220 -11560
rect -19608 -10840 -18808 -10800
rect -19608 -11560 -19568 -10840
rect -18848 -11560 -18808 -10840
rect -19608 -11600 -18808 -11560
rect -18196 -10840 -17396 -10800
rect -18196 -11560 -18156 -10840
rect -17436 -11560 -17396 -10840
rect -18196 -11600 -17396 -11560
rect -16784 -10840 -15984 -10800
rect -16784 -11560 -16744 -10840
rect -16024 -11560 -15984 -10840
rect -16784 -11600 -15984 -11560
rect -15372 -10840 -14572 -10800
rect -15372 -11560 -15332 -10840
rect -14612 -11560 -14572 -10840
rect -15372 -11600 -14572 -11560
rect -13960 -10840 -13160 -10800
rect -13960 -11560 -13920 -10840
rect -13200 -11560 -13160 -10840
rect -13960 -11600 -13160 -11560
rect -12548 -10840 -11748 -10800
rect -12548 -11560 -12508 -10840
rect -11788 -11560 -11748 -10840
rect -12548 -11600 -11748 -11560
rect -11136 -10840 -10336 -10800
rect -11136 -11560 -11096 -10840
rect -10376 -11560 -10336 -10840
rect -11136 -11600 -10336 -11560
rect -9724 -10840 -8924 -10800
rect -9724 -11560 -9684 -10840
rect -8964 -11560 -8924 -10840
rect -9724 -11600 -8924 -11560
rect -8312 -10840 -7512 -10800
rect -8312 -11560 -8272 -10840
rect -7552 -11560 -7512 -10840
rect -8312 -11600 -7512 -11560
rect -6900 -10840 -6100 -10800
rect -6900 -11560 -6860 -10840
rect -6140 -11560 -6100 -10840
rect -6900 -11600 -6100 -11560
rect -5488 -10840 -4688 -10800
rect -5488 -11560 -5448 -10840
rect -4728 -11560 -4688 -10840
rect -5488 -11600 -4688 -11560
rect -4076 -10840 -3276 -10800
rect -4076 -11560 -4036 -10840
rect -3316 -11560 -3276 -10840
rect -4076 -11600 -3276 -11560
rect -2664 -10840 -1864 -10800
rect -2664 -11560 -2624 -10840
rect -1904 -11560 -1864 -10840
rect -2664 -11600 -1864 -11560
rect -1252 -10840 -452 -10800
rect -1252 -11560 -1212 -10840
rect -492 -11560 -452 -10840
rect -1252 -11600 -452 -11560
rect 160 -10840 960 -10800
rect 160 -11560 200 -10840
rect 920 -11560 960 -10840
rect 160 -11600 960 -11560
rect 1572 -10840 2372 -10800
rect 1572 -11560 1612 -10840
rect 2332 -11560 2372 -10840
rect 1572 -11600 2372 -11560
rect 2984 -10840 3784 -10800
rect 2984 -11560 3024 -10840
rect 3744 -11560 3784 -10840
rect 2984 -11600 3784 -11560
rect 4396 -10840 5196 -10800
rect 4396 -11560 4436 -10840
rect 5156 -11560 5196 -10840
rect 4396 -11600 5196 -11560
rect 5808 -10840 6608 -10800
rect 5808 -11560 5848 -10840
rect 6568 -11560 6608 -10840
rect 5808 -11600 6608 -11560
rect 7220 -10840 8020 -10800
rect 7220 -11560 7260 -10840
rect 7980 -11560 8020 -10840
rect 7220 -11600 8020 -11560
rect 8632 -10840 9432 -10800
rect 8632 -11560 8672 -10840
rect 9392 -11560 9432 -10840
rect 8632 -11600 9432 -11560
rect 10044 -10840 10844 -10800
rect 10044 -11560 10084 -10840
rect 10804 -11560 10844 -10840
rect 10044 -11600 10844 -11560
rect 11456 -10840 12256 -10800
rect 11456 -11560 11496 -10840
rect 12216 -11560 12256 -10840
rect 11456 -11600 12256 -11560
rect 12868 -10840 13668 -10800
rect 12868 -11560 12908 -10840
rect 13628 -11560 13668 -10840
rect 12868 -11600 13668 -11560
rect 14280 -10840 15080 -10800
rect 14280 -11560 14320 -10840
rect 15040 -11560 15080 -10840
rect 14280 -11600 15080 -11560
rect 15692 -10840 16492 -10800
rect 15692 -11560 15732 -10840
rect 16452 -11560 16492 -10840
rect 15692 -11600 16492 -11560
rect 17104 -10840 17904 -10800
rect 17104 -11560 17144 -10840
rect 17864 -11560 17904 -10840
rect 17104 -11600 17904 -11560
rect 18516 -10840 19316 -10800
rect 18516 -11560 18556 -10840
rect 19276 -11560 19316 -10840
rect 18516 -11600 19316 -11560
rect 19928 -10840 20728 -10800
rect 19928 -11560 19968 -10840
rect 20688 -11560 20728 -10840
rect 19928 -11600 20728 -11560
rect 21340 -10840 22140 -10800
rect 21340 -11560 21380 -10840
rect 22100 -11560 22140 -10840
rect 21340 -11600 22140 -11560
rect 22752 -10840 23552 -10800
rect 22752 -11560 22792 -10840
rect 23512 -11560 23552 -10840
rect 22752 -11600 23552 -11560
rect -23844 -11960 -23044 -11920
rect -23844 -12680 -23804 -11960
rect -23084 -12680 -23044 -11960
rect -23844 -12720 -23044 -12680
rect -22432 -11960 -21632 -11920
rect -22432 -12680 -22392 -11960
rect -21672 -12680 -21632 -11960
rect -22432 -12720 -21632 -12680
rect -21020 -11960 -20220 -11920
rect -21020 -12680 -20980 -11960
rect -20260 -12680 -20220 -11960
rect -21020 -12720 -20220 -12680
rect -19608 -11960 -18808 -11920
rect -19608 -12680 -19568 -11960
rect -18848 -12680 -18808 -11960
rect -19608 -12720 -18808 -12680
rect -18196 -11960 -17396 -11920
rect -18196 -12680 -18156 -11960
rect -17436 -12680 -17396 -11960
rect -18196 -12720 -17396 -12680
rect -16784 -11960 -15984 -11920
rect -16784 -12680 -16744 -11960
rect -16024 -12680 -15984 -11960
rect -16784 -12720 -15984 -12680
rect -15372 -11960 -14572 -11920
rect -15372 -12680 -15332 -11960
rect -14612 -12680 -14572 -11960
rect -15372 -12720 -14572 -12680
rect -13960 -11960 -13160 -11920
rect -13960 -12680 -13920 -11960
rect -13200 -12680 -13160 -11960
rect -13960 -12720 -13160 -12680
rect -12548 -11960 -11748 -11920
rect -12548 -12680 -12508 -11960
rect -11788 -12680 -11748 -11960
rect -12548 -12720 -11748 -12680
rect -11136 -11960 -10336 -11920
rect -11136 -12680 -11096 -11960
rect -10376 -12680 -10336 -11960
rect -11136 -12720 -10336 -12680
rect -9724 -11960 -8924 -11920
rect -9724 -12680 -9684 -11960
rect -8964 -12680 -8924 -11960
rect -9724 -12720 -8924 -12680
rect -8312 -11960 -7512 -11920
rect -8312 -12680 -8272 -11960
rect -7552 -12680 -7512 -11960
rect -8312 -12720 -7512 -12680
rect -6900 -11960 -6100 -11920
rect -6900 -12680 -6860 -11960
rect -6140 -12680 -6100 -11960
rect -6900 -12720 -6100 -12680
rect -5488 -11960 -4688 -11920
rect -5488 -12680 -5448 -11960
rect -4728 -12680 -4688 -11960
rect -5488 -12720 -4688 -12680
rect -4076 -11960 -3276 -11920
rect -4076 -12680 -4036 -11960
rect -3316 -12680 -3276 -11960
rect -4076 -12720 -3276 -12680
rect -2664 -11960 -1864 -11920
rect -2664 -12680 -2624 -11960
rect -1904 -12680 -1864 -11960
rect -2664 -12720 -1864 -12680
rect -1252 -11960 -452 -11920
rect -1252 -12680 -1212 -11960
rect -492 -12680 -452 -11960
rect -1252 -12720 -452 -12680
rect 160 -11960 960 -11920
rect 160 -12680 200 -11960
rect 920 -12680 960 -11960
rect 160 -12720 960 -12680
rect 1572 -11960 2372 -11920
rect 1572 -12680 1612 -11960
rect 2332 -12680 2372 -11960
rect 1572 -12720 2372 -12680
rect 2984 -11960 3784 -11920
rect 2984 -12680 3024 -11960
rect 3744 -12680 3784 -11960
rect 2984 -12720 3784 -12680
rect 4396 -11960 5196 -11920
rect 4396 -12680 4436 -11960
rect 5156 -12680 5196 -11960
rect 4396 -12720 5196 -12680
rect 5808 -11960 6608 -11920
rect 5808 -12680 5848 -11960
rect 6568 -12680 6608 -11960
rect 5808 -12720 6608 -12680
rect 7220 -11960 8020 -11920
rect 7220 -12680 7260 -11960
rect 7980 -12680 8020 -11960
rect 7220 -12720 8020 -12680
rect 8632 -11960 9432 -11920
rect 8632 -12680 8672 -11960
rect 9392 -12680 9432 -11960
rect 8632 -12720 9432 -12680
rect 10044 -11960 10844 -11920
rect 10044 -12680 10084 -11960
rect 10804 -12680 10844 -11960
rect 10044 -12720 10844 -12680
rect 11456 -11960 12256 -11920
rect 11456 -12680 11496 -11960
rect 12216 -12680 12256 -11960
rect 11456 -12720 12256 -12680
rect 12868 -11960 13668 -11920
rect 12868 -12680 12908 -11960
rect 13628 -12680 13668 -11960
rect 12868 -12720 13668 -12680
rect 14280 -11960 15080 -11920
rect 14280 -12680 14320 -11960
rect 15040 -12680 15080 -11960
rect 14280 -12720 15080 -12680
rect 15692 -11960 16492 -11920
rect 15692 -12680 15732 -11960
rect 16452 -12680 16492 -11960
rect 15692 -12720 16492 -12680
rect 17104 -11960 17904 -11920
rect 17104 -12680 17144 -11960
rect 17864 -12680 17904 -11960
rect 17104 -12720 17904 -12680
rect 18516 -11960 19316 -11920
rect 18516 -12680 18556 -11960
rect 19276 -12680 19316 -11960
rect 18516 -12720 19316 -12680
rect 19928 -11960 20728 -11920
rect 19928 -12680 19968 -11960
rect 20688 -12680 20728 -11960
rect 19928 -12720 20728 -12680
rect 21340 -11960 22140 -11920
rect 21340 -12680 21380 -11960
rect 22100 -12680 22140 -11960
rect 21340 -12720 22140 -12680
rect 22752 -11960 23552 -11920
rect 22752 -12680 22792 -11960
rect 23512 -12680 23552 -11960
rect 22752 -12720 23552 -12680
rect -23844 -13080 -23044 -13040
rect -23844 -13800 -23804 -13080
rect -23084 -13800 -23044 -13080
rect -23844 -13840 -23044 -13800
rect -22432 -13080 -21632 -13040
rect -22432 -13800 -22392 -13080
rect -21672 -13800 -21632 -13080
rect -22432 -13840 -21632 -13800
rect -21020 -13080 -20220 -13040
rect -21020 -13800 -20980 -13080
rect -20260 -13800 -20220 -13080
rect -21020 -13840 -20220 -13800
rect -19608 -13080 -18808 -13040
rect -19608 -13800 -19568 -13080
rect -18848 -13800 -18808 -13080
rect -19608 -13840 -18808 -13800
rect -18196 -13080 -17396 -13040
rect -18196 -13800 -18156 -13080
rect -17436 -13800 -17396 -13080
rect -18196 -13840 -17396 -13800
rect -16784 -13080 -15984 -13040
rect -16784 -13800 -16744 -13080
rect -16024 -13800 -15984 -13080
rect -16784 -13840 -15984 -13800
rect -15372 -13080 -14572 -13040
rect -15372 -13800 -15332 -13080
rect -14612 -13800 -14572 -13080
rect -15372 -13840 -14572 -13800
rect -13960 -13080 -13160 -13040
rect -13960 -13800 -13920 -13080
rect -13200 -13800 -13160 -13080
rect -13960 -13840 -13160 -13800
rect -12548 -13080 -11748 -13040
rect -12548 -13800 -12508 -13080
rect -11788 -13800 -11748 -13080
rect -12548 -13840 -11748 -13800
rect -11136 -13080 -10336 -13040
rect -11136 -13800 -11096 -13080
rect -10376 -13800 -10336 -13080
rect -11136 -13840 -10336 -13800
rect -9724 -13080 -8924 -13040
rect -9724 -13800 -9684 -13080
rect -8964 -13800 -8924 -13080
rect -9724 -13840 -8924 -13800
rect -8312 -13080 -7512 -13040
rect -8312 -13800 -8272 -13080
rect -7552 -13800 -7512 -13080
rect -8312 -13840 -7512 -13800
rect -6900 -13080 -6100 -13040
rect -6900 -13800 -6860 -13080
rect -6140 -13800 -6100 -13080
rect -6900 -13840 -6100 -13800
rect -5488 -13080 -4688 -13040
rect -5488 -13800 -5448 -13080
rect -4728 -13800 -4688 -13080
rect -5488 -13840 -4688 -13800
rect -4076 -13080 -3276 -13040
rect -4076 -13800 -4036 -13080
rect -3316 -13800 -3276 -13080
rect -4076 -13840 -3276 -13800
rect -2664 -13080 -1864 -13040
rect -2664 -13800 -2624 -13080
rect -1904 -13800 -1864 -13080
rect -2664 -13840 -1864 -13800
rect -1252 -13080 -452 -13040
rect -1252 -13800 -1212 -13080
rect -492 -13800 -452 -13080
rect -1252 -13840 -452 -13800
rect 160 -13080 960 -13040
rect 160 -13800 200 -13080
rect 920 -13800 960 -13080
rect 160 -13840 960 -13800
rect 1572 -13080 2372 -13040
rect 1572 -13800 1612 -13080
rect 2332 -13800 2372 -13080
rect 1572 -13840 2372 -13800
rect 2984 -13080 3784 -13040
rect 2984 -13800 3024 -13080
rect 3744 -13800 3784 -13080
rect 2984 -13840 3784 -13800
rect 4396 -13080 5196 -13040
rect 4396 -13800 4436 -13080
rect 5156 -13800 5196 -13080
rect 4396 -13840 5196 -13800
rect 5808 -13080 6608 -13040
rect 5808 -13800 5848 -13080
rect 6568 -13800 6608 -13080
rect 5808 -13840 6608 -13800
rect 7220 -13080 8020 -13040
rect 7220 -13800 7260 -13080
rect 7980 -13800 8020 -13080
rect 7220 -13840 8020 -13800
rect 8632 -13080 9432 -13040
rect 8632 -13800 8672 -13080
rect 9392 -13800 9432 -13080
rect 8632 -13840 9432 -13800
rect 10044 -13080 10844 -13040
rect 10044 -13800 10084 -13080
rect 10804 -13800 10844 -13080
rect 10044 -13840 10844 -13800
rect 11456 -13080 12256 -13040
rect 11456 -13800 11496 -13080
rect 12216 -13800 12256 -13080
rect 11456 -13840 12256 -13800
rect 12868 -13080 13668 -13040
rect 12868 -13800 12908 -13080
rect 13628 -13800 13668 -13080
rect 12868 -13840 13668 -13800
rect 14280 -13080 15080 -13040
rect 14280 -13800 14320 -13080
rect 15040 -13800 15080 -13080
rect 14280 -13840 15080 -13800
rect 15692 -13080 16492 -13040
rect 15692 -13800 15732 -13080
rect 16452 -13800 16492 -13080
rect 15692 -13840 16492 -13800
rect 17104 -13080 17904 -13040
rect 17104 -13800 17144 -13080
rect 17864 -13800 17904 -13080
rect 17104 -13840 17904 -13800
rect 18516 -13080 19316 -13040
rect 18516 -13800 18556 -13080
rect 19276 -13800 19316 -13080
rect 18516 -13840 19316 -13800
rect 19928 -13080 20728 -13040
rect 19928 -13800 19968 -13080
rect 20688 -13800 20728 -13080
rect 19928 -13840 20728 -13800
rect 21340 -13080 22140 -13040
rect 21340 -13800 21380 -13080
rect 22100 -13800 22140 -13080
rect 21340 -13840 22140 -13800
rect 22752 -13080 23552 -13040
rect 22752 -13800 22792 -13080
rect 23512 -13800 23552 -13080
rect 22752 -13840 23552 -13800
rect -23844 -14200 -23044 -14160
rect -23844 -14920 -23804 -14200
rect -23084 -14920 -23044 -14200
rect -23844 -14960 -23044 -14920
rect -22432 -14200 -21632 -14160
rect -22432 -14920 -22392 -14200
rect -21672 -14920 -21632 -14200
rect -22432 -14960 -21632 -14920
rect -21020 -14200 -20220 -14160
rect -21020 -14920 -20980 -14200
rect -20260 -14920 -20220 -14200
rect -21020 -14960 -20220 -14920
rect -19608 -14200 -18808 -14160
rect -19608 -14920 -19568 -14200
rect -18848 -14920 -18808 -14200
rect -19608 -14960 -18808 -14920
rect -18196 -14200 -17396 -14160
rect -18196 -14920 -18156 -14200
rect -17436 -14920 -17396 -14200
rect -18196 -14960 -17396 -14920
rect -16784 -14200 -15984 -14160
rect -16784 -14920 -16744 -14200
rect -16024 -14920 -15984 -14200
rect -16784 -14960 -15984 -14920
rect -15372 -14200 -14572 -14160
rect -15372 -14920 -15332 -14200
rect -14612 -14920 -14572 -14200
rect -15372 -14960 -14572 -14920
rect -13960 -14200 -13160 -14160
rect -13960 -14920 -13920 -14200
rect -13200 -14920 -13160 -14200
rect -13960 -14960 -13160 -14920
rect -12548 -14200 -11748 -14160
rect -12548 -14920 -12508 -14200
rect -11788 -14920 -11748 -14200
rect -12548 -14960 -11748 -14920
rect -11136 -14200 -10336 -14160
rect -11136 -14920 -11096 -14200
rect -10376 -14920 -10336 -14200
rect -11136 -14960 -10336 -14920
rect -9724 -14200 -8924 -14160
rect -9724 -14920 -9684 -14200
rect -8964 -14920 -8924 -14200
rect -9724 -14960 -8924 -14920
rect -8312 -14200 -7512 -14160
rect -8312 -14920 -8272 -14200
rect -7552 -14920 -7512 -14200
rect -8312 -14960 -7512 -14920
rect -6900 -14200 -6100 -14160
rect -6900 -14920 -6860 -14200
rect -6140 -14920 -6100 -14200
rect -6900 -14960 -6100 -14920
rect -5488 -14200 -4688 -14160
rect -5488 -14920 -5448 -14200
rect -4728 -14920 -4688 -14200
rect -5488 -14960 -4688 -14920
rect -4076 -14200 -3276 -14160
rect -4076 -14920 -4036 -14200
rect -3316 -14920 -3276 -14200
rect -4076 -14960 -3276 -14920
rect -2664 -14200 -1864 -14160
rect -2664 -14920 -2624 -14200
rect -1904 -14920 -1864 -14200
rect -2664 -14960 -1864 -14920
rect -1252 -14200 -452 -14160
rect -1252 -14920 -1212 -14200
rect -492 -14920 -452 -14200
rect -1252 -14960 -452 -14920
rect 160 -14200 960 -14160
rect 160 -14920 200 -14200
rect 920 -14920 960 -14200
rect 160 -14960 960 -14920
rect 1572 -14200 2372 -14160
rect 1572 -14920 1612 -14200
rect 2332 -14920 2372 -14200
rect 1572 -14960 2372 -14920
rect 2984 -14200 3784 -14160
rect 2984 -14920 3024 -14200
rect 3744 -14920 3784 -14200
rect 2984 -14960 3784 -14920
rect 4396 -14200 5196 -14160
rect 4396 -14920 4436 -14200
rect 5156 -14920 5196 -14200
rect 4396 -14960 5196 -14920
rect 5808 -14200 6608 -14160
rect 5808 -14920 5848 -14200
rect 6568 -14920 6608 -14200
rect 5808 -14960 6608 -14920
rect 7220 -14200 8020 -14160
rect 7220 -14920 7260 -14200
rect 7980 -14920 8020 -14200
rect 7220 -14960 8020 -14920
rect 8632 -14200 9432 -14160
rect 8632 -14920 8672 -14200
rect 9392 -14920 9432 -14200
rect 8632 -14960 9432 -14920
rect 10044 -14200 10844 -14160
rect 10044 -14920 10084 -14200
rect 10804 -14920 10844 -14200
rect 10044 -14960 10844 -14920
rect 11456 -14200 12256 -14160
rect 11456 -14920 11496 -14200
rect 12216 -14920 12256 -14200
rect 11456 -14960 12256 -14920
rect 12868 -14200 13668 -14160
rect 12868 -14920 12908 -14200
rect 13628 -14920 13668 -14200
rect 12868 -14960 13668 -14920
rect 14280 -14200 15080 -14160
rect 14280 -14920 14320 -14200
rect 15040 -14920 15080 -14200
rect 14280 -14960 15080 -14920
rect 15692 -14200 16492 -14160
rect 15692 -14920 15732 -14200
rect 16452 -14920 16492 -14200
rect 15692 -14960 16492 -14920
rect 17104 -14200 17904 -14160
rect 17104 -14920 17144 -14200
rect 17864 -14920 17904 -14200
rect 17104 -14960 17904 -14920
rect 18516 -14200 19316 -14160
rect 18516 -14920 18556 -14200
rect 19276 -14920 19316 -14200
rect 18516 -14960 19316 -14920
rect 19928 -14200 20728 -14160
rect 19928 -14920 19968 -14200
rect 20688 -14920 20728 -14200
rect 19928 -14960 20728 -14920
rect 21340 -14200 22140 -14160
rect 21340 -14920 21380 -14200
rect 22100 -14920 22140 -14200
rect 21340 -14960 22140 -14920
rect 22752 -14200 23552 -14160
rect 22752 -14920 22792 -14200
rect 23512 -14920 23552 -14200
rect 22752 -14960 23552 -14920
rect -23844 -15320 -23044 -15280
rect -23844 -16040 -23804 -15320
rect -23084 -16040 -23044 -15320
rect -23844 -16080 -23044 -16040
rect -22432 -15320 -21632 -15280
rect -22432 -16040 -22392 -15320
rect -21672 -16040 -21632 -15320
rect -22432 -16080 -21632 -16040
rect -21020 -15320 -20220 -15280
rect -21020 -16040 -20980 -15320
rect -20260 -16040 -20220 -15320
rect -21020 -16080 -20220 -16040
rect -19608 -15320 -18808 -15280
rect -19608 -16040 -19568 -15320
rect -18848 -16040 -18808 -15320
rect -19608 -16080 -18808 -16040
rect -18196 -15320 -17396 -15280
rect -18196 -16040 -18156 -15320
rect -17436 -16040 -17396 -15320
rect -18196 -16080 -17396 -16040
rect -16784 -15320 -15984 -15280
rect -16784 -16040 -16744 -15320
rect -16024 -16040 -15984 -15320
rect -16784 -16080 -15984 -16040
rect -15372 -15320 -14572 -15280
rect -15372 -16040 -15332 -15320
rect -14612 -16040 -14572 -15320
rect -15372 -16080 -14572 -16040
rect -13960 -15320 -13160 -15280
rect -13960 -16040 -13920 -15320
rect -13200 -16040 -13160 -15320
rect -13960 -16080 -13160 -16040
rect -12548 -15320 -11748 -15280
rect -12548 -16040 -12508 -15320
rect -11788 -16040 -11748 -15320
rect -12548 -16080 -11748 -16040
rect -11136 -15320 -10336 -15280
rect -11136 -16040 -11096 -15320
rect -10376 -16040 -10336 -15320
rect -11136 -16080 -10336 -16040
rect -9724 -15320 -8924 -15280
rect -9724 -16040 -9684 -15320
rect -8964 -16040 -8924 -15320
rect -9724 -16080 -8924 -16040
rect -8312 -15320 -7512 -15280
rect -8312 -16040 -8272 -15320
rect -7552 -16040 -7512 -15320
rect -8312 -16080 -7512 -16040
rect -6900 -15320 -6100 -15280
rect -6900 -16040 -6860 -15320
rect -6140 -16040 -6100 -15320
rect -6900 -16080 -6100 -16040
rect -5488 -15320 -4688 -15280
rect -5488 -16040 -5448 -15320
rect -4728 -16040 -4688 -15320
rect -5488 -16080 -4688 -16040
rect -4076 -15320 -3276 -15280
rect -4076 -16040 -4036 -15320
rect -3316 -16040 -3276 -15320
rect -4076 -16080 -3276 -16040
rect -2664 -15320 -1864 -15280
rect -2664 -16040 -2624 -15320
rect -1904 -16040 -1864 -15320
rect -2664 -16080 -1864 -16040
rect -1252 -15320 -452 -15280
rect -1252 -16040 -1212 -15320
rect -492 -16040 -452 -15320
rect -1252 -16080 -452 -16040
rect 160 -15320 960 -15280
rect 160 -16040 200 -15320
rect 920 -16040 960 -15320
rect 160 -16080 960 -16040
rect 1572 -15320 2372 -15280
rect 1572 -16040 1612 -15320
rect 2332 -16040 2372 -15320
rect 1572 -16080 2372 -16040
rect 2984 -15320 3784 -15280
rect 2984 -16040 3024 -15320
rect 3744 -16040 3784 -15320
rect 2984 -16080 3784 -16040
rect 4396 -15320 5196 -15280
rect 4396 -16040 4436 -15320
rect 5156 -16040 5196 -15320
rect 4396 -16080 5196 -16040
rect 5808 -15320 6608 -15280
rect 5808 -16040 5848 -15320
rect 6568 -16040 6608 -15320
rect 5808 -16080 6608 -16040
rect 7220 -15320 8020 -15280
rect 7220 -16040 7260 -15320
rect 7980 -16040 8020 -15320
rect 7220 -16080 8020 -16040
rect 8632 -15320 9432 -15280
rect 8632 -16040 8672 -15320
rect 9392 -16040 9432 -15320
rect 8632 -16080 9432 -16040
rect 10044 -15320 10844 -15280
rect 10044 -16040 10084 -15320
rect 10804 -16040 10844 -15320
rect 10044 -16080 10844 -16040
rect 11456 -15320 12256 -15280
rect 11456 -16040 11496 -15320
rect 12216 -16040 12256 -15320
rect 11456 -16080 12256 -16040
rect 12868 -15320 13668 -15280
rect 12868 -16040 12908 -15320
rect 13628 -16040 13668 -15320
rect 12868 -16080 13668 -16040
rect 14280 -15320 15080 -15280
rect 14280 -16040 14320 -15320
rect 15040 -16040 15080 -15320
rect 14280 -16080 15080 -16040
rect 15692 -15320 16492 -15280
rect 15692 -16040 15732 -15320
rect 16452 -16040 16492 -15320
rect 15692 -16080 16492 -16040
rect 17104 -15320 17904 -15280
rect 17104 -16040 17144 -15320
rect 17864 -16040 17904 -15320
rect 17104 -16080 17904 -16040
rect 18516 -15320 19316 -15280
rect 18516 -16040 18556 -15320
rect 19276 -16040 19316 -15320
rect 18516 -16080 19316 -16040
rect 19928 -15320 20728 -15280
rect 19928 -16040 19968 -15320
rect 20688 -16040 20728 -15320
rect 19928 -16080 20728 -16040
rect 21340 -15320 22140 -15280
rect 21340 -16040 21380 -15320
rect 22100 -16040 22140 -15320
rect 21340 -16080 22140 -16040
rect 22752 -15320 23552 -15280
rect 22752 -16040 22792 -15320
rect 23512 -16040 23552 -15320
rect 22752 -16080 23552 -16040
rect -23844 -16440 -23044 -16400
rect -23844 -17160 -23804 -16440
rect -23084 -17160 -23044 -16440
rect -23844 -17200 -23044 -17160
rect -22432 -16440 -21632 -16400
rect -22432 -17160 -22392 -16440
rect -21672 -17160 -21632 -16440
rect -22432 -17200 -21632 -17160
rect -21020 -16440 -20220 -16400
rect -21020 -17160 -20980 -16440
rect -20260 -17160 -20220 -16440
rect -21020 -17200 -20220 -17160
rect -19608 -16440 -18808 -16400
rect -19608 -17160 -19568 -16440
rect -18848 -17160 -18808 -16440
rect -19608 -17200 -18808 -17160
rect -18196 -16440 -17396 -16400
rect -18196 -17160 -18156 -16440
rect -17436 -17160 -17396 -16440
rect -18196 -17200 -17396 -17160
rect -16784 -16440 -15984 -16400
rect -16784 -17160 -16744 -16440
rect -16024 -17160 -15984 -16440
rect -16784 -17200 -15984 -17160
rect -15372 -16440 -14572 -16400
rect -15372 -17160 -15332 -16440
rect -14612 -17160 -14572 -16440
rect -15372 -17200 -14572 -17160
rect -13960 -16440 -13160 -16400
rect -13960 -17160 -13920 -16440
rect -13200 -17160 -13160 -16440
rect -13960 -17200 -13160 -17160
rect -12548 -16440 -11748 -16400
rect -12548 -17160 -12508 -16440
rect -11788 -17160 -11748 -16440
rect -12548 -17200 -11748 -17160
rect -11136 -16440 -10336 -16400
rect -11136 -17160 -11096 -16440
rect -10376 -17160 -10336 -16440
rect -11136 -17200 -10336 -17160
rect -9724 -16440 -8924 -16400
rect -9724 -17160 -9684 -16440
rect -8964 -17160 -8924 -16440
rect -9724 -17200 -8924 -17160
rect -8312 -16440 -7512 -16400
rect -8312 -17160 -8272 -16440
rect -7552 -17160 -7512 -16440
rect -8312 -17200 -7512 -17160
rect -6900 -16440 -6100 -16400
rect -6900 -17160 -6860 -16440
rect -6140 -17160 -6100 -16440
rect -6900 -17200 -6100 -17160
rect -5488 -16440 -4688 -16400
rect -5488 -17160 -5448 -16440
rect -4728 -17160 -4688 -16440
rect -5488 -17200 -4688 -17160
rect -4076 -16440 -3276 -16400
rect -4076 -17160 -4036 -16440
rect -3316 -17160 -3276 -16440
rect -4076 -17200 -3276 -17160
rect -2664 -16440 -1864 -16400
rect -2664 -17160 -2624 -16440
rect -1904 -17160 -1864 -16440
rect -2664 -17200 -1864 -17160
rect -1252 -16440 -452 -16400
rect -1252 -17160 -1212 -16440
rect -492 -17160 -452 -16440
rect -1252 -17200 -452 -17160
rect 160 -16440 960 -16400
rect 160 -17160 200 -16440
rect 920 -17160 960 -16440
rect 160 -17200 960 -17160
rect 1572 -16440 2372 -16400
rect 1572 -17160 1612 -16440
rect 2332 -17160 2372 -16440
rect 1572 -17200 2372 -17160
rect 2984 -16440 3784 -16400
rect 2984 -17160 3024 -16440
rect 3744 -17160 3784 -16440
rect 2984 -17200 3784 -17160
rect 4396 -16440 5196 -16400
rect 4396 -17160 4436 -16440
rect 5156 -17160 5196 -16440
rect 4396 -17200 5196 -17160
rect 5808 -16440 6608 -16400
rect 5808 -17160 5848 -16440
rect 6568 -17160 6608 -16440
rect 5808 -17200 6608 -17160
rect 7220 -16440 8020 -16400
rect 7220 -17160 7260 -16440
rect 7980 -17160 8020 -16440
rect 7220 -17200 8020 -17160
rect 8632 -16440 9432 -16400
rect 8632 -17160 8672 -16440
rect 9392 -17160 9432 -16440
rect 8632 -17200 9432 -17160
rect 10044 -16440 10844 -16400
rect 10044 -17160 10084 -16440
rect 10804 -17160 10844 -16440
rect 10044 -17200 10844 -17160
rect 11456 -16440 12256 -16400
rect 11456 -17160 11496 -16440
rect 12216 -17160 12256 -16440
rect 11456 -17200 12256 -17160
rect 12868 -16440 13668 -16400
rect 12868 -17160 12908 -16440
rect 13628 -17160 13668 -16440
rect 12868 -17200 13668 -17160
rect 14280 -16440 15080 -16400
rect 14280 -17160 14320 -16440
rect 15040 -17160 15080 -16440
rect 14280 -17200 15080 -17160
rect 15692 -16440 16492 -16400
rect 15692 -17160 15732 -16440
rect 16452 -17160 16492 -16440
rect 15692 -17200 16492 -17160
rect 17104 -16440 17904 -16400
rect 17104 -17160 17144 -16440
rect 17864 -17160 17904 -16440
rect 17104 -17200 17904 -17160
rect 18516 -16440 19316 -16400
rect 18516 -17160 18556 -16440
rect 19276 -17160 19316 -16440
rect 18516 -17200 19316 -17160
rect 19928 -16440 20728 -16400
rect 19928 -17160 19968 -16440
rect 20688 -17160 20728 -16440
rect 19928 -17200 20728 -17160
rect 21340 -16440 22140 -16400
rect 21340 -17160 21380 -16440
rect 22100 -17160 22140 -16440
rect 21340 -17200 22140 -17160
rect 22752 -16440 23552 -16400
rect 22752 -17160 22792 -16440
rect 23512 -17160 23552 -16440
rect 22752 -17200 23552 -17160
rect -23844 -17560 -23044 -17520
rect -23844 -18280 -23804 -17560
rect -23084 -18280 -23044 -17560
rect -23844 -18320 -23044 -18280
rect -22432 -17560 -21632 -17520
rect -22432 -18280 -22392 -17560
rect -21672 -18280 -21632 -17560
rect -22432 -18320 -21632 -18280
rect -21020 -17560 -20220 -17520
rect -21020 -18280 -20980 -17560
rect -20260 -18280 -20220 -17560
rect -21020 -18320 -20220 -18280
rect -19608 -17560 -18808 -17520
rect -19608 -18280 -19568 -17560
rect -18848 -18280 -18808 -17560
rect -19608 -18320 -18808 -18280
rect -18196 -17560 -17396 -17520
rect -18196 -18280 -18156 -17560
rect -17436 -18280 -17396 -17560
rect -18196 -18320 -17396 -18280
rect -16784 -17560 -15984 -17520
rect -16784 -18280 -16744 -17560
rect -16024 -18280 -15984 -17560
rect -16784 -18320 -15984 -18280
rect -15372 -17560 -14572 -17520
rect -15372 -18280 -15332 -17560
rect -14612 -18280 -14572 -17560
rect -15372 -18320 -14572 -18280
rect -13960 -17560 -13160 -17520
rect -13960 -18280 -13920 -17560
rect -13200 -18280 -13160 -17560
rect -13960 -18320 -13160 -18280
rect -12548 -17560 -11748 -17520
rect -12548 -18280 -12508 -17560
rect -11788 -18280 -11748 -17560
rect -12548 -18320 -11748 -18280
rect -11136 -17560 -10336 -17520
rect -11136 -18280 -11096 -17560
rect -10376 -18280 -10336 -17560
rect -11136 -18320 -10336 -18280
rect -9724 -17560 -8924 -17520
rect -9724 -18280 -9684 -17560
rect -8964 -18280 -8924 -17560
rect -9724 -18320 -8924 -18280
rect -8312 -17560 -7512 -17520
rect -8312 -18280 -8272 -17560
rect -7552 -18280 -7512 -17560
rect -8312 -18320 -7512 -18280
rect -6900 -17560 -6100 -17520
rect -6900 -18280 -6860 -17560
rect -6140 -18280 -6100 -17560
rect -6900 -18320 -6100 -18280
rect -5488 -17560 -4688 -17520
rect -5488 -18280 -5448 -17560
rect -4728 -18280 -4688 -17560
rect -5488 -18320 -4688 -18280
rect -4076 -17560 -3276 -17520
rect -4076 -18280 -4036 -17560
rect -3316 -18280 -3276 -17560
rect -4076 -18320 -3276 -18280
rect -2664 -17560 -1864 -17520
rect -2664 -18280 -2624 -17560
rect -1904 -18280 -1864 -17560
rect -2664 -18320 -1864 -18280
rect -1252 -17560 -452 -17520
rect -1252 -18280 -1212 -17560
rect -492 -18280 -452 -17560
rect -1252 -18320 -452 -18280
rect 160 -17560 960 -17520
rect 160 -18280 200 -17560
rect 920 -18280 960 -17560
rect 160 -18320 960 -18280
rect 1572 -17560 2372 -17520
rect 1572 -18280 1612 -17560
rect 2332 -18280 2372 -17560
rect 1572 -18320 2372 -18280
rect 2984 -17560 3784 -17520
rect 2984 -18280 3024 -17560
rect 3744 -18280 3784 -17560
rect 2984 -18320 3784 -18280
rect 4396 -17560 5196 -17520
rect 4396 -18280 4436 -17560
rect 5156 -18280 5196 -17560
rect 4396 -18320 5196 -18280
rect 5808 -17560 6608 -17520
rect 5808 -18280 5848 -17560
rect 6568 -18280 6608 -17560
rect 5808 -18320 6608 -18280
rect 7220 -17560 8020 -17520
rect 7220 -18280 7260 -17560
rect 7980 -18280 8020 -17560
rect 7220 -18320 8020 -18280
rect 8632 -17560 9432 -17520
rect 8632 -18280 8672 -17560
rect 9392 -18280 9432 -17560
rect 8632 -18320 9432 -18280
rect 10044 -17560 10844 -17520
rect 10044 -18280 10084 -17560
rect 10804 -18280 10844 -17560
rect 10044 -18320 10844 -18280
rect 11456 -17560 12256 -17520
rect 11456 -18280 11496 -17560
rect 12216 -18280 12256 -17560
rect 11456 -18320 12256 -18280
rect 12868 -17560 13668 -17520
rect 12868 -18280 12908 -17560
rect 13628 -18280 13668 -17560
rect 12868 -18320 13668 -18280
rect 14280 -17560 15080 -17520
rect 14280 -18280 14320 -17560
rect 15040 -18280 15080 -17560
rect 14280 -18320 15080 -18280
rect 15692 -17560 16492 -17520
rect 15692 -18280 15732 -17560
rect 16452 -18280 16492 -17560
rect 15692 -18320 16492 -18280
rect 17104 -17560 17904 -17520
rect 17104 -18280 17144 -17560
rect 17864 -18280 17904 -17560
rect 17104 -18320 17904 -18280
rect 18516 -17560 19316 -17520
rect 18516 -18280 18556 -17560
rect 19276 -18280 19316 -17560
rect 18516 -18320 19316 -18280
rect 19928 -17560 20728 -17520
rect 19928 -18280 19968 -17560
rect 20688 -18280 20728 -17560
rect 19928 -18320 20728 -18280
rect 21340 -17560 22140 -17520
rect 21340 -18280 21380 -17560
rect 22100 -18280 22140 -17560
rect 21340 -18320 22140 -18280
rect 22752 -17560 23552 -17520
rect 22752 -18280 22792 -17560
rect 23512 -18280 23552 -17560
rect 22752 -18320 23552 -18280
<< mimcapcontact >>
rect -23804 17560 -23084 18280
rect -22392 17560 -21672 18280
rect -20980 17560 -20260 18280
rect -19568 17560 -18848 18280
rect -18156 17560 -17436 18280
rect -16744 17560 -16024 18280
rect -15332 17560 -14612 18280
rect -13920 17560 -13200 18280
rect -12508 17560 -11788 18280
rect -11096 17560 -10376 18280
rect -9684 17560 -8964 18280
rect -8272 17560 -7552 18280
rect -6860 17560 -6140 18280
rect -5448 17560 -4728 18280
rect -4036 17560 -3316 18280
rect -2624 17560 -1904 18280
rect -1212 17560 -492 18280
rect 200 17560 920 18280
rect 1612 17560 2332 18280
rect 3024 17560 3744 18280
rect 4436 17560 5156 18280
rect 5848 17560 6568 18280
rect 7260 17560 7980 18280
rect 8672 17560 9392 18280
rect 10084 17560 10804 18280
rect 11496 17560 12216 18280
rect 12908 17560 13628 18280
rect 14320 17560 15040 18280
rect 15732 17560 16452 18280
rect 17144 17560 17864 18280
rect 18556 17560 19276 18280
rect 19968 17560 20688 18280
rect 21380 17560 22100 18280
rect 22792 17560 23512 18280
rect -23804 16440 -23084 17160
rect -22392 16440 -21672 17160
rect -20980 16440 -20260 17160
rect -19568 16440 -18848 17160
rect -18156 16440 -17436 17160
rect -16744 16440 -16024 17160
rect -15332 16440 -14612 17160
rect -13920 16440 -13200 17160
rect -12508 16440 -11788 17160
rect -11096 16440 -10376 17160
rect -9684 16440 -8964 17160
rect -8272 16440 -7552 17160
rect -6860 16440 -6140 17160
rect -5448 16440 -4728 17160
rect -4036 16440 -3316 17160
rect -2624 16440 -1904 17160
rect -1212 16440 -492 17160
rect 200 16440 920 17160
rect 1612 16440 2332 17160
rect 3024 16440 3744 17160
rect 4436 16440 5156 17160
rect 5848 16440 6568 17160
rect 7260 16440 7980 17160
rect 8672 16440 9392 17160
rect 10084 16440 10804 17160
rect 11496 16440 12216 17160
rect 12908 16440 13628 17160
rect 14320 16440 15040 17160
rect 15732 16440 16452 17160
rect 17144 16440 17864 17160
rect 18556 16440 19276 17160
rect 19968 16440 20688 17160
rect 21380 16440 22100 17160
rect 22792 16440 23512 17160
rect -23804 15320 -23084 16040
rect -22392 15320 -21672 16040
rect -20980 15320 -20260 16040
rect -19568 15320 -18848 16040
rect -18156 15320 -17436 16040
rect -16744 15320 -16024 16040
rect -15332 15320 -14612 16040
rect -13920 15320 -13200 16040
rect -12508 15320 -11788 16040
rect -11096 15320 -10376 16040
rect -9684 15320 -8964 16040
rect -8272 15320 -7552 16040
rect -6860 15320 -6140 16040
rect -5448 15320 -4728 16040
rect -4036 15320 -3316 16040
rect -2624 15320 -1904 16040
rect -1212 15320 -492 16040
rect 200 15320 920 16040
rect 1612 15320 2332 16040
rect 3024 15320 3744 16040
rect 4436 15320 5156 16040
rect 5848 15320 6568 16040
rect 7260 15320 7980 16040
rect 8672 15320 9392 16040
rect 10084 15320 10804 16040
rect 11496 15320 12216 16040
rect 12908 15320 13628 16040
rect 14320 15320 15040 16040
rect 15732 15320 16452 16040
rect 17144 15320 17864 16040
rect 18556 15320 19276 16040
rect 19968 15320 20688 16040
rect 21380 15320 22100 16040
rect 22792 15320 23512 16040
rect -23804 14200 -23084 14920
rect -22392 14200 -21672 14920
rect -20980 14200 -20260 14920
rect -19568 14200 -18848 14920
rect -18156 14200 -17436 14920
rect -16744 14200 -16024 14920
rect -15332 14200 -14612 14920
rect -13920 14200 -13200 14920
rect -12508 14200 -11788 14920
rect -11096 14200 -10376 14920
rect -9684 14200 -8964 14920
rect -8272 14200 -7552 14920
rect -6860 14200 -6140 14920
rect -5448 14200 -4728 14920
rect -4036 14200 -3316 14920
rect -2624 14200 -1904 14920
rect -1212 14200 -492 14920
rect 200 14200 920 14920
rect 1612 14200 2332 14920
rect 3024 14200 3744 14920
rect 4436 14200 5156 14920
rect 5848 14200 6568 14920
rect 7260 14200 7980 14920
rect 8672 14200 9392 14920
rect 10084 14200 10804 14920
rect 11496 14200 12216 14920
rect 12908 14200 13628 14920
rect 14320 14200 15040 14920
rect 15732 14200 16452 14920
rect 17144 14200 17864 14920
rect 18556 14200 19276 14920
rect 19968 14200 20688 14920
rect 21380 14200 22100 14920
rect 22792 14200 23512 14920
rect -23804 13080 -23084 13800
rect -22392 13080 -21672 13800
rect -20980 13080 -20260 13800
rect -19568 13080 -18848 13800
rect -18156 13080 -17436 13800
rect -16744 13080 -16024 13800
rect -15332 13080 -14612 13800
rect -13920 13080 -13200 13800
rect -12508 13080 -11788 13800
rect -11096 13080 -10376 13800
rect -9684 13080 -8964 13800
rect -8272 13080 -7552 13800
rect -6860 13080 -6140 13800
rect -5448 13080 -4728 13800
rect -4036 13080 -3316 13800
rect -2624 13080 -1904 13800
rect -1212 13080 -492 13800
rect 200 13080 920 13800
rect 1612 13080 2332 13800
rect 3024 13080 3744 13800
rect 4436 13080 5156 13800
rect 5848 13080 6568 13800
rect 7260 13080 7980 13800
rect 8672 13080 9392 13800
rect 10084 13080 10804 13800
rect 11496 13080 12216 13800
rect 12908 13080 13628 13800
rect 14320 13080 15040 13800
rect 15732 13080 16452 13800
rect 17144 13080 17864 13800
rect 18556 13080 19276 13800
rect 19968 13080 20688 13800
rect 21380 13080 22100 13800
rect 22792 13080 23512 13800
rect -23804 11960 -23084 12680
rect -22392 11960 -21672 12680
rect -20980 11960 -20260 12680
rect -19568 11960 -18848 12680
rect -18156 11960 -17436 12680
rect -16744 11960 -16024 12680
rect -15332 11960 -14612 12680
rect -13920 11960 -13200 12680
rect -12508 11960 -11788 12680
rect -11096 11960 -10376 12680
rect -9684 11960 -8964 12680
rect -8272 11960 -7552 12680
rect -6860 11960 -6140 12680
rect -5448 11960 -4728 12680
rect -4036 11960 -3316 12680
rect -2624 11960 -1904 12680
rect -1212 11960 -492 12680
rect 200 11960 920 12680
rect 1612 11960 2332 12680
rect 3024 11960 3744 12680
rect 4436 11960 5156 12680
rect 5848 11960 6568 12680
rect 7260 11960 7980 12680
rect 8672 11960 9392 12680
rect 10084 11960 10804 12680
rect 11496 11960 12216 12680
rect 12908 11960 13628 12680
rect 14320 11960 15040 12680
rect 15732 11960 16452 12680
rect 17144 11960 17864 12680
rect 18556 11960 19276 12680
rect 19968 11960 20688 12680
rect 21380 11960 22100 12680
rect 22792 11960 23512 12680
rect -23804 10840 -23084 11560
rect -22392 10840 -21672 11560
rect -20980 10840 -20260 11560
rect -19568 10840 -18848 11560
rect -18156 10840 -17436 11560
rect -16744 10840 -16024 11560
rect -15332 10840 -14612 11560
rect -13920 10840 -13200 11560
rect -12508 10840 -11788 11560
rect -11096 10840 -10376 11560
rect -9684 10840 -8964 11560
rect -8272 10840 -7552 11560
rect -6860 10840 -6140 11560
rect -5448 10840 -4728 11560
rect -4036 10840 -3316 11560
rect -2624 10840 -1904 11560
rect -1212 10840 -492 11560
rect 200 10840 920 11560
rect 1612 10840 2332 11560
rect 3024 10840 3744 11560
rect 4436 10840 5156 11560
rect 5848 10840 6568 11560
rect 7260 10840 7980 11560
rect 8672 10840 9392 11560
rect 10084 10840 10804 11560
rect 11496 10840 12216 11560
rect 12908 10840 13628 11560
rect 14320 10840 15040 11560
rect 15732 10840 16452 11560
rect 17144 10840 17864 11560
rect 18556 10840 19276 11560
rect 19968 10840 20688 11560
rect 21380 10840 22100 11560
rect 22792 10840 23512 11560
rect -23804 9720 -23084 10440
rect -22392 9720 -21672 10440
rect -20980 9720 -20260 10440
rect -19568 9720 -18848 10440
rect -18156 9720 -17436 10440
rect -16744 9720 -16024 10440
rect -15332 9720 -14612 10440
rect -13920 9720 -13200 10440
rect -12508 9720 -11788 10440
rect -11096 9720 -10376 10440
rect -9684 9720 -8964 10440
rect -8272 9720 -7552 10440
rect -6860 9720 -6140 10440
rect -5448 9720 -4728 10440
rect -4036 9720 -3316 10440
rect -2624 9720 -1904 10440
rect -1212 9720 -492 10440
rect 200 9720 920 10440
rect 1612 9720 2332 10440
rect 3024 9720 3744 10440
rect 4436 9720 5156 10440
rect 5848 9720 6568 10440
rect 7260 9720 7980 10440
rect 8672 9720 9392 10440
rect 10084 9720 10804 10440
rect 11496 9720 12216 10440
rect 12908 9720 13628 10440
rect 14320 9720 15040 10440
rect 15732 9720 16452 10440
rect 17144 9720 17864 10440
rect 18556 9720 19276 10440
rect 19968 9720 20688 10440
rect 21380 9720 22100 10440
rect 22792 9720 23512 10440
rect -23804 8600 -23084 9320
rect -22392 8600 -21672 9320
rect -20980 8600 -20260 9320
rect -19568 8600 -18848 9320
rect -18156 8600 -17436 9320
rect -16744 8600 -16024 9320
rect -15332 8600 -14612 9320
rect -13920 8600 -13200 9320
rect -12508 8600 -11788 9320
rect -11096 8600 -10376 9320
rect -9684 8600 -8964 9320
rect -8272 8600 -7552 9320
rect -6860 8600 -6140 9320
rect -5448 8600 -4728 9320
rect -4036 8600 -3316 9320
rect -2624 8600 -1904 9320
rect -1212 8600 -492 9320
rect 200 8600 920 9320
rect 1612 8600 2332 9320
rect 3024 8600 3744 9320
rect 4436 8600 5156 9320
rect 5848 8600 6568 9320
rect 7260 8600 7980 9320
rect 8672 8600 9392 9320
rect 10084 8600 10804 9320
rect 11496 8600 12216 9320
rect 12908 8600 13628 9320
rect 14320 8600 15040 9320
rect 15732 8600 16452 9320
rect 17144 8600 17864 9320
rect 18556 8600 19276 9320
rect 19968 8600 20688 9320
rect 21380 8600 22100 9320
rect 22792 8600 23512 9320
rect -23804 7480 -23084 8200
rect -22392 7480 -21672 8200
rect -20980 7480 -20260 8200
rect -19568 7480 -18848 8200
rect -18156 7480 -17436 8200
rect -16744 7480 -16024 8200
rect -15332 7480 -14612 8200
rect -13920 7480 -13200 8200
rect -12508 7480 -11788 8200
rect -11096 7480 -10376 8200
rect -9684 7480 -8964 8200
rect -8272 7480 -7552 8200
rect -6860 7480 -6140 8200
rect -5448 7480 -4728 8200
rect -4036 7480 -3316 8200
rect -2624 7480 -1904 8200
rect -1212 7480 -492 8200
rect 200 7480 920 8200
rect 1612 7480 2332 8200
rect 3024 7480 3744 8200
rect 4436 7480 5156 8200
rect 5848 7480 6568 8200
rect 7260 7480 7980 8200
rect 8672 7480 9392 8200
rect 10084 7480 10804 8200
rect 11496 7480 12216 8200
rect 12908 7480 13628 8200
rect 14320 7480 15040 8200
rect 15732 7480 16452 8200
rect 17144 7480 17864 8200
rect 18556 7480 19276 8200
rect 19968 7480 20688 8200
rect 21380 7480 22100 8200
rect 22792 7480 23512 8200
rect -23804 6360 -23084 7080
rect -22392 6360 -21672 7080
rect -20980 6360 -20260 7080
rect -19568 6360 -18848 7080
rect -18156 6360 -17436 7080
rect -16744 6360 -16024 7080
rect -15332 6360 -14612 7080
rect -13920 6360 -13200 7080
rect -12508 6360 -11788 7080
rect -11096 6360 -10376 7080
rect -9684 6360 -8964 7080
rect -8272 6360 -7552 7080
rect -6860 6360 -6140 7080
rect -5448 6360 -4728 7080
rect -4036 6360 -3316 7080
rect -2624 6360 -1904 7080
rect -1212 6360 -492 7080
rect 200 6360 920 7080
rect 1612 6360 2332 7080
rect 3024 6360 3744 7080
rect 4436 6360 5156 7080
rect 5848 6360 6568 7080
rect 7260 6360 7980 7080
rect 8672 6360 9392 7080
rect 10084 6360 10804 7080
rect 11496 6360 12216 7080
rect 12908 6360 13628 7080
rect 14320 6360 15040 7080
rect 15732 6360 16452 7080
rect 17144 6360 17864 7080
rect 18556 6360 19276 7080
rect 19968 6360 20688 7080
rect 21380 6360 22100 7080
rect 22792 6360 23512 7080
rect -23804 5240 -23084 5960
rect -22392 5240 -21672 5960
rect -20980 5240 -20260 5960
rect -19568 5240 -18848 5960
rect -18156 5240 -17436 5960
rect -16744 5240 -16024 5960
rect -15332 5240 -14612 5960
rect -13920 5240 -13200 5960
rect -12508 5240 -11788 5960
rect -11096 5240 -10376 5960
rect -9684 5240 -8964 5960
rect -8272 5240 -7552 5960
rect -6860 5240 -6140 5960
rect -5448 5240 -4728 5960
rect -4036 5240 -3316 5960
rect -2624 5240 -1904 5960
rect -1212 5240 -492 5960
rect 200 5240 920 5960
rect 1612 5240 2332 5960
rect 3024 5240 3744 5960
rect 4436 5240 5156 5960
rect 5848 5240 6568 5960
rect 7260 5240 7980 5960
rect 8672 5240 9392 5960
rect 10084 5240 10804 5960
rect 11496 5240 12216 5960
rect 12908 5240 13628 5960
rect 14320 5240 15040 5960
rect 15732 5240 16452 5960
rect 17144 5240 17864 5960
rect 18556 5240 19276 5960
rect 19968 5240 20688 5960
rect 21380 5240 22100 5960
rect 22792 5240 23512 5960
rect -23804 4120 -23084 4840
rect -22392 4120 -21672 4840
rect -20980 4120 -20260 4840
rect -19568 4120 -18848 4840
rect -18156 4120 -17436 4840
rect -16744 4120 -16024 4840
rect -15332 4120 -14612 4840
rect -13920 4120 -13200 4840
rect -12508 4120 -11788 4840
rect -11096 4120 -10376 4840
rect -9684 4120 -8964 4840
rect -8272 4120 -7552 4840
rect -6860 4120 -6140 4840
rect -5448 4120 -4728 4840
rect -4036 4120 -3316 4840
rect -2624 4120 -1904 4840
rect -1212 4120 -492 4840
rect 200 4120 920 4840
rect 1612 4120 2332 4840
rect 3024 4120 3744 4840
rect 4436 4120 5156 4840
rect 5848 4120 6568 4840
rect 7260 4120 7980 4840
rect 8672 4120 9392 4840
rect 10084 4120 10804 4840
rect 11496 4120 12216 4840
rect 12908 4120 13628 4840
rect 14320 4120 15040 4840
rect 15732 4120 16452 4840
rect 17144 4120 17864 4840
rect 18556 4120 19276 4840
rect 19968 4120 20688 4840
rect 21380 4120 22100 4840
rect 22792 4120 23512 4840
rect -23804 3000 -23084 3720
rect -22392 3000 -21672 3720
rect -20980 3000 -20260 3720
rect -19568 3000 -18848 3720
rect -18156 3000 -17436 3720
rect -16744 3000 -16024 3720
rect -15332 3000 -14612 3720
rect -13920 3000 -13200 3720
rect -12508 3000 -11788 3720
rect -11096 3000 -10376 3720
rect -9684 3000 -8964 3720
rect -8272 3000 -7552 3720
rect -6860 3000 -6140 3720
rect -5448 3000 -4728 3720
rect -4036 3000 -3316 3720
rect -2624 3000 -1904 3720
rect -1212 3000 -492 3720
rect 200 3000 920 3720
rect 1612 3000 2332 3720
rect 3024 3000 3744 3720
rect 4436 3000 5156 3720
rect 5848 3000 6568 3720
rect 7260 3000 7980 3720
rect 8672 3000 9392 3720
rect 10084 3000 10804 3720
rect 11496 3000 12216 3720
rect 12908 3000 13628 3720
rect 14320 3000 15040 3720
rect 15732 3000 16452 3720
rect 17144 3000 17864 3720
rect 18556 3000 19276 3720
rect 19968 3000 20688 3720
rect 21380 3000 22100 3720
rect 22792 3000 23512 3720
rect -23804 1880 -23084 2600
rect -22392 1880 -21672 2600
rect -20980 1880 -20260 2600
rect -19568 1880 -18848 2600
rect -18156 1880 -17436 2600
rect -16744 1880 -16024 2600
rect -15332 1880 -14612 2600
rect -13920 1880 -13200 2600
rect -12508 1880 -11788 2600
rect -11096 1880 -10376 2600
rect -9684 1880 -8964 2600
rect -8272 1880 -7552 2600
rect -6860 1880 -6140 2600
rect -5448 1880 -4728 2600
rect -4036 1880 -3316 2600
rect -2624 1880 -1904 2600
rect -1212 1880 -492 2600
rect 200 1880 920 2600
rect 1612 1880 2332 2600
rect 3024 1880 3744 2600
rect 4436 1880 5156 2600
rect 5848 1880 6568 2600
rect 7260 1880 7980 2600
rect 8672 1880 9392 2600
rect 10084 1880 10804 2600
rect 11496 1880 12216 2600
rect 12908 1880 13628 2600
rect 14320 1880 15040 2600
rect 15732 1880 16452 2600
rect 17144 1880 17864 2600
rect 18556 1880 19276 2600
rect 19968 1880 20688 2600
rect 21380 1880 22100 2600
rect 22792 1880 23512 2600
rect -23804 760 -23084 1480
rect -22392 760 -21672 1480
rect -20980 760 -20260 1480
rect -19568 760 -18848 1480
rect -18156 760 -17436 1480
rect -16744 760 -16024 1480
rect -15332 760 -14612 1480
rect -13920 760 -13200 1480
rect -12508 760 -11788 1480
rect -11096 760 -10376 1480
rect -9684 760 -8964 1480
rect -8272 760 -7552 1480
rect -6860 760 -6140 1480
rect -5448 760 -4728 1480
rect -4036 760 -3316 1480
rect -2624 760 -1904 1480
rect -1212 760 -492 1480
rect 200 760 920 1480
rect 1612 760 2332 1480
rect 3024 760 3744 1480
rect 4436 760 5156 1480
rect 5848 760 6568 1480
rect 7260 760 7980 1480
rect 8672 760 9392 1480
rect 10084 760 10804 1480
rect 11496 760 12216 1480
rect 12908 760 13628 1480
rect 14320 760 15040 1480
rect 15732 760 16452 1480
rect 17144 760 17864 1480
rect 18556 760 19276 1480
rect 19968 760 20688 1480
rect 21380 760 22100 1480
rect 22792 760 23512 1480
rect -23804 -360 -23084 360
rect -22392 -360 -21672 360
rect -20980 -360 -20260 360
rect -19568 -360 -18848 360
rect -18156 -360 -17436 360
rect -16744 -360 -16024 360
rect -15332 -360 -14612 360
rect -13920 -360 -13200 360
rect -12508 -360 -11788 360
rect -11096 -360 -10376 360
rect -9684 -360 -8964 360
rect -8272 -360 -7552 360
rect -6860 -360 -6140 360
rect -5448 -360 -4728 360
rect -4036 -360 -3316 360
rect -2624 -360 -1904 360
rect -1212 -360 -492 360
rect 200 -360 920 360
rect 1612 -360 2332 360
rect 3024 -360 3744 360
rect 4436 -360 5156 360
rect 5848 -360 6568 360
rect 7260 -360 7980 360
rect 8672 -360 9392 360
rect 10084 -360 10804 360
rect 11496 -360 12216 360
rect 12908 -360 13628 360
rect 14320 -360 15040 360
rect 15732 -360 16452 360
rect 17144 -360 17864 360
rect 18556 -360 19276 360
rect 19968 -360 20688 360
rect 21380 -360 22100 360
rect 22792 -360 23512 360
rect -23804 -1480 -23084 -760
rect -22392 -1480 -21672 -760
rect -20980 -1480 -20260 -760
rect -19568 -1480 -18848 -760
rect -18156 -1480 -17436 -760
rect -16744 -1480 -16024 -760
rect -15332 -1480 -14612 -760
rect -13920 -1480 -13200 -760
rect -12508 -1480 -11788 -760
rect -11096 -1480 -10376 -760
rect -9684 -1480 -8964 -760
rect -8272 -1480 -7552 -760
rect -6860 -1480 -6140 -760
rect -5448 -1480 -4728 -760
rect -4036 -1480 -3316 -760
rect -2624 -1480 -1904 -760
rect -1212 -1480 -492 -760
rect 200 -1480 920 -760
rect 1612 -1480 2332 -760
rect 3024 -1480 3744 -760
rect 4436 -1480 5156 -760
rect 5848 -1480 6568 -760
rect 7260 -1480 7980 -760
rect 8672 -1480 9392 -760
rect 10084 -1480 10804 -760
rect 11496 -1480 12216 -760
rect 12908 -1480 13628 -760
rect 14320 -1480 15040 -760
rect 15732 -1480 16452 -760
rect 17144 -1480 17864 -760
rect 18556 -1480 19276 -760
rect 19968 -1480 20688 -760
rect 21380 -1480 22100 -760
rect 22792 -1480 23512 -760
rect -23804 -2600 -23084 -1880
rect -22392 -2600 -21672 -1880
rect -20980 -2600 -20260 -1880
rect -19568 -2600 -18848 -1880
rect -18156 -2600 -17436 -1880
rect -16744 -2600 -16024 -1880
rect -15332 -2600 -14612 -1880
rect -13920 -2600 -13200 -1880
rect -12508 -2600 -11788 -1880
rect -11096 -2600 -10376 -1880
rect -9684 -2600 -8964 -1880
rect -8272 -2600 -7552 -1880
rect -6860 -2600 -6140 -1880
rect -5448 -2600 -4728 -1880
rect -4036 -2600 -3316 -1880
rect -2624 -2600 -1904 -1880
rect -1212 -2600 -492 -1880
rect 200 -2600 920 -1880
rect 1612 -2600 2332 -1880
rect 3024 -2600 3744 -1880
rect 4436 -2600 5156 -1880
rect 5848 -2600 6568 -1880
rect 7260 -2600 7980 -1880
rect 8672 -2600 9392 -1880
rect 10084 -2600 10804 -1880
rect 11496 -2600 12216 -1880
rect 12908 -2600 13628 -1880
rect 14320 -2600 15040 -1880
rect 15732 -2600 16452 -1880
rect 17144 -2600 17864 -1880
rect 18556 -2600 19276 -1880
rect 19968 -2600 20688 -1880
rect 21380 -2600 22100 -1880
rect 22792 -2600 23512 -1880
rect -23804 -3720 -23084 -3000
rect -22392 -3720 -21672 -3000
rect -20980 -3720 -20260 -3000
rect -19568 -3720 -18848 -3000
rect -18156 -3720 -17436 -3000
rect -16744 -3720 -16024 -3000
rect -15332 -3720 -14612 -3000
rect -13920 -3720 -13200 -3000
rect -12508 -3720 -11788 -3000
rect -11096 -3720 -10376 -3000
rect -9684 -3720 -8964 -3000
rect -8272 -3720 -7552 -3000
rect -6860 -3720 -6140 -3000
rect -5448 -3720 -4728 -3000
rect -4036 -3720 -3316 -3000
rect -2624 -3720 -1904 -3000
rect -1212 -3720 -492 -3000
rect 200 -3720 920 -3000
rect 1612 -3720 2332 -3000
rect 3024 -3720 3744 -3000
rect 4436 -3720 5156 -3000
rect 5848 -3720 6568 -3000
rect 7260 -3720 7980 -3000
rect 8672 -3720 9392 -3000
rect 10084 -3720 10804 -3000
rect 11496 -3720 12216 -3000
rect 12908 -3720 13628 -3000
rect 14320 -3720 15040 -3000
rect 15732 -3720 16452 -3000
rect 17144 -3720 17864 -3000
rect 18556 -3720 19276 -3000
rect 19968 -3720 20688 -3000
rect 21380 -3720 22100 -3000
rect 22792 -3720 23512 -3000
rect -23804 -4840 -23084 -4120
rect -22392 -4840 -21672 -4120
rect -20980 -4840 -20260 -4120
rect -19568 -4840 -18848 -4120
rect -18156 -4840 -17436 -4120
rect -16744 -4840 -16024 -4120
rect -15332 -4840 -14612 -4120
rect -13920 -4840 -13200 -4120
rect -12508 -4840 -11788 -4120
rect -11096 -4840 -10376 -4120
rect -9684 -4840 -8964 -4120
rect -8272 -4840 -7552 -4120
rect -6860 -4840 -6140 -4120
rect -5448 -4840 -4728 -4120
rect -4036 -4840 -3316 -4120
rect -2624 -4840 -1904 -4120
rect -1212 -4840 -492 -4120
rect 200 -4840 920 -4120
rect 1612 -4840 2332 -4120
rect 3024 -4840 3744 -4120
rect 4436 -4840 5156 -4120
rect 5848 -4840 6568 -4120
rect 7260 -4840 7980 -4120
rect 8672 -4840 9392 -4120
rect 10084 -4840 10804 -4120
rect 11496 -4840 12216 -4120
rect 12908 -4840 13628 -4120
rect 14320 -4840 15040 -4120
rect 15732 -4840 16452 -4120
rect 17144 -4840 17864 -4120
rect 18556 -4840 19276 -4120
rect 19968 -4840 20688 -4120
rect 21380 -4840 22100 -4120
rect 22792 -4840 23512 -4120
rect -23804 -5960 -23084 -5240
rect -22392 -5960 -21672 -5240
rect -20980 -5960 -20260 -5240
rect -19568 -5960 -18848 -5240
rect -18156 -5960 -17436 -5240
rect -16744 -5960 -16024 -5240
rect -15332 -5960 -14612 -5240
rect -13920 -5960 -13200 -5240
rect -12508 -5960 -11788 -5240
rect -11096 -5960 -10376 -5240
rect -9684 -5960 -8964 -5240
rect -8272 -5960 -7552 -5240
rect -6860 -5960 -6140 -5240
rect -5448 -5960 -4728 -5240
rect -4036 -5960 -3316 -5240
rect -2624 -5960 -1904 -5240
rect -1212 -5960 -492 -5240
rect 200 -5960 920 -5240
rect 1612 -5960 2332 -5240
rect 3024 -5960 3744 -5240
rect 4436 -5960 5156 -5240
rect 5848 -5960 6568 -5240
rect 7260 -5960 7980 -5240
rect 8672 -5960 9392 -5240
rect 10084 -5960 10804 -5240
rect 11496 -5960 12216 -5240
rect 12908 -5960 13628 -5240
rect 14320 -5960 15040 -5240
rect 15732 -5960 16452 -5240
rect 17144 -5960 17864 -5240
rect 18556 -5960 19276 -5240
rect 19968 -5960 20688 -5240
rect 21380 -5960 22100 -5240
rect 22792 -5960 23512 -5240
rect -23804 -7080 -23084 -6360
rect -22392 -7080 -21672 -6360
rect -20980 -7080 -20260 -6360
rect -19568 -7080 -18848 -6360
rect -18156 -7080 -17436 -6360
rect -16744 -7080 -16024 -6360
rect -15332 -7080 -14612 -6360
rect -13920 -7080 -13200 -6360
rect -12508 -7080 -11788 -6360
rect -11096 -7080 -10376 -6360
rect -9684 -7080 -8964 -6360
rect -8272 -7080 -7552 -6360
rect -6860 -7080 -6140 -6360
rect -5448 -7080 -4728 -6360
rect -4036 -7080 -3316 -6360
rect -2624 -7080 -1904 -6360
rect -1212 -7080 -492 -6360
rect 200 -7080 920 -6360
rect 1612 -7080 2332 -6360
rect 3024 -7080 3744 -6360
rect 4436 -7080 5156 -6360
rect 5848 -7080 6568 -6360
rect 7260 -7080 7980 -6360
rect 8672 -7080 9392 -6360
rect 10084 -7080 10804 -6360
rect 11496 -7080 12216 -6360
rect 12908 -7080 13628 -6360
rect 14320 -7080 15040 -6360
rect 15732 -7080 16452 -6360
rect 17144 -7080 17864 -6360
rect 18556 -7080 19276 -6360
rect 19968 -7080 20688 -6360
rect 21380 -7080 22100 -6360
rect 22792 -7080 23512 -6360
rect -23804 -8200 -23084 -7480
rect -22392 -8200 -21672 -7480
rect -20980 -8200 -20260 -7480
rect -19568 -8200 -18848 -7480
rect -18156 -8200 -17436 -7480
rect -16744 -8200 -16024 -7480
rect -15332 -8200 -14612 -7480
rect -13920 -8200 -13200 -7480
rect -12508 -8200 -11788 -7480
rect -11096 -8200 -10376 -7480
rect -9684 -8200 -8964 -7480
rect -8272 -8200 -7552 -7480
rect -6860 -8200 -6140 -7480
rect -5448 -8200 -4728 -7480
rect -4036 -8200 -3316 -7480
rect -2624 -8200 -1904 -7480
rect -1212 -8200 -492 -7480
rect 200 -8200 920 -7480
rect 1612 -8200 2332 -7480
rect 3024 -8200 3744 -7480
rect 4436 -8200 5156 -7480
rect 5848 -8200 6568 -7480
rect 7260 -8200 7980 -7480
rect 8672 -8200 9392 -7480
rect 10084 -8200 10804 -7480
rect 11496 -8200 12216 -7480
rect 12908 -8200 13628 -7480
rect 14320 -8200 15040 -7480
rect 15732 -8200 16452 -7480
rect 17144 -8200 17864 -7480
rect 18556 -8200 19276 -7480
rect 19968 -8200 20688 -7480
rect 21380 -8200 22100 -7480
rect 22792 -8200 23512 -7480
rect -23804 -9320 -23084 -8600
rect -22392 -9320 -21672 -8600
rect -20980 -9320 -20260 -8600
rect -19568 -9320 -18848 -8600
rect -18156 -9320 -17436 -8600
rect -16744 -9320 -16024 -8600
rect -15332 -9320 -14612 -8600
rect -13920 -9320 -13200 -8600
rect -12508 -9320 -11788 -8600
rect -11096 -9320 -10376 -8600
rect -9684 -9320 -8964 -8600
rect -8272 -9320 -7552 -8600
rect -6860 -9320 -6140 -8600
rect -5448 -9320 -4728 -8600
rect -4036 -9320 -3316 -8600
rect -2624 -9320 -1904 -8600
rect -1212 -9320 -492 -8600
rect 200 -9320 920 -8600
rect 1612 -9320 2332 -8600
rect 3024 -9320 3744 -8600
rect 4436 -9320 5156 -8600
rect 5848 -9320 6568 -8600
rect 7260 -9320 7980 -8600
rect 8672 -9320 9392 -8600
rect 10084 -9320 10804 -8600
rect 11496 -9320 12216 -8600
rect 12908 -9320 13628 -8600
rect 14320 -9320 15040 -8600
rect 15732 -9320 16452 -8600
rect 17144 -9320 17864 -8600
rect 18556 -9320 19276 -8600
rect 19968 -9320 20688 -8600
rect 21380 -9320 22100 -8600
rect 22792 -9320 23512 -8600
rect -23804 -10440 -23084 -9720
rect -22392 -10440 -21672 -9720
rect -20980 -10440 -20260 -9720
rect -19568 -10440 -18848 -9720
rect -18156 -10440 -17436 -9720
rect -16744 -10440 -16024 -9720
rect -15332 -10440 -14612 -9720
rect -13920 -10440 -13200 -9720
rect -12508 -10440 -11788 -9720
rect -11096 -10440 -10376 -9720
rect -9684 -10440 -8964 -9720
rect -8272 -10440 -7552 -9720
rect -6860 -10440 -6140 -9720
rect -5448 -10440 -4728 -9720
rect -4036 -10440 -3316 -9720
rect -2624 -10440 -1904 -9720
rect -1212 -10440 -492 -9720
rect 200 -10440 920 -9720
rect 1612 -10440 2332 -9720
rect 3024 -10440 3744 -9720
rect 4436 -10440 5156 -9720
rect 5848 -10440 6568 -9720
rect 7260 -10440 7980 -9720
rect 8672 -10440 9392 -9720
rect 10084 -10440 10804 -9720
rect 11496 -10440 12216 -9720
rect 12908 -10440 13628 -9720
rect 14320 -10440 15040 -9720
rect 15732 -10440 16452 -9720
rect 17144 -10440 17864 -9720
rect 18556 -10440 19276 -9720
rect 19968 -10440 20688 -9720
rect 21380 -10440 22100 -9720
rect 22792 -10440 23512 -9720
rect -23804 -11560 -23084 -10840
rect -22392 -11560 -21672 -10840
rect -20980 -11560 -20260 -10840
rect -19568 -11560 -18848 -10840
rect -18156 -11560 -17436 -10840
rect -16744 -11560 -16024 -10840
rect -15332 -11560 -14612 -10840
rect -13920 -11560 -13200 -10840
rect -12508 -11560 -11788 -10840
rect -11096 -11560 -10376 -10840
rect -9684 -11560 -8964 -10840
rect -8272 -11560 -7552 -10840
rect -6860 -11560 -6140 -10840
rect -5448 -11560 -4728 -10840
rect -4036 -11560 -3316 -10840
rect -2624 -11560 -1904 -10840
rect -1212 -11560 -492 -10840
rect 200 -11560 920 -10840
rect 1612 -11560 2332 -10840
rect 3024 -11560 3744 -10840
rect 4436 -11560 5156 -10840
rect 5848 -11560 6568 -10840
rect 7260 -11560 7980 -10840
rect 8672 -11560 9392 -10840
rect 10084 -11560 10804 -10840
rect 11496 -11560 12216 -10840
rect 12908 -11560 13628 -10840
rect 14320 -11560 15040 -10840
rect 15732 -11560 16452 -10840
rect 17144 -11560 17864 -10840
rect 18556 -11560 19276 -10840
rect 19968 -11560 20688 -10840
rect 21380 -11560 22100 -10840
rect 22792 -11560 23512 -10840
rect -23804 -12680 -23084 -11960
rect -22392 -12680 -21672 -11960
rect -20980 -12680 -20260 -11960
rect -19568 -12680 -18848 -11960
rect -18156 -12680 -17436 -11960
rect -16744 -12680 -16024 -11960
rect -15332 -12680 -14612 -11960
rect -13920 -12680 -13200 -11960
rect -12508 -12680 -11788 -11960
rect -11096 -12680 -10376 -11960
rect -9684 -12680 -8964 -11960
rect -8272 -12680 -7552 -11960
rect -6860 -12680 -6140 -11960
rect -5448 -12680 -4728 -11960
rect -4036 -12680 -3316 -11960
rect -2624 -12680 -1904 -11960
rect -1212 -12680 -492 -11960
rect 200 -12680 920 -11960
rect 1612 -12680 2332 -11960
rect 3024 -12680 3744 -11960
rect 4436 -12680 5156 -11960
rect 5848 -12680 6568 -11960
rect 7260 -12680 7980 -11960
rect 8672 -12680 9392 -11960
rect 10084 -12680 10804 -11960
rect 11496 -12680 12216 -11960
rect 12908 -12680 13628 -11960
rect 14320 -12680 15040 -11960
rect 15732 -12680 16452 -11960
rect 17144 -12680 17864 -11960
rect 18556 -12680 19276 -11960
rect 19968 -12680 20688 -11960
rect 21380 -12680 22100 -11960
rect 22792 -12680 23512 -11960
rect -23804 -13800 -23084 -13080
rect -22392 -13800 -21672 -13080
rect -20980 -13800 -20260 -13080
rect -19568 -13800 -18848 -13080
rect -18156 -13800 -17436 -13080
rect -16744 -13800 -16024 -13080
rect -15332 -13800 -14612 -13080
rect -13920 -13800 -13200 -13080
rect -12508 -13800 -11788 -13080
rect -11096 -13800 -10376 -13080
rect -9684 -13800 -8964 -13080
rect -8272 -13800 -7552 -13080
rect -6860 -13800 -6140 -13080
rect -5448 -13800 -4728 -13080
rect -4036 -13800 -3316 -13080
rect -2624 -13800 -1904 -13080
rect -1212 -13800 -492 -13080
rect 200 -13800 920 -13080
rect 1612 -13800 2332 -13080
rect 3024 -13800 3744 -13080
rect 4436 -13800 5156 -13080
rect 5848 -13800 6568 -13080
rect 7260 -13800 7980 -13080
rect 8672 -13800 9392 -13080
rect 10084 -13800 10804 -13080
rect 11496 -13800 12216 -13080
rect 12908 -13800 13628 -13080
rect 14320 -13800 15040 -13080
rect 15732 -13800 16452 -13080
rect 17144 -13800 17864 -13080
rect 18556 -13800 19276 -13080
rect 19968 -13800 20688 -13080
rect 21380 -13800 22100 -13080
rect 22792 -13800 23512 -13080
rect -23804 -14920 -23084 -14200
rect -22392 -14920 -21672 -14200
rect -20980 -14920 -20260 -14200
rect -19568 -14920 -18848 -14200
rect -18156 -14920 -17436 -14200
rect -16744 -14920 -16024 -14200
rect -15332 -14920 -14612 -14200
rect -13920 -14920 -13200 -14200
rect -12508 -14920 -11788 -14200
rect -11096 -14920 -10376 -14200
rect -9684 -14920 -8964 -14200
rect -8272 -14920 -7552 -14200
rect -6860 -14920 -6140 -14200
rect -5448 -14920 -4728 -14200
rect -4036 -14920 -3316 -14200
rect -2624 -14920 -1904 -14200
rect -1212 -14920 -492 -14200
rect 200 -14920 920 -14200
rect 1612 -14920 2332 -14200
rect 3024 -14920 3744 -14200
rect 4436 -14920 5156 -14200
rect 5848 -14920 6568 -14200
rect 7260 -14920 7980 -14200
rect 8672 -14920 9392 -14200
rect 10084 -14920 10804 -14200
rect 11496 -14920 12216 -14200
rect 12908 -14920 13628 -14200
rect 14320 -14920 15040 -14200
rect 15732 -14920 16452 -14200
rect 17144 -14920 17864 -14200
rect 18556 -14920 19276 -14200
rect 19968 -14920 20688 -14200
rect 21380 -14920 22100 -14200
rect 22792 -14920 23512 -14200
rect -23804 -16040 -23084 -15320
rect -22392 -16040 -21672 -15320
rect -20980 -16040 -20260 -15320
rect -19568 -16040 -18848 -15320
rect -18156 -16040 -17436 -15320
rect -16744 -16040 -16024 -15320
rect -15332 -16040 -14612 -15320
rect -13920 -16040 -13200 -15320
rect -12508 -16040 -11788 -15320
rect -11096 -16040 -10376 -15320
rect -9684 -16040 -8964 -15320
rect -8272 -16040 -7552 -15320
rect -6860 -16040 -6140 -15320
rect -5448 -16040 -4728 -15320
rect -4036 -16040 -3316 -15320
rect -2624 -16040 -1904 -15320
rect -1212 -16040 -492 -15320
rect 200 -16040 920 -15320
rect 1612 -16040 2332 -15320
rect 3024 -16040 3744 -15320
rect 4436 -16040 5156 -15320
rect 5848 -16040 6568 -15320
rect 7260 -16040 7980 -15320
rect 8672 -16040 9392 -15320
rect 10084 -16040 10804 -15320
rect 11496 -16040 12216 -15320
rect 12908 -16040 13628 -15320
rect 14320 -16040 15040 -15320
rect 15732 -16040 16452 -15320
rect 17144 -16040 17864 -15320
rect 18556 -16040 19276 -15320
rect 19968 -16040 20688 -15320
rect 21380 -16040 22100 -15320
rect 22792 -16040 23512 -15320
rect -23804 -17160 -23084 -16440
rect -22392 -17160 -21672 -16440
rect -20980 -17160 -20260 -16440
rect -19568 -17160 -18848 -16440
rect -18156 -17160 -17436 -16440
rect -16744 -17160 -16024 -16440
rect -15332 -17160 -14612 -16440
rect -13920 -17160 -13200 -16440
rect -12508 -17160 -11788 -16440
rect -11096 -17160 -10376 -16440
rect -9684 -17160 -8964 -16440
rect -8272 -17160 -7552 -16440
rect -6860 -17160 -6140 -16440
rect -5448 -17160 -4728 -16440
rect -4036 -17160 -3316 -16440
rect -2624 -17160 -1904 -16440
rect -1212 -17160 -492 -16440
rect 200 -17160 920 -16440
rect 1612 -17160 2332 -16440
rect 3024 -17160 3744 -16440
rect 4436 -17160 5156 -16440
rect 5848 -17160 6568 -16440
rect 7260 -17160 7980 -16440
rect 8672 -17160 9392 -16440
rect 10084 -17160 10804 -16440
rect 11496 -17160 12216 -16440
rect 12908 -17160 13628 -16440
rect 14320 -17160 15040 -16440
rect 15732 -17160 16452 -16440
rect 17144 -17160 17864 -16440
rect 18556 -17160 19276 -16440
rect 19968 -17160 20688 -16440
rect 21380 -17160 22100 -16440
rect 22792 -17160 23512 -16440
rect -23804 -18280 -23084 -17560
rect -22392 -18280 -21672 -17560
rect -20980 -18280 -20260 -17560
rect -19568 -18280 -18848 -17560
rect -18156 -18280 -17436 -17560
rect -16744 -18280 -16024 -17560
rect -15332 -18280 -14612 -17560
rect -13920 -18280 -13200 -17560
rect -12508 -18280 -11788 -17560
rect -11096 -18280 -10376 -17560
rect -9684 -18280 -8964 -17560
rect -8272 -18280 -7552 -17560
rect -6860 -18280 -6140 -17560
rect -5448 -18280 -4728 -17560
rect -4036 -18280 -3316 -17560
rect -2624 -18280 -1904 -17560
rect -1212 -18280 -492 -17560
rect 200 -18280 920 -17560
rect 1612 -18280 2332 -17560
rect 3024 -18280 3744 -17560
rect 4436 -18280 5156 -17560
rect 5848 -18280 6568 -17560
rect 7260 -18280 7980 -17560
rect 8672 -18280 9392 -17560
rect 10084 -18280 10804 -17560
rect 11496 -18280 12216 -17560
rect 12908 -18280 13628 -17560
rect 14320 -18280 15040 -17560
rect 15732 -18280 16452 -17560
rect 17144 -18280 17864 -17560
rect 18556 -18280 19276 -17560
rect 19968 -18280 20688 -17560
rect 21380 -18280 22100 -17560
rect 22792 -18280 23512 -17560
<< metal4 >>
rect -22812 18332 -22716 18348
rect -23805 18280 -23083 18281
rect -23805 17560 -23804 18280
rect -23084 17560 -23083 18280
rect -23805 17559 -23083 17560
rect -22812 17508 -22796 18332
rect -22732 17508 -22716 18332
rect -21400 18332 -21304 18348
rect -22393 18280 -21671 18281
rect -22393 17560 -22392 18280
rect -21672 17560 -21671 18280
rect -22393 17559 -21671 17560
rect -22812 17492 -22716 17508
rect -21400 17508 -21384 18332
rect -21320 17508 -21304 18332
rect -19988 18332 -19892 18348
rect -20981 18280 -20259 18281
rect -20981 17560 -20980 18280
rect -20260 17560 -20259 18280
rect -20981 17559 -20259 17560
rect -21400 17492 -21304 17508
rect -19988 17508 -19972 18332
rect -19908 17508 -19892 18332
rect -18576 18332 -18480 18348
rect -19569 18280 -18847 18281
rect -19569 17560 -19568 18280
rect -18848 17560 -18847 18280
rect -19569 17559 -18847 17560
rect -19988 17492 -19892 17508
rect -18576 17508 -18560 18332
rect -18496 17508 -18480 18332
rect -17164 18332 -17068 18348
rect -18157 18280 -17435 18281
rect -18157 17560 -18156 18280
rect -17436 17560 -17435 18280
rect -18157 17559 -17435 17560
rect -18576 17492 -18480 17508
rect -17164 17508 -17148 18332
rect -17084 17508 -17068 18332
rect -15752 18332 -15656 18348
rect -16745 18280 -16023 18281
rect -16745 17560 -16744 18280
rect -16024 17560 -16023 18280
rect -16745 17559 -16023 17560
rect -17164 17492 -17068 17508
rect -15752 17508 -15736 18332
rect -15672 17508 -15656 18332
rect -14340 18332 -14244 18348
rect -15333 18280 -14611 18281
rect -15333 17560 -15332 18280
rect -14612 17560 -14611 18280
rect -15333 17559 -14611 17560
rect -15752 17492 -15656 17508
rect -14340 17508 -14324 18332
rect -14260 17508 -14244 18332
rect -12928 18332 -12832 18348
rect -13921 18280 -13199 18281
rect -13921 17560 -13920 18280
rect -13200 17560 -13199 18280
rect -13921 17559 -13199 17560
rect -14340 17492 -14244 17508
rect -12928 17508 -12912 18332
rect -12848 17508 -12832 18332
rect -11516 18332 -11420 18348
rect -12509 18280 -11787 18281
rect -12509 17560 -12508 18280
rect -11788 17560 -11787 18280
rect -12509 17559 -11787 17560
rect -12928 17492 -12832 17508
rect -11516 17508 -11500 18332
rect -11436 17508 -11420 18332
rect -10104 18332 -10008 18348
rect -11097 18280 -10375 18281
rect -11097 17560 -11096 18280
rect -10376 17560 -10375 18280
rect -11097 17559 -10375 17560
rect -11516 17492 -11420 17508
rect -10104 17508 -10088 18332
rect -10024 17508 -10008 18332
rect -8692 18332 -8596 18348
rect -9685 18280 -8963 18281
rect -9685 17560 -9684 18280
rect -8964 17560 -8963 18280
rect -9685 17559 -8963 17560
rect -10104 17492 -10008 17508
rect -8692 17508 -8676 18332
rect -8612 17508 -8596 18332
rect -7280 18332 -7184 18348
rect -8273 18280 -7551 18281
rect -8273 17560 -8272 18280
rect -7552 17560 -7551 18280
rect -8273 17559 -7551 17560
rect -8692 17492 -8596 17508
rect -7280 17508 -7264 18332
rect -7200 17508 -7184 18332
rect -5868 18332 -5772 18348
rect -6861 18280 -6139 18281
rect -6861 17560 -6860 18280
rect -6140 17560 -6139 18280
rect -6861 17559 -6139 17560
rect -7280 17492 -7184 17508
rect -5868 17508 -5852 18332
rect -5788 17508 -5772 18332
rect -4456 18332 -4360 18348
rect -5449 18280 -4727 18281
rect -5449 17560 -5448 18280
rect -4728 17560 -4727 18280
rect -5449 17559 -4727 17560
rect -5868 17492 -5772 17508
rect -4456 17508 -4440 18332
rect -4376 17508 -4360 18332
rect -3044 18332 -2948 18348
rect -4037 18280 -3315 18281
rect -4037 17560 -4036 18280
rect -3316 17560 -3315 18280
rect -4037 17559 -3315 17560
rect -4456 17492 -4360 17508
rect -3044 17508 -3028 18332
rect -2964 17508 -2948 18332
rect -1632 18332 -1536 18348
rect -2625 18280 -1903 18281
rect -2625 17560 -2624 18280
rect -1904 17560 -1903 18280
rect -2625 17559 -1903 17560
rect -3044 17492 -2948 17508
rect -1632 17508 -1616 18332
rect -1552 17508 -1536 18332
rect -220 18332 -124 18348
rect -1213 18280 -491 18281
rect -1213 17560 -1212 18280
rect -492 17560 -491 18280
rect -1213 17559 -491 17560
rect -1632 17492 -1536 17508
rect -220 17508 -204 18332
rect -140 17508 -124 18332
rect 1192 18332 1288 18348
rect 199 18280 921 18281
rect 199 17560 200 18280
rect 920 17560 921 18280
rect 199 17559 921 17560
rect -220 17492 -124 17508
rect 1192 17508 1208 18332
rect 1272 17508 1288 18332
rect 2604 18332 2700 18348
rect 1611 18280 2333 18281
rect 1611 17560 1612 18280
rect 2332 17560 2333 18280
rect 1611 17559 2333 17560
rect 1192 17492 1288 17508
rect 2604 17508 2620 18332
rect 2684 17508 2700 18332
rect 4016 18332 4112 18348
rect 3023 18280 3745 18281
rect 3023 17560 3024 18280
rect 3744 17560 3745 18280
rect 3023 17559 3745 17560
rect 2604 17492 2700 17508
rect 4016 17508 4032 18332
rect 4096 17508 4112 18332
rect 5428 18332 5524 18348
rect 4435 18280 5157 18281
rect 4435 17560 4436 18280
rect 5156 17560 5157 18280
rect 4435 17559 5157 17560
rect 4016 17492 4112 17508
rect 5428 17508 5444 18332
rect 5508 17508 5524 18332
rect 6840 18332 6936 18348
rect 5847 18280 6569 18281
rect 5847 17560 5848 18280
rect 6568 17560 6569 18280
rect 5847 17559 6569 17560
rect 5428 17492 5524 17508
rect 6840 17508 6856 18332
rect 6920 17508 6936 18332
rect 8252 18332 8348 18348
rect 7259 18280 7981 18281
rect 7259 17560 7260 18280
rect 7980 17560 7981 18280
rect 7259 17559 7981 17560
rect 6840 17492 6936 17508
rect 8252 17508 8268 18332
rect 8332 17508 8348 18332
rect 9664 18332 9760 18348
rect 8671 18280 9393 18281
rect 8671 17560 8672 18280
rect 9392 17560 9393 18280
rect 8671 17559 9393 17560
rect 8252 17492 8348 17508
rect 9664 17508 9680 18332
rect 9744 17508 9760 18332
rect 11076 18332 11172 18348
rect 10083 18280 10805 18281
rect 10083 17560 10084 18280
rect 10804 17560 10805 18280
rect 10083 17559 10805 17560
rect 9664 17492 9760 17508
rect 11076 17508 11092 18332
rect 11156 17508 11172 18332
rect 12488 18332 12584 18348
rect 11495 18280 12217 18281
rect 11495 17560 11496 18280
rect 12216 17560 12217 18280
rect 11495 17559 12217 17560
rect 11076 17492 11172 17508
rect 12488 17508 12504 18332
rect 12568 17508 12584 18332
rect 13900 18332 13996 18348
rect 12907 18280 13629 18281
rect 12907 17560 12908 18280
rect 13628 17560 13629 18280
rect 12907 17559 13629 17560
rect 12488 17492 12584 17508
rect 13900 17508 13916 18332
rect 13980 17508 13996 18332
rect 15312 18332 15408 18348
rect 14319 18280 15041 18281
rect 14319 17560 14320 18280
rect 15040 17560 15041 18280
rect 14319 17559 15041 17560
rect 13900 17492 13996 17508
rect 15312 17508 15328 18332
rect 15392 17508 15408 18332
rect 16724 18332 16820 18348
rect 15731 18280 16453 18281
rect 15731 17560 15732 18280
rect 16452 17560 16453 18280
rect 15731 17559 16453 17560
rect 15312 17492 15408 17508
rect 16724 17508 16740 18332
rect 16804 17508 16820 18332
rect 18136 18332 18232 18348
rect 17143 18280 17865 18281
rect 17143 17560 17144 18280
rect 17864 17560 17865 18280
rect 17143 17559 17865 17560
rect 16724 17492 16820 17508
rect 18136 17508 18152 18332
rect 18216 17508 18232 18332
rect 19548 18332 19644 18348
rect 18555 18280 19277 18281
rect 18555 17560 18556 18280
rect 19276 17560 19277 18280
rect 18555 17559 19277 17560
rect 18136 17492 18232 17508
rect 19548 17508 19564 18332
rect 19628 17508 19644 18332
rect 20960 18332 21056 18348
rect 19967 18280 20689 18281
rect 19967 17560 19968 18280
rect 20688 17560 20689 18280
rect 19967 17559 20689 17560
rect 19548 17492 19644 17508
rect 20960 17508 20976 18332
rect 21040 17508 21056 18332
rect 22372 18332 22468 18348
rect 21379 18280 22101 18281
rect 21379 17560 21380 18280
rect 22100 17560 22101 18280
rect 21379 17559 22101 17560
rect 20960 17492 21056 17508
rect 22372 17508 22388 18332
rect 22452 17508 22468 18332
rect 23784 18332 23880 18348
rect 22791 18280 23513 18281
rect 22791 17560 22792 18280
rect 23512 17560 23513 18280
rect 22791 17559 23513 17560
rect 22372 17492 22468 17508
rect 23784 17508 23800 18332
rect 23864 17508 23880 18332
rect 23784 17492 23880 17508
rect -22812 17212 -22716 17228
rect -23805 17160 -23083 17161
rect -23805 16440 -23804 17160
rect -23084 16440 -23083 17160
rect -23805 16439 -23083 16440
rect -22812 16388 -22796 17212
rect -22732 16388 -22716 17212
rect -21400 17212 -21304 17228
rect -22393 17160 -21671 17161
rect -22393 16440 -22392 17160
rect -21672 16440 -21671 17160
rect -22393 16439 -21671 16440
rect -22812 16372 -22716 16388
rect -21400 16388 -21384 17212
rect -21320 16388 -21304 17212
rect -19988 17212 -19892 17228
rect -20981 17160 -20259 17161
rect -20981 16440 -20980 17160
rect -20260 16440 -20259 17160
rect -20981 16439 -20259 16440
rect -21400 16372 -21304 16388
rect -19988 16388 -19972 17212
rect -19908 16388 -19892 17212
rect -18576 17212 -18480 17228
rect -19569 17160 -18847 17161
rect -19569 16440 -19568 17160
rect -18848 16440 -18847 17160
rect -19569 16439 -18847 16440
rect -19988 16372 -19892 16388
rect -18576 16388 -18560 17212
rect -18496 16388 -18480 17212
rect -17164 17212 -17068 17228
rect -18157 17160 -17435 17161
rect -18157 16440 -18156 17160
rect -17436 16440 -17435 17160
rect -18157 16439 -17435 16440
rect -18576 16372 -18480 16388
rect -17164 16388 -17148 17212
rect -17084 16388 -17068 17212
rect -15752 17212 -15656 17228
rect -16745 17160 -16023 17161
rect -16745 16440 -16744 17160
rect -16024 16440 -16023 17160
rect -16745 16439 -16023 16440
rect -17164 16372 -17068 16388
rect -15752 16388 -15736 17212
rect -15672 16388 -15656 17212
rect -14340 17212 -14244 17228
rect -15333 17160 -14611 17161
rect -15333 16440 -15332 17160
rect -14612 16440 -14611 17160
rect -15333 16439 -14611 16440
rect -15752 16372 -15656 16388
rect -14340 16388 -14324 17212
rect -14260 16388 -14244 17212
rect -12928 17212 -12832 17228
rect -13921 17160 -13199 17161
rect -13921 16440 -13920 17160
rect -13200 16440 -13199 17160
rect -13921 16439 -13199 16440
rect -14340 16372 -14244 16388
rect -12928 16388 -12912 17212
rect -12848 16388 -12832 17212
rect -11516 17212 -11420 17228
rect -12509 17160 -11787 17161
rect -12509 16440 -12508 17160
rect -11788 16440 -11787 17160
rect -12509 16439 -11787 16440
rect -12928 16372 -12832 16388
rect -11516 16388 -11500 17212
rect -11436 16388 -11420 17212
rect -10104 17212 -10008 17228
rect -11097 17160 -10375 17161
rect -11097 16440 -11096 17160
rect -10376 16440 -10375 17160
rect -11097 16439 -10375 16440
rect -11516 16372 -11420 16388
rect -10104 16388 -10088 17212
rect -10024 16388 -10008 17212
rect -8692 17212 -8596 17228
rect -9685 17160 -8963 17161
rect -9685 16440 -9684 17160
rect -8964 16440 -8963 17160
rect -9685 16439 -8963 16440
rect -10104 16372 -10008 16388
rect -8692 16388 -8676 17212
rect -8612 16388 -8596 17212
rect -7280 17212 -7184 17228
rect -8273 17160 -7551 17161
rect -8273 16440 -8272 17160
rect -7552 16440 -7551 17160
rect -8273 16439 -7551 16440
rect -8692 16372 -8596 16388
rect -7280 16388 -7264 17212
rect -7200 16388 -7184 17212
rect -5868 17212 -5772 17228
rect -6861 17160 -6139 17161
rect -6861 16440 -6860 17160
rect -6140 16440 -6139 17160
rect -6861 16439 -6139 16440
rect -7280 16372 -7184 16388
rect -5868 16388 -5852 17212
rect -5788 16388 -5772 17212
rect -4456 17212 -4360 17228
rect -5449 17160 -4727 17161
rect -5449 16440 -5448 17160
rect -4728 16440 -4727 17160
rect -5449 16439 -4727 16440
rect -5868 16372 -5772 16388
rect -4456 16388 -4440 17212
rect -4376 16388 -4360 17212
rect -3044 17212 -2948 17228
rect -4037 17160 -3315 17161
rect -4037 16440 -4036 17160
rect -3316 16440 -3315 17160
rect -4037 16439 -3315 16440
rect -4456 16372 -4360 16388
rect -3044 16388 -3028 17212
rect -2964 16388 -2948 17212
rect -1632 17212 -1536 17228
rect -2625 17160 -1903 17161
rect -2625 16440 -2624 17160
rect -1904 16440 -1903 17160
rect -2625 16439 -1903 16440
rect -3044 16372 -2948 16388
rect -1632 16388 -1616 17212
rect -1552 16388 -1536 17212
rect -220 17212 -124 17228
rect -1213 17160 -491 17161
rect -1213 16440 -1212 17160
rect -492 16440 -491 17160
rect -1213 16439 -491 16440
rect -1632 16372 -1536 16388
rect -220 16388 -204 17212
rect -140 16388 -124 17212
rect 1192 17212 1288 17228
rect 199 17160 921 17161
rect 199 16440 200 17160
rect 920 16440 921 17160
rect 199 16439 921 16440
rect -220 16372 -124 16388
rect 1192 16388 1208 17212
rect 1272 16388 1288 17212
rect 2604 17212 2700 17228
rect 1611 17160 2333 17161
rect 1611 16440 1612 17160
rect 2332 16440 2333 17160
rect 1611 16439 2333 16440
rect 1192 16372 1288 16388
rect 2604 16388 2620 17212
rect 2684 16388 2700 17212
rect 4016 17212 4112 17228
rect 3023 17160 3745 17161
rect 3023 16440 3024 17160
rect 3744 16440 3745 17160
rect 3023 16439 3745 16440
rect 2604 16372 2700 16388
rect 4016 16388 4032 17212
rect 4096 16388 4112 17212
rect 5428 17212 5524 17228
rect 4435 17160 5157 17161
rect 4435 16440 4436 17160
rect 5156 16440 5157 17160
rect 4435 16439 5157 16440
rect 4016 16372 4112 16388
rect 5428 16388 5444 17212
rect 5508 16388 5524 17212
rect 6840 17212 6936 17228
rect 5847 17160 6569 17161
rect 5847 16440 5848 17160
rect 6568 16440 6569 17160
rect 5847 16439 6569 16440
rect 5428 16372 5524 16388
rect 6840 16388 6856 17212
rect 6920 16388 6936 17212
rect 8252 17212 8348 17228
rect 7259 17160 7981 17161
rect 7259 16440 7260 17160
rect 7980 16440 7981 17160
rect 7259 16439 7981 16440
rect 6840 16372 6936 16388
rect 8252 16388 8268 17212
rect 8332 16388 8348 17212
rect 9664 17212 9760 17228
rect 8671 17160 9393 17161
rect 8671 16440 8672 17160
rect 9392 16440 9393 17160
rect 8671 16439 9393 16440
rect 8252 16372 8348 16388
rect 9664 16388 9680 17212
rect 9744 16388 9760 17212
rect 11076 17212 11172 17228
rect 10083 17160 10805 17161
rect 10083 16440 10084 17160
rect 10804 16440 10805 17160
rect 10083 16439 10805 16440
rect 9664 16372 9760 16388
rect 11076 16388 11092 17212
rect 11156 16388 11172 17212
rect 12488 17212 12584 17228
rect 11495 17160 12217 17161
rect 11495 16440 11496 17160
rect 12216 16440 12217 17160
rect 11495 16439 12217 16440
rect 11076 16372 11172 16388
rect 12488 16388 12504 17212
rect 12568 16388 12584 17212
rect 13900 17212 13996 17228
rect 12907 17160 13629 17161
rect 12907 16440 12908 17160
rect 13628 16440 13629 17160
rect 12907 16439 13629 16440
rect 12488 16372 12584 16388
rect 13900 16388 13916 17212
rect 13980 16388 13996 17212
rect 15312 17212 15408 17228
rect 14319 17160 15041 17161
rect 14319 16440 14320 17160
rect 15040 16440 15041 17160
rect 14319 16439 15041 16440
rect 13900 16372 13996 16388
rect 15312 16388 15328 17212
rect 15392 16388 15408 17212
rect 16724 17212 16820 17228
rect 15731 17160 16453 17161
rect 15731 16440 15732 17160
rect 16452 16440 16453 17160
rect 15731 16439 16453 16440
rect 15312 16372 15408 16388
rect 16724 16388 16740 17212
rect 16804 16388 16820 17212
rect 18136 17212 18232 17228
rect 17143 17160 17865 17161
rect 17143 16440 17144 17160
rect 17864 16440 17865 17160
rect 17143 16439 17865 16440
rect 16724 16372 16820 16388
rect 18136 16388 18152 17212
rect 18216 16388 18232 17212
rect 19548 17212 19644 17228
rect 18555 17160 19277 17161
rect 18555 16440 18556 17160
rect 19276 16440 19277 17160
rect 18555 16439 19277 16440
rect 18136 16372 18232 16388
rect 19548 16388 19564 17212
rect 19628 16388 19644 17212
rect 20960 17212 21056 17228
rect 19967 17160 20689 17161
rect 19967 16440 19968 17160
rect 20688 16440 20689 17160
rect 19967 16439 20689 16440
rect 19548 16372 19644 16388
rect 20960 16388 20976 17212
rect 21040 16388 21056 17212
rect 22372 17212 22468 17228
rect 21379 17160 22101 17161
rect 21379 16440 21380 17160
rect 22100 16440 22101 17160
rect 21379 16439 22101 16440
rect 20960 16372 21056 16388
rect 22372 16388 22388 17212
rect 22452 16388 22468 17212
rect 23784 17212 23880 17228
rect 22791 17160 23513 17161
rect 22791 16440 22792 17160
rect 23512 16440 23513 17160
rect 22791 16439 23513 16440
rect 22372 16372 22468 16388
rect 23784 16388 23800 17212
rect 23864 16388 23880 17212
rect 23784 16372 23880 16388
rect -22812 16092 -22716 16108
rect -23805 16040 -23083 16041
rect -23805 15320 -23804 16040
rect -23084 15320 -23083 16040
rect -23805 15319 -23083 15320
rect -22812 15268 -22796 16092
rect -22732 15268 -22716 16092
rect -21400 16092 -21304 16108
rect -22393 16040 -21671 16041
rect -22393 15320 -22392 16040
rect -21672 15320 -21671 16040
rect -22393 15319 -21671 15320
rect -22812 15252 -22716 15268
rect -21400 15268 -21384 16092
rect -21320 15268 -21304 16092
rect -19988 16092 -19892 16108
rect -20981 16040 -20259 16041
rect -20981 15320 -20980 16040
rect -20260 15320 -20259 16040
rect -20981 15319 -20259 15320
rect -21400 15252 -21304 15268
rect -19988 15268 -19972 16092
rect -19908 15268 -19892 16092
rect -18576 16092 -18480 16108
rect -19569 16040 -18847 16041
rect -19569 15320 -19568 16040
rect -18848 15320 -18847 16040
rect -19569 15319 -18847 15320
rect -19988 15252 -19892 15268
rect -18576 15268 -18560 16092
rect -18496 15268 -18480 16092
rect -17164 16092 -17068 16108
rect -18157 16040 -17435 16041
rect -18157 15320 -18156 16040
rect -17436 15320 -17435 16040
rect -18157 15319 -17435 15320
rect -18576 15252 -18480 15268
rect -17164 15268 -17148 16092
rect -17084 15268 -17068 16092
rect -15752 16092 -15656 16108
rect -16745 16040 -16023 16041
rect -16745 15320 -16744 16040
rect -16024 15320 -16023 16040
rect -16745 15319 -16023 15320
rect -17164 15252 -17068 15268
rect -15752 15268 -15736 16092
rect -15672 15268 -15656 16092
rect -14340 16092 -14244 16108
rect -15333 16040 -14611 16041
rect -15333 15320 -15332 16040
rect -14612 15320 -14611 16040
rect -15333 15319 -14611 15320
rect -15752 15252 -15656 15268
rect -14340 15268 -14324 16092
rect -14260 15268 -14244 16092
rect -12928 16092 -12832 16108
rect -13921 16040 -13199 16041
rect -13921 15320 -13920 16040
rect -13200 15320 -13199 16040
rect -13921 15319 -13199 15320
rect -14340 15252 -14244 15268
rect -12928 15268 -12912 16092
rect -12848 15268 -12832 16092
rect -11516 16092 -11420 16108
rect -12509 16040 -11787 16041
rect -12509 15320 -12508 16040
rect -11788 15320 -11787 16040
rect -12509 15319 -11787 15320
rect -12928 15252 -12832 15268
rect -11516 15268 -11500 16092
rect -11436 15268 -11420 16092
rect -10104 16092 -10008 16108
rect -11097 16040 -10375 16041
rect -11097 15320 -11096 16040
rect -10376 15320 -10375 16040
rect -11097 15319 -10375 15320
rect -11516 15252 -11420 15268
rect -10104 15268 -10088 16092
rect -10024 15268 -10008 16092
rect -8692 16092 -8596 16108
rect -9685 16040 -8963 16041
rect -9685 15320 -9684 16040
rect -8964 15320 -8963 16040
rect -9685 15319 -8963 15320
rect -10104 15252 -10008 15268
rect -8692 15268 -8676 16092
rect -8612 15268 -8596 16092
rect -7280 16092 -7184 16108
rect -8273 16040 -7551 16041
rect -8273 15320 -8272 16040
rect -7552 15320 -7551 16040
rect -8273 15319 -7551 15320
rect -8692 15252 -8596 15268
rect -7280 15268 -7264 16092
rect -7200 15268 -7184 16092
rect -5868 16092 -5772 16108
rect -6861 16040 -6139 16041
rect -6861 15320 -6860 16040
rect -6140 15320 -6139 16040
rect -6861 15319 -6139 15320
rect -7280 15252 -7184 15268
rect -5868 15268 -5852 16092
rect -5788 15268 -5772 16092
rect -4456 16092 -4360 16108
rect -5449 16040 -4727 16041
rect -5449 15320 -5448 16040
rect -4728 15320 -4727 16040
rect -5449 15319 -4727 15320
rect -5868 15252 -5772 15268
rect -4456 15268 -4440 16092
rect -4376 15268 -4360 16092
rect -3044 16092 -2948 16108
rect -4037 16040 -3315 16041
rect -4037 15320 -4036 16040
rect -3316 15320 -3315 16040
rect -4037 15319 -3315 15320
rect -4456 15252 -4360 15268
rect -3044 15268 -3028 16092
rect -2964 15268 -2948 16092
rect -1632 16092 -1536 16108
rect -2625 16040 -1903 16041
rect -2625 15320 -2624 16040
rect -1904 15320 -1903 16040
rect -2625 15319 -1903 15320
rect -3044 15252 -2948 15268
rect -1632 15268 -1616 16092
rect -1552 15268 -1536 16092
rect -220 16092 -124 16108
rect -1213 16040 -491 16041
rect -1213 15320 -1212 16040
rect -492 15320 -491 16040
rect -1213 15319 -491 15320
rect -1632 15252 -1536 15268
rect -220 15268 -204 16092
rect -140 15268 -124 16092
rect 1192 16092 1288 16108
rect 199 16040 921 16041
rect 199 15320 200 16040
rect 920 15320 921 16040
rect 199 15319 921 15320
rect -220 15252 -124 15268
rect 1192 15268 1208 16092
rect 1272 15268 1288 16092
rect 2604 16092 2700 16108
rect 1611 16040 2333 16041
rect 1611 15320 1612 16040
rect 2332 15320 2333 16040
rect 1611 15319 2333 15320
rect 1192 15252 1288 15268
rect 2604 15268 2620 16092
rect 2684 15268 2700 16092
rect 4016 16092 4112 16108
rect 3023 16040 3745 16041
rect 3023 15320 3024 16040
rect 3744 15320 3745 16040
rect 3023 15319 3745 15320
rect 2604 15252 2700 15268
rect 4016 15268 4032 16092
rect 4096 15268 4112 16092
rect 5428 16092 5524 16108
rect 4435 16040 5157 16041
rect 4435 15320 4436 16040
rect 5156 15320 5157 16040
rect 4435 15319 5157 15320
rect 4016 15252 4112 15268
rect 5428 15268 5444 16092
rect 5508 15268 5524 16092
rect 6840 16092 6936 16108
rect 5847 16040 6569 16041
rect 5847 15320 5848 16040
rect 6568 15320 6569 16040
rect 5847 15319 6569 15320
rect 5428 15252 5524 15268
rect 6840 15268 6856 16092
rect 6920 15268 6936 16092
rect 8252 16092 8348 16108
rect 7259 16040 7981 16041
rect 7259 15320 7260 16040
rect 7980 15320 7981 16040
rect 7259 15319 7981 15320
rect 6840 15252 6936 15268
rect 8252 15268 8268 16092
rect 8332 15268 8348 16092
rect 9664 16092 9760 16108
rect 8671 16040 9393 16041
rect 8671 15320 8672 16040
rect 9392 15320 9393 16040
rect 8671 15319 9393 15320
rect 8252 15252 8348 15268
rect 9664 15268 9680 16092
rect 9744 15268 9760 16092
rect 11076 16092 11172 16108
rect 10083 16040 10805 16041
rect 10083 15320 10084 16040
rect 10804 15320 10805 16040
rect 10083 15319 10805 15320
rect 9664 15252 9760 15268
rect 11076 15268 11092 16092
rect 11156 15268 11172 16092
rect 12488 16092 12584 16108
rect 11495 16040 12217 16041
rect 11495 15320 11496 16040
rect 12216 15320 12217 16040
rect 11495 15319 12217 15320
rect 11076 15252 11172 15268
rect 12488 15268 12504 16092
rect 12568 15268 12584 16092
rect 13900 16092 13996 16108
rect 12907 16040 13629 16041
rect 12907 15320 12908 16040
rect 13628 15320 13629 16040
rect 12907 15319 13629 15320
rect 12488 15252 12584 15268
rect 13900 15268 13916 16092
rect 13980 15268 13996 16092
rect 15312 16092 15408 16108
rect 14319 16040 15041 16041
rect 14319 15320 14320 16040
rect 15040 15320 15041 16040
rect 14319 15319 15041 15320
rect 13900 15252 13996 15268
rect 15312 15268 15328 16092
rect 15392 15268 15408 16092
rect 16724 16092 16820 16108
rect 15731 16040 16453 16041
rect 15731 15320 15732 16040
rect 16452 15320 16453 16040
rect 15731 15319 16453 15320
rect 15312 15252 15408 15268
rect 16724 15268 16740 16092
rect 16804 15268 16820 16092
rect 18136 16092 18232 16108
rect 17143 16040 17865 16041
rect 17143 15320 17144 16040
rect 17864 15320 17865 16040
rect 17143 15319 17865 15320
rect 16724 15252 16820 15268
rect 18136 15268 18152 16092
rect 18216 15268 18232 16092
rect 19548 16092 19644 16108
rect 18555 16040 19277 16041
rect 18555 15320 18556 16040
rect 19276 15320 19277 16040
rect 18555 15319 19277 15320
rect 18136 15252 18232 15268
rect 19548 15268 19564 16092
rect 19628 15268 19644 16092
rect 20960 16092 21056 16108
rect 19967 16040 20689 16041
rect 19967 15320 19968 16040
rect 20688 15320 20689 16040
rect 19967 15319 20689 15320
rect 19548 15252 19644 15268
rect 20960 15268 20976 16092
rect 21040 15268 21056 16092
rect 22372 16092 22468 16108
rect 21379 16040 22101 16041
rect 21379 15320 21380 16040
rect 22100 15320 22101 16040
rect 21379 15319 22101 15320
rect 20960 15252 21056 15268
rect 22372 15268 22388 16092
rect 22452 15268 22468 16092
rect 23784 16092 23880 16108
rect 22791 16040 23513 16041
rect 22791 15320 22792 16040
rect 23512 15320 23513 16040
rect 22791 15319 23513 15320
rect 22372 15252 22468 15268
rect 23784 15268 23800 16092
rect 23864 15268 23880 16092
rect 23784 15252 23880 15268
rect -22812 14972 -22716 14988
rect -23805 14920 -23083 14921
rect -23805 14200 -23804 14920
rect -23084 14200 -23083 14920
rect -23805 14199 -23083 14200
rect -22812 14148 -22796 14972
rect -22732 14148 -22716 14972
rect -21400 14972 -21304 14988
rect -22393 14920 -21671 14921
rect -22393 14200 -22392 14920
rect -21672 14200 -21671 14920
rect -22393 14199 -21671 14200
rect -22812 14132 -22716 14148
rect -21400 14148 -21384 14972
rect -21320 14148 -21304 14972
rect -19988 14972 -19892 14988
rect -20981 14920 -20259 14921
rect -20981 14200 -20980 14920
rect -20260 14200 -20259 14920
rect -20981 14199 -20259 14200
rect -21400 14132 -21304 14148
rect -19988 14148 -19972 14972
rect -19908 14148 -19892 14972
rect -18576 14972 -18480 14988
rect -19569 14920 -18847 14921
rect -19569 14200 -19568 14920
rect -18848 14200 -18847 14920
rect -19569 14199 -18847 14200
rect -19988 14132 -19892 14148
rect -18576 14148 -18560 14972
rect -18496 14148 -18480 14972
rect -17164 14972 -17068 14988
rect -18157 14920 -17435 14921
rect -18157 14200 -18156 14920
rect -17436 14200 -17435 14920
rect -18157 14199 -17435 14200
rect -18576 14132 -18480 14148
rect -17164 14148 -17148 14972
rect -17084 14148 -17068 14972
rect -15752 14972 -15656 14988
rect -16745 14920 -16023 14921
rect -16745 14200 -16744 14920
rect -16024 14200 -16023 14920
rect -16745 14199 -16023 14200
rect -17164 14132 -17068 14148
rect -15752 14148 -15736 14972
rect -15672 14148 -15656 14972
rect -14340 14972 -14244 14988
rect -15333 14920 -14611 14921
rect -15333 14200 -15332 14920
rect -14612 14200 -14611 14920
rect -15333 14199 -14611 14200
rect -15752 14132 -15656 14148
rect -14340 14148 -14324 14972
rect -14260 14148 -14244 14972
rect -12928 14972 -12832 14988
rect -13921 14920 -13199 14921
rect -13921 14200 -13920 14920
rect -13200 14200 -13199 14920
rect -13921 14199 -13199 14200
rect -14340 14132 -14244 14148
rect -12928 14148 -12912 14972
rect -12848 14148 -12832 14972
rect -11516 14972 -11420 14988
rect -12509 14920 -11787 14921
rect -12509 14200 -12508 14920
rect -11788 14200 -11787 14920
rect -12509 14199 -11787 14200
rect -12928 14132 -12832 14148
rect -11516 14148 -11500 14972
rect -11436 14148 -11420 14972
rect -10104 14972 -10008 14988
rect -11097 14920 -10375 14921
rect -11097 14200 -11096 14920
rect -10376 14200 -10375 14920
rect -11097 14199 -10375 14200
rect -11516 14132 -11420 14148
rect -10104 14148 -10088 14972
rect -10024 14148 -10008 14972
rect -8692 14972 -8596 14988
rect -9685 14920 -8963 14921
rect -9685 14200 -9684 14920
rect -8964 14200 -8963 14920
rect -9685 14199 -8963 14200
rect -10104 14132 -10008 14148
rect -8692 14148 -8676 14972
rect -8612 14148 -8596 14972
rect -7280 14972 -7184 14988
rect -8273 14920 -7551 14921
rect -8273 14200 -8272 14920
rect -7552 14200 -7551 14920
rect -8273 14199 -7551 14200
rect -8692 14132 -8596 14148
rect -7280 14148 -7264 14972
rect -7200 14148 -7184 14972
rect -5868 14972 -5772 14988
rect -6861 14920 -6139 14921
rect -6861 14200 -6860 14920
rect -6140 14200 -6139 14920
rect -6861 14199 -6139 14200
rect -7280 14132 -7184 14148
rect -5868 14148 -5852 14972
rect -5788 14148 -5772 14972
rect -4456 14972 -4360 14988
rect -5449 14920 -4727 14921
rect -5449 14200 -5448 14920
rect -4728 14200 -4727 14920
rect -5449 14199 -4727 14200
rect -5868 14132 -5772 14148
rect -4456 14148 -4440 14972
rect -4376 14148 -4360 14972
rect -3044 14972 -2948 14988
rect -4037 14920 -3315 14921
rect -4037 14200 -4036 14920
rect -3316 14200 -3315 14920
rect -4037 14199 -3315 14200
rect -4456 14132 -4360 14148
rect -3044 14148 -3028 14972
rect -2964 14148 -2948 14972
rect -1632 14972 -1536 14988
rect -2625 14920 -1903 14921
rect -2625 14200 -2624 14920
rect -1904 14200 -1903 14920
rect -2625 14199 -1903 14200
rect -3044 14132 -2948 14148
rect -1632 14148 -1616 14972
rect -1552 14148 -1536 14972
rect -220 14972 -124 14988
rect -1213 14920 -491 14921
rect -1213 14200 -1212 14920
rect -492 14200 -491 14920
rect -1213 14199 -491 14200
rect -1632 14132 -1536 14148
rect -220 14148 -204 14972
rect -140 14148 -124 14972
rect 1192 14972 1288 14988
rect 199 14920 921 14921
rect 199 14200 200 14920
rect 920 14200 921 14920
rect 199 14199 921 14200
rect -220 14132 -124 14148
rect 1192 14148 1208 14972
rect 1272 14148 1288 14972
rect 2604 14972 2700 14988
rect 1611 14920 2333 14921
rect 1611 14200 1612 14920
rect 2332 14200 2333 14920
rect 1611 14199 2333 14200
rect 1192 14132 1288 14148
rect 2604 14148 2620 14972
rect 2684 14148 2700 14972
rect 4016 14972 4112 14988
rect 3023 14920 3745 14921
rect 3023 14200 3024 14920
rect 3744 14200 3745 14920
rect 3023 14199 3745 14200
rect 2604 14132 2700 14148
rect 4016 14148 4032 14972
rect 4096 14148 4112 14972
rect 5428 14972 5524 14988
rect 4435 14920 5157 14921
rect 4435 14200 4436 14920
rect 5156 14200 5157 14920
rect 4435 14199 5157 14200
rect 4016 14132 4112 14148
rect 5428 14148 5444 14972
rect 5508 14148 5524 14972
rect 6840 14972 6936 14988
rect 5847 14920 6569 14921
rect 5847 14200 5848 14920
rect 6568 14200 6569 14920
rect 5847 14199 6569 14200
rect 5428 14132 5524 14148
rect 6840 14148 6856 14972
rect 6920 14148 6936 14972
rect 8252 14972 8348 14988
rect 7259 14920 7981 14921
rect 7259 14200 7260 14920
rect 7980 14200 7981 14920
rect 7259 14199 7981 14200
rect 6840 14132 6936 14148
rect 8252 14148 8268 14972
rect 8332 14148 8348 14972
rect 9664 14972 9760 14988
rect 8671 14920 9393 14921
rect 8671 14200 8672 14920
rect 9392 14200 9393 14920
rect 8671 14199 9393 14200
rect 8252 14132 8348 14148
rect 9664 14148 9680 14972
rect 9744 14148 9760 14972
rect 11076 14972 11172 14988
rect 10083 14920 10805 14921
rect 10083 14200 10084 14920
rect 10804 14200 10805 14920
rect 10083 14199 10805 14200
rect 9664 14132 9760 14148
rect 11076 14148 11092 14972
rect 11156 14148 11172 14972
rect 12488 14972 12584 14988
rect 11495 14920 12217 14921
rect 11495 14200 11496 14920
rect 12216 14200 12217 14920
rect 11495 14199 12217 14200
rect 11076 14132 11172 14148
rect 12488 14148 12504 14972
rect 12568 14148 12584 14972
rect 13900 14972 13996 14988
rect 12907 14920 13629 14921
rect 12907 14200 12908 14920
rect 13628 14200 13629 14920
rect 12907 14199 13629 14200
rect 12488 14132 12584 14148
rect 13900 14148 13916 14972
rect 13980 14148 13996 14972
rect 15312 14972 15408 14988
rect 14319 14920 15041 14921
rect 14319 14200 14320 14920
rect 15040 14200 15041 14920
rect 14319 14199 15041 14200
rect 13900 14132 13996 14148
rect 15312 14148 15328 14972
rect 15392 14148 15408 14972
rect 16724 14972 16820 14988
rect 15731 14920 16453 14921
rect 15731 14200 15732 14920
rect 16452 14200 16453 14920
rect 15731 14199 16453 14200
rect 15312 14132 15408 14148
rect 16724 14148 16740 14972
rect 16804 14148 16820 14972
rect 18136 14972 18232 14988
rect 17143 14920 17865 14921
rect 17143 14200 17144 14920
rect 17864 14200 17865 14920
rect 17143 14199 17865 14200
rect 16724 14132 16820 14148
rect 18136 14148 18152 14972
rect 18216 14148 18232 14972
rect 19548 14972 19644 14988
rect 18555 14920 19277 14921
rect 18555 14200 18556 14920
rect 19276 14200 19277 14920
rect 18555 14199 19277 14200
rect 18136 14132 18232 14148
rect 19548 14148 19564 14972
rect 19628 14148 19644 14972
rect 20960 14972 21056 14988
rect 19967 14920 20689 14921
rect 19967 14200 19968 14920
rect 20688 14200 20689 14920
rect 19967 14199 20689 14200
rect 19548 14132 19644 14148
rect 20960 14148 20976 14972
rect 21040 14148 21056 14972
rect 22372 14972 22468 14988
rect 21379 14920 22101 14921
rect 21379 14200 21380 14920
rect 22100 14200 22101 14920
rect 21379 14199 22101 14200
rect 20960 14132 21056 14148
rect 22372 14148 22388 14972
rect 22452 14148 22468 14972
rect 23784 14972 23880 14988
rect 22791 14920 23513 14921
rect 22791 14200 22792 14920
rect 23512 14200 23513 14920
rect 22791 14199 23513 14200
rect 22372 14132 22468 14148
rect 23784 14148 23800 14972
rect 23864 14148 23880 14972
rect 23784 14132 23880 14148
rect -22812 13852 -22716 13868
rect -23805 13800 -23083 13801
rect -23805 13080 -23804 13800
rect -23084 13080 -23083 13800
rect -23805 13079 -23083 13080
rect -22812 13028 -22796 13852
rect -22732 13028 -22716 13852
rect -21400 13852 -21304 13868
rect -22393 13800 -21671 13801
rect -22393 13080 -22392 13800
rect -21672 13080 -21671 13800
rect -22393 13079 -21671 13080
rect -22812 13012 -22716 13028
rect -21400 13028 -21384 13852
rect -21320 13028 -21304 13852
rect -19988 13852 -19892 13868
rect -20981 13800 -20259 13801
rect -20981 13080 -20980 13800
rect -20260 13080 -20259 13800
rect -20981 13079 -20259 13080
rect -21400 13012 -21304 13028
rect -19988 13028 -19972 13852
rect -19908 13028 -19892 13852
rect -18576 13852 -18480 13868
rect -19569 13800 -18847 13801
rect -19569 13080 -19568 13800
rect -18848 13080 -18847 13800
rect -19569 13079 -18847 13080
rect -19988 13012 -19892 13028
rect -18576 13028 -18560 13852
rect -18496 13028 -18480 13852
rect -17164 13852 -17068 13868
rect -18157 13800 -17435 13801
rect -18157 13080 -18156 13800
rect -17436 13080 -17435 13800
rect -18157 13079 -17435 13080
rect -18576 13012 -18480 13028
rect -17164 13028 -17148 13852
rect -17084 13028 -17068 13852
rect -15752 13852 -15656 13868
rect -16745 13800 -16023 13801
rect -16745 13080 -16744 13800
rect -16024 13080 -16023 13800
rect -16745 13079 -16023 13080
rect -17164 13012 -17068 13028
rect -15752 13028 -15736 13852
rect -15672 13028 -15656 13852
rect -14340 13852 -14244 13868
rect -15333 13800 -14611 13801
rect -15333 13080 -15332 13800
rect -14612 13080 -14611 13800
rect -15333 13079 -14611 13080
rect -15752 13012 -15656 13028
rect -14340 13028 -14324 13852
rect -14260 13028 -14244 13852
rect -12928 13852 -12832 13868
rect -13921 13800 -13199 13801
rect -13921 13080 -13920 13800
rect -13200 13080 -13199 13800
rect -13921 13079 -13199 13080
rect -14340 13012 -14244 13028
rect -12928 13028 -12912 13852
rect -12848 13028 -12832 13852
rect -11516 13852 -11420 13868
rect -12509 13800 -11787 13801
rect -12509 13080 -12508 13800
rect -11788 13080 -11787 13800
rect -12509 13079 -11787 13080
rect -12928 13012 -12832 13028
rect -11516 13028 -11500 13852
rect -11436 13028 -11420 13852
rect -10104 13852 -10008 13868
rect -11097 13800 -10375 13801
rect -11097 13080 -11096 13800
rect -10376 13080 -10375 13800
rect -11097 13079 -10375 13080
rect -11516 13012 -11420 13028
rect -10104 13028 -10088 13852
rect -10024 13028 -10008 13852
rect -8692 13852 -8596 13868
rect -9685 13800 -8963 13801
rect -9685 13080 -9684 13800
rect -8964 13080 -8963 13800
rect -9685 13079 -8963 13080
rect -10104 13012 -10008 13028
rect -8692 13028 -8676 13852
rect -8612 13028 -8596 13852
rect -7280 13852 -7184 13868
rect -8273 13800 -7551 13801
rect -8273 13080 -8272 13800
rect -7552 13080 -7551 13800
rect -8273 13079 -7551 13080
rect -8692 13012 -8596 13028
rect -7280 13028 -7264 13852
rect -7200 13028 -7184 13852
rect -5868 13852 -5772 13868
rect -6861 13800 -6139 13801
rect -6861 13080 -6860 13800
rect -6140 13080 -6139 13800
rect -6861 13079 -6139 13080
rect -7280 13012 -7184 13028
rect -5868 13028 -5852 13852
rect -5788 13028 -5772 13852
rect -4456 13852 -4360 13868
rect -5449 13800 -4727 13801
rect -5449 13080 -5448 13800
rect -4728 13080 -4727 13800
rect -5449 13079 -4727 13080
rect -5868 13012 -5772 13028
rect -4456 13028 -4440 13852
rect -4376 13028 -4360 13852
rect -3044 13852 -2948 13868
rect -4037 13800 -3315 13801
rect -4037 13080 -4036 13800
rect -3316 13080 -3315 13800
rect -4037 13079 -3315 13080
rect -4456 13012 -4360 13028
rect -3044 13028 -3028 13852
rect -2964 13028 -2948 13852
rect -1632 13852 -1536 13868
rect -2625 13800 -1903 13801
rect -2625 13080 -2624 13800
rect -1904 13080 -1903 13800
rect -2625 13079 -1903 13080
rect -3044 13012 -2948 13028
rect -1632 13028 -1616 13852
rect -1552 13028 -1536 13852
rect -220 13852 -124 13868
rect -1213 13800 -491 13801
rect -1213 13080 -1212 13800
rect -492 13080 -491 13800
rect -1213 13079 -491 13080
rect -1632 13012 -1536 13028
rect -220 13028 -204 13852
rect -140 13028 -124 13852
rect 1192 13852 1288 13868
rect 199 13800 921 13801
rect 199 13080 200 13800
rect 920 13080 921 13800
rect 199 13079 921 13080
rect -220 13012 -124 13028
rect 1192 13028 1208 13852
rect 1272 13028 1288 13852
rect 2604 13852 2700 13868
rect 1611 13800 2333 13801
rect 1611 13080 1612 13800
rect 2332 13080 2333 13800
rect 1611 13079 2333 13080
rect 1192 13012 1288 13028
rect 2604 13028 2620 13852
rect 2684 13028 2700 13852
rect 4016 13852 4112 13868
rect 3023 13800 3745 13801
rect 3023 13080 3024 13800
rect 3744 13080 3745 13800
rect 3023 13079 3745 13080
rect 2604 13012 2700 13028
rect 4016 13028 4032 13852
rect 4096 13028 4112 13852
rect 5428 13852 5524 13868
rect 4435 13800 5157 13801
rect 4435 13080 4436 13800
rect 5156 13080 5157 13800
rect 4435 13079 5157 13080
rect 4016 13012 4112 13028
rect 5428 13028 5444 13852
rect 5508 13028 5524 13852
rect 6840 13852 6936 13868
rect 5847 13800 6569 13801
rect 5847 13080 5848 13800
rect 6568 13080 6569 13800
rect 5847 13079 6569 13080
rect 5428 13012 5524 13028
rect 6840 13028 6856 13852
rect 6920 13028 6936 13852
rect 8252 13852 8348 13868
rect 7259 13800 7981 13801
rect 7259 13080 7260 13800
rect 7980 13080 7981 13800
rect 7259 13079 7981 13080
rect 6840 13012 6936 13028
rect 8252 13028 8268 13852
rect 8332 13028 8348 13852
rect 9664 13852 9760 13868
rect 8671 13800 9393 13801
rect 8671 13080 8672 13800
rect 9392 13080 9393 13800
rect 8671 13079 9393 13080
rect 8252 13012 8348 13028
rect 9664 13028 9680 13852
rect 9744 13028 9760 13852
rect 11076 13852 11172 13868
rect 10083 13800 10805 13801
rect 10083 13080 10084 13800
rect 10804 13080 10805 13800
rect 10083 13079 10805 13080
rect 9664 13012 9760 13028
rect 11076 13028 11092 13852
rect 11156 13028 11172 13852
rect 12488 13852 12584 13868
rect 11495 13800 12217 13801
rect 11495 13080 11496 13800
rect 12216 13080 12217 13800
rect 11495 13079 12217 13080
rect 11076 13012 11172 13028
rect 12488 13028 12504 13852
rect 12568 13028 12584 13852
rect 13900 13852 13996 13868
rect 12907 13800 13629 13801
rect 12907 13080 12908 13800
rect 13628 13080 13629 13800
rect 12907 13079 13629 13080
rect 12488 13012 12584 13028
rect 13900 13028 13916 13852
rect 13980 13028 13996 13852
rect 15312 13852 15408 13868
rect 14319 13800 15041 13801
rect 14319 13080 14320 13800
rect 15040 13080 15041 13800
rect 14319 13079 15041 13080
rect 13900 13012 13996 13028
rect 15312 13028 15328 13852
rect 15392 13028 15408 13852
rect 16724 13852 16820 13868
rect 15731 13800 16453 13801
rect 15731 13080 15732 13800
rect 16452 13080 16453 13800
rect 15731 13079 16453 13080
rect 15312 13012 15408 13028
rect 16724 13028 16740 13852
rect 16804 13028 16820 13852
rect 18136 13852 18232 13868
rect 17143 13800 17865 13801
rect 17143 13080 17144 13800
rect 17864 13080 17865 13800
rect 17143 13079 17865 13080
rect 16724 13012 16820 13028
rect 18136 13028 18152 13852
rect 18216 13028 18232 13852
rect 19548 13852 19644 13868
rect 18555 13800 19277 13801
rect 18555 13080 18556 13800
rect 19276 13080 19277 13800
rect 18555 13079 19277 13080
rect 18136 13012 18232 13028
rect 19548 13028 19564 13852
rect 19628 13028 19644 13852
rect 20960 13852 21056 13868
rect 19967 13800 20689 13801
rect 19967 13080 19968 13800
rect 20688 13080 20689 13800
rect 19967 13079 20689 13080
rect 19548 13012 19644 13028
rect 20960 13028 20976 13852
rect 21040 13028 21056 13852
rect 22372 13852 22468 13868
rect 21379 13800 22101 13801
rect 21379 13080 21380 13800
rect 22100 13080 22101 13800
rect 21379 13079 22101 13080
rect 20960 13012 21056 13028
rect 22372 13028 22388 13852
rect 22452 13028 22468 13852
rect 23784 13852 23880 13868
rect 22791 13800 23513 13801
rect 22791 13080 22792 13800
rect 23512 13080 23513 13800
rect 22791 13079 23513 13080
rect 22372 13012 22468 13028
rect 23784 13028 23800 13852
rect 23864 13028 23880 13852
rect 23784 13012 23880 13028
rect -22812 12732 -22716 12748
rect -23805 12680 -23083 12681
rect -23805 11960 -23804 12680
rect -23084 11960 -23083 12680
rect -23805 11959 -23083 11960
rect -22812 11908 -22796 12732
rect -22732 11908 -22716 12732
rect -21400 12732 -21304 12748
rect -22393 12680 -21671 12681
rect -22393 11960 -22392 12680
rect -21672 11960 -21671 12680
rect -22393 11959 -21671 11960
rect -22812 11892 -22716 11908
rect -21400 11908 -21384 12732
rect -21320 11908 -21304 12732
rect -19988 12732 -19892 12748
rect -20981 12680 -20259 12681
rect -20981 11960 -20980 12680
rect -20260 11960 -20259 12680
rect -20981 11959 -20259 11960
rect -21400 11892 -21304 11908
rect -19988 11908 -19972 12732
rect -19908 11908 -19892 12732
rect -18576 12732 -18480 12748
rect -19569 12680 -18847 12681
rect -19569 11960 -19568 12680
rect -18848 11960 -18847 12680
rect -19569 11959 -18847 11960
rect -19988 11892 -19892 11908
rect -18576 11908 -18560 12732
rect -18496 11908 -18480 12732
rect -17164 12732 -17068 12748
rect -18157 12680 -17435 12681
rect -18157 11960 -18156 12680
rect -17436 11960 -17435 12680
rect -18157 11959 -17435 11960
rect -18576 11892 -18480 11908
rect -17164 11908 -17148 12732
rect -17084 11908 -17068 12732
rect -15752 12732 -15656 12748
rect -16745 12680 -16023 12681
rect -16745 11960 -16744 12680
rect -16024 11960 -16023 12680
rect -16745 11959 -16023 11960
rect -17164 11892 -17068 11908
rect -15752 11908 -15736 12732
rect -15672 11908 -15656 12732
rect -14340 12732 -14244 12748
rect -15333 12680 -14611 12681
rect -15333 11960 -15332 12680
rect -14612 11960 -14611 12680
rect -15333 11959 -14611 11960
rect -15752 11892 -15656 11908
rect -14340 11908 -14324 12732
rect -14260 11908 -14244 12732
rect -12928 12732 -12832 12748
rect -13921 12680 -13199 12681
rect -13921 11960 -13920 12680
rect -13200 11960 -13199 12680
rect -13921 11959 -13199 11960
rect -14340 11892 -14244 11908
rect -12928 11908 -12912 12732
rect -12848 11908 -12832 12732
rect -11516 12732 -11420 12748
rect -12509 12680 -11787 12681
rect -12509 11960 -12508 12680
rect -11788 11960 -11787 12680
rect -12509 11959 -11787 11960
rect -12928 11892 -12832 11908
rect -11516 11908 -11500 12732
rect -11436 11908 -11420 12732
rect -10104 12732 -10008 12748
rect -11097 12680 -10375 12681
rect -11097 11960 -11096 12680
rect -10376 11960 -10375 12680
rect -11097 11959 -10375 11960
rect -11516 11892 -11420 11908
rect -10104 11908 -10088 12732
rect -10024 11908 -10008 12732
rect -8692 12732 -8596 12748
rect -9685 12680 -8963 12681
rect -9685 11960 -9684 12680
rect -8964 11960 -8963 12680
rect -9685 11959 -8963 11960
rect -10104 11892 -10008 11908
rect -8692 11908 -8676 12732
rect -8612 11908 -8596 12732
rect -7280 12732 -7184 12748
rect -8273 12680 -7551 12681
rect -8273 11960 -8272 12680
rect -7552 11960 -7551 12680
rect -8273 11959 -7551 11960
rect -8692 11892 -8596 11908
rect -7280 11908 -7264 12732
rect -7200 11908 -7184 12732
rect -5868 12732 -5772 12748
rect -6861 12680 -6139 12681
rect -6861 11960 -6860 12680
rect -6140 11960 -6139 12680
rect -6861 11959 -6139 11960
rect -7280 11892 -7184 11908
rect -5868 11908 -5852 12732
rect -5788 11908 -5772 12732
rect -4456 12732 -4360 12748
rect -5449 12680 -4727 12681
rect -5449 11960 -5448 12680
rect -4728 11960 -4727 12680
rect -5449 11959 -4727 11960
rect -5868 11892 -5772 11908
rect -4456 11908 -4440 12732
rect -4376 11908 -4360 12732
rect -3044 12732 -2948 12748
rect -4037 12680 -3315 12681
rect -4037 11960 -4036 12680
rect -3316 11960 -3315 12680
rect -4037 11959 -3315 11960
rect -4456 11892 -4360 11908
rect -3044 11908 -3028 12732
rect -2964 11908 -2948 12732
rect -1632 12732 -1536 12748
rect -2625 12680 -1903 12681
rect -2625 11960 -2624 12680
rect -1904 11960 -1903 12680
rect -2625 11959 -1903 11960
rect -3044 11892 -2948 11908
rect -1632 11908 -1616 12732
rect -1552 11908 -1536 12732
rect -220 12732 -124 12748
rect -1213 12680 -491 12681
rect -1213 11960 -1212 12680
rect -492 11960 -491 12680
rect -1213 11959 -491 11960
rect -1632 11892 -1536 11908
rect -220 11908 -204 12732
rect -140 11908 -124 12732
rect 1192 12732 1288 12748
rect 199 12680 921 12681
rect 199 11960 200 12680
rect 920 11960 921 12680
rect 199 11959 921 11960
rect -220 11892 -124 11908
rect 1192 11908 1208 12732
rect 1272 11908 1288 12732
rect 2604 12732 2700 12748
rect 1611 12680 2333 12681
rect 1611 11960 1612 12680
rect 2332 11960 2333 12680
rect 1611 11959 2333 11960
rect 1192 11892 1288 11908
rect 2604 11908 2620 12732
rect 2684 11908 2700 12732
rect 4016 12732 4112 12748
rect 3023 12680 3745 12681
rect 3023 11960 3024 12680
rect 3744 11960 3745 12680
rect 3023 11959 3745 11960
rect 2604 11892 2700 11908
rect 4016 11908 4032 12732
rect 4096 11908 4112 12732
rect 5428 12732 5524 12748
rect 4435 12680 5157 12681
rect 4435 11960 4436 12680
rect 5156 11960 5157 12680
rect 4435 11959 5157 11960
rect 4016 11892 4112 11908
rect 5428 11908 5444 12732
rect 5508 11908 5524 12732
rect 6840 12732 6936 12748
rect 5847 12680 6569 12681
rect 5847 11960 5848 12680
rect 6568 11960 6569 12680
rect 5847 11959 6569 11960
rect 5428 11892 5524 11908
rect 6840 11908 6856 12732
rect 6920 11908 6936 12732
rect 8252 12732 8348 12748
rect 7259 12680 7981 12681
rect 7259 11960 7260 12680
rect 7980 11960 7981 12680
rect 7259 11959 7981 11960
rect 6840 11892 6936 11908
rect 8252 11908 8268 12732
rect 8332 11908 8348 12732
rect 9664 12732 9760 12748
rect 8671 12680 9393 12681
rect 8671 11960 8672 12680
rect 9392 11960 9393 12680
rect 8671 11959 9393 11960
rect 8252 11892 8348 11908
rect 9664 11908 9680 12732
rect 9744 11908 9760 12732
rect 11076 12732 11172 12748
rect 10083 12680 10805 12681
rect 10083 11960 10084 12680
rect 10804 11960 10805 12680
rect 10083 11959 10805 11960
rect 9664 11892 9760 11908
rect 11076 11908 11092 12732
rect 11156 11908 11172 12732
rect 12488 12732 12584 12748
rect 11495 12680 12217 12681
rect 11495 11960 11496 12680
rect 12216 11960 12217 12680
rect 11495 11959 12217 11960
rect 11076 11892 11172 11908
rect 12488 11908 12504 12732
rect 12568 11908 12584 12732
rect 13900 12732 13996 12748
rect 12907 12680 13629 12681
rect 12907 11960 12908 12680
rect 13628 11960 13629 12680
rect 12907 11959 13629 11960
rect 12488 11892 12584 11908
rect 13900 11908 13916 12732
rect 13980 11908 13996 12732
rect 15312 12732 15408 12748
rect 14319 12680 15041 12681
rect 14319 11960 14320 12680
rect 15040 11960 15041 12680
rect 14319 11959 15041 11960
rect 13900 11892 13996 11908
rect 15312 11908 15328 12732
rect 15392 11908 15408 12732
rect 16724 12732 16820 12748
rect 15731 12680 16453 12681
rect 15731 11960 15732 12680
rect 16452 11960 16453 12680
rect 15731 11959 16453 11960
rect 15312 11892 15408 11908
rect 16724 11908 16740 12732
rect 16804 11908 16820 12732
rect 18136 12732 18232 12748
rect 17143 12680 17865 12681
rect 17143 11960 17144 12680
rect 17864 11960 17865 12680
rect 17143 11959 17865 11960
rect 16724 11892 16820 11908
rect 18136 11908 18152 12732
rect 18216 11908 18232 12732
rect 19548 12732 19644 12748
rect 18555 12680 19277 12681
rect 18555 11960 18556 12680
rect 19276 11960 19277 12680
rect 18555 11959 19277 11960
rect 18136 11892 18232 11908
rect 19548 11908 19564 12732
rect 19628 11908 19644 12732
rect 20960 12732 21056 12748
rect 19967 12680 20689 12681
rect 19967 11960 19968 12680
rect 20688 11960 20689 12680
rect 19967 11959 20689 11960
rect 19548 11892 19644 11908
rect 20960 11908 20976 12732
rect 21040 11908 21056 12732
rect 22372 12732 22468 12748
rect 21379 12680 22101 12681
rect 21379 11960 21380 12680
rect 22100 11960 22101 12680
rect 21379 11959 22101 11960
rect 20960 11892 21056 11908
rect 22372 11908 22388 12732
rect 22452 11908 22468 12732
rect 23784 12732 23880 12748
rect 22791 12680 23513 12681
rect 22791 11960 22792 12680
rect 23512 11960 23513 12680
rect 22791 11959 23513 11960
rect 22372 11892 22468 11908
rect 23784 11908 23800 12732
rect 23864 11908 23880 12732
rect 23784 11892 23880 11908
rect -22812 11612 -22716 11628
rect -23805 11560 -23083 11561
rect -23805 10840 -23804 11560
rect -23084 10840 -23083 11560
rect -23805 10839 -23083 10840
rect -22812 10788 -22796 11612
rect -22732 10788 -22716 11612
rect -21400 11612 -21304 11628
rect -22393 11560 -21671 11561
rect -22393 10840 -22392 11560
rect -21672 10840 -21671 11560
rect -22393 10839 -21671 10840
rect -22812 10772 -22716 10788
rect -21400 10788 -21384 11612
rect -21320 10788 -21304 11612
rect -19988 11612 -19892 11628
rect -20981 11560 -20259 11561
rect -20981 10840 -20980 11560
rect -20260 10840 -20259 11560
rect -20981 10839 -20259 10840
rect -21400 10772 -21304 10788
rect -19988 10788 -19972 11612
rect -19908 10788 -19892 11612
rect -18576 11612 -18480 11628
rect -19569 11560 -18847 11561
rect -19569 10840 -19568 11560
rect -18848 10840 -18847 11560
rect -19569 10839 -18847 10840
rect -19988 10772 -19892 10788
rect -18576 10788 -18560 11612
rect -18496 10788 -18480 11612
rect -17164 11612 -17068 11628
rect -18157 11560 -17435 11561
rect -18157 10840 -18156 11560
rect -17436 10840 -17435 11560
rect -18157 10839 -17435 10840
rect -18576 10772 -18480 10788
rect -17164 10788 -17148 11612
rect -17084 10788 -17068 11612
rect -15752 11612 -15656 11628
rect -16745 11560 -16023 11561
rect -16745 10840 -16744 11560
rect -16024 10840 -16023 11560
rect -16745 10839 -16023 10840
rect -17164 10772 -17068 10788
rect -15752 10788 -15736 11612
rect -15672 10788 -15656 11612
rect -14340 11612 -14244 11628
rect -15333 11560 -14611 11561
rect -15333 10840 -15332 11560
rect -14612 10840 -14611 11560
rect -15333 10839 -14611 10840
rect -15752 10772 -15656 10788
rect -14340 10788 -14324 11612
rect -14260 10788 -14244 11612
rect -12928 11612 -12832 11628
rect -13921 11560 -13199 11561
rect -13921 10840 -13920 11560
rect -13200 10840 -13199 11560
rect -13921 10839 -13199 10840
rect -14340 10772 -14244 10788
rect -12928 10788 -12912 11612
rect -12848 10788 -12832 11612
rect -11516 11612 -11420 11628
rect -12509 11560 -11787 11561
rect -12509 10840 -12508 11560
rect -11788 10840 -11787 11560
rect -12509 10839 -11787 10840
rect -12928 10772 -12832 10788
rect -11516 10788 -11500 11612
rect -11436 10788 -11420 11612
rect -10104 11612 -10008 11628
rect -11097 11560 -10375 11561
rect -11097 10840 -11096 11560
rect -10376 10840 -10375 11560
rect -11097 10839 -10375 10840
rect -11516 10772 -11420 10788
rect -10104 10788 -10088 11612
rect -10024 10788 -10008 11612
rect -8692 11612 -8596 11628
rect -9685 11560 -8963 11561
rect -9685 10840 -9684 11560
rect -8964 10840 -8963 11560
rect -9685 10839 -8963 10840
rect -10104 10772 -10008 10788
rect -8692 10788 -8676 11612
rect -8612 10788 -8596 11612
rect -7280 11612 -7184 11628
rect -8273 11560 -7551 11561
rect -8273 10840 -8272 11560
rect -7552 10840 -7551 11560
rect -8273 10839 -7551 10840
rect -8692 10772 -8596 10788
rect -7280 10788 -7264 11612
rect -7200 10788 -7184 11612
rect -5868 11612 -5772 11628
rect -6861 11560 -6139 11561
rect -6861 10840 -6860 11560
rect -6140 10840 -6139 11560
rect -6861 10839 -6139 10840
rect -7280 10772 -7184 10788
rect -5868 10788 -5852 11612
rect -5788 10788 -5772 11612
rect -4456 11612 -4360 11628
rect -5449 11560 -4727 11561
rect -5449 10840 -5448 11560
rect -4728 10840 -4727 11560
rect -5449 10839 -4727 10840
rect -5868 10772 -5772 10788
rect -4456 10788 -4440 11612
rect -4376 10788 -4360 11612
rect -3044 11612 -2948 11628
rect -4037 11560 -3315 11561
rect -4037 10840 -4036 11560
rect -3316 10840 -3315 11560
rect -4037 10839 -3315 10840
rect -4456 10772 -4360 10788
rect -3044 10788 -3028 11612
rect -2964 10788 -2948 11612
rect -1632 11612 -1536 11628
rect -2625 11560 -1903 11561
rect -2625 10840 -2624 11560
rect -1904 10840 -1903 11560
rect -2625 10839 -1903 10840
rect -3044 10772 -2948 10788
rect -1632 10788 -1616 11612
rect -1552 10788 -1536 11612
rect -220 11612 -124 11628
rect -1213 11560 -491 11561
rect -1213 10840 -1212 11560
rect -492 10840 -491 11560
rect -1213 10839 -491 10840
rect -1632 10772 -1536 10788
rect -220 10788 -204 11612
rect -140 10788 -124 11612
rect 1192 11612 1288 11628
rect 199 11560 921 11561
rect 199 10840 200 11560
rect 920 10840 921 11560
rect 199 10839 921 10840
rect -220 10772 -124 10788
rect 1192 10788 1208 11612
rect 1272 10788 1288 11612
rect 2604 11612 2700 11628
rect 1611 11560 2333 11561
rect 1611 10840 1612 11560
rect 2332 10840 2333 11560
rect 1611 10839 2333 10840
rect 1192 10772 1288 10788
rect 2604 10788 2620 11612
rect 2684 10788 2700 11612
rect 4016 11612 4112 11628
rect 3023 11560 3745 11561
rect 3023 10840 3024 11560
rect 3744 10840 3745 11560
rect 3023 10839 3745 10840
rect 2604 10772 2700 10788
rect 4016 10788 4032 11612
rect 4096 10788 4112 11612
rect 5428 11612 5524 11628
rect 4435 11560 5157 11561
rect 4435 10840 4436 11560
rect 5156 10840 5157 11560
rect 4435 10839 5157 10840
rect 4016 10772 4112 10788
rect 5428 10788 5444 11612
rect 5508 10788 5524 11612
rect 6840 11612 6936 11628
rect 5847 11560 6569 11561
rect 5847 10840 5848 11560
rect 6568 10840 6569 11560
rect 5847 10839 6569 10840
rect 5428 10772 5524 10788
rect 6840 10788 6856 11612
rect 6920 10788 6936 11612
rect 8252 11612 8348 11628
rect 7259 11560 7981 11561
rect 7259 10840 7260 11560
rect 7980 10840 7981 11560
rect 7259 10839 7981 10840
rect 6840 10772 6936 10788
rect 8252 10788 8268 11612
rect 8332 10788 8348 11612
rect 9664 11612 9760 11628
rect 8671 11560 9393 11561
rect 8671 10840 8672 11560
rect 9392 10840 9393 11560
rect 8671 10839 9393 10840
rect 8252 10772 8348 10788
rect 9664 10788 9680 11612
rect 9744 10788 9760 11612
rect 11076 11612 11172 11628
rect 10083 11560 10805 11561
rect 10083 10840 10084 11560
rect 10804 10840 10805 11560
rect 10083 10839 10805 10840
rect 9664 10772 9760 10788
rect 11076 10788 11092 11612
rect 11156 10788 11172 11612
rect 12488 11612 12584 11628
rect 11495 11560 12217 11561
rect 11495 10840 11496 11560
rect 12216 10840 12217 11560
rect 11495 10839 12217 10840
rect 11076 10772 11172 10788
rect 12488 10788 12504 11612
rect 12568 10788 12584 11612
rect 13900 11612 13996 11628
rect 12907 11560 13629 11561
rect 12907 10840 12908 11560
rect 13628 10840 13629 11560
rect 12907 10839 13629 10840
rect 12488 10772 12584 10788
rect 13900 10788 13916 11612
rect 13980 10788 13996 11612
rect 15312 11612 15408 11628
rect 14319 11560 15041 11561
rect 14319 10840 14320 11560
rect 15040 10840 15041 11560
rect 14319 10839 15041 10840
rect 13900 10772 13996 10788
rect 15312 10788 15328 11612
rect 15392 10788 15408 11612
rect 16724 11612 16820 11628
rect 15731 11560 16453 11561
rect 15731 10840 15732 11560
rect 16452 10840 16453 11560
rect 15731 10839 16453 10840
rect 15312 10772 15408 10788
rect 16724 10788 16740 11612
rect 16804 10788 16820 11612
rect 18136 11612 18232 11628
rect 17143 11560 17865 11561
rect 17143 10840 17144 11560
rect 17864 10840 17865 11560
rect 17143 10839 17865 10840
rect 16724 10772 16820 10788
rect 18136 10788 18152 11612
rect 18216 10788 18232 11612
rect 19548 11612 19644 11628
rect 18555 11560 19277 11561
rect 18555 10840 18556 11560
rect 19276 10840 19277 11560
rect 18555 10839 19277 10840
rect 18136 10772 18232 10788
rect 19548 10788 19564 11612
rect 19628 10788 19644 11612
rect 20960 11612 21056 11628
rect 19967 11560 20689 11561
rect 19967 10840 19968 11560
rect 20688 10840 20689 11560
rect 19967 10839 20689 10840
rect 19548 10772 19644 10788
rect 20960 10788 20976 11612
rect 21040 10788 21056 11612
rect 22372 11612 22468 11628
rect 21379 11560 22101 11561
rect 21379 10840 21380 11560
rect 22100 10840 22101 11560
rect 21379 10839 22101 10840
rect 20960 10772 21056 10788
rect 22372 10788 22388 11612
rect 22452 10788 22468 11612
rect 23784 11612 23880 11628
rect 22791 11560 23513 11561
rect 22791 10840 22792 11560
rect 23512 10840 23513 11560
rect 22791 10839 23513 10840
rect 22372 10772 22468 10788
rect 23784 10788 23800 11612
rect 23864 10788 23880 11612
rect 23784 10772 23880 10788
rect -22812 10492 -22716 10508
rect -23805 10440 -23083 10441
rect -23805 9720 -23804 10440
rect -23084 9720 -23083 10440
rect -23805 9719 -23083 9720
rect -22812 9668 -22796 10492
rect -22732 9668 -22716 10492
rect -21400 10492 -21304 10508
rect -22393 10440 -21671 10441
rect -22393 9720 -22392 10440
rect -21672 9720 -21671 10440
rect -22393 9719 -21671 9720
rect -22812 9652 -22716 9668
rect -21400 9668 -21384 10492
rect -21320 9668 -21304 10492
rect -19988 10492 -19892 10508
rect -20981 10440 -20259 10441
rect -20981 9720 -20980 10440
rect -20260 9720 -20259 10440
rect -20981 9719 -20259 9720
rect -21400 9652 -21304 9668
rect -19988 9668 -19972 10492
rect -19908 9668 -19892 10492
rect -18576 10492 -18480 10508
rect -19569 10440 -18847 10441
rect -19569 9720 -19568 10440
rect -18848 9720 -18847 10440
rect -19569 9719 -18847 9720
rect -19988 9652 -19892 9668
rect -18576 9668 -18560 10492
rect -18496 9668 -18480 10492
rect -17164 10492 -17068 10508
rect -18157 10440 -17435 10441
rect -18157 9720 -18156 10440
rect -17436 9720 -17435 10440
rect -18157 9719 -17435 9720
rect -18576 9652 -18480 9668
rect -17164 9668 -17148 10492
rect -17084 9668 -17068 10492
rect -15752 10492 -15656 10508
rect -16745 10440 -16023 10441
rect -16745 9720 -16744 10440
rect -16024 9720 -16023 10440
rect -16745 9719 -16023 9720
rect -17164 9652 -17068 9668
rect -15752 9668 -15736 10492
rect -15672 9668 -15656 10492
rect -14340 10492 -14244 10508
rect -15333 10440 -14611 10441
rect -15333 9720 -15332 10440
rect -14612 9720 -14611 10440
rect -15333 9719 -14611 9720
rect -15752 9652 -15656 9668
rect -14340 9668 -14324 10492
rect -14260 9668 -14244 10492
rect -12928 10492 -12832 10508
rect -13921 10440 -13199 10441
rect -13921 9720 -13920 10440
rect -13200 9720 -13199 10440
rect -13921 9719 -13199 9720
rect -14340 9652 -14244 9668
rect -12928 9668 -12912 10492
rect -12848 9668 -12832 10492
rect -11516 10492 -11420 10508
rect -12509 10440 -11787 10441
rect -12509 9720 -12508 10440
rect -11788 9720 -11787 10440
rect -12509 9719 -11787 9720
rect -12928 9652 -12832 9668
rect -11516 9668 -11500 10492
rect -11436 9668 -11420 10492
rect -10104 10492 -10008 10508
rect -11097 10440 -10375 10441
rect -11097 9720 -11096 10440
rect -10376 9720 -10375 10440
rect -11097 9719 -10375 9720
rect -11516 9652 -11420 9668
rect -10104 9668 -10088 10492
rect -10024 9668 -10008 10492
rect -8692 10492 -8596 10508
rect -9685 10440 -8963 10441
rect -9685 9720 -9684 10440
rect -8964 9720 -8963 10440
rect -9685 9719 -8963 9720
rect -10104 9652 -10008 9668
rect -8692 9668 -8676 10492
rect -8612 9668 -8596 10492
rect -7280 10492 -7184 10508
rect -8273 10440 -7551 10441
rect -8273 9720 -8272 10440
rect -7552 9720 -7551 10440
rect -8273 9719 -7551 9720
rect -8692 9652 -8596 9668
rect -7280 9668 -7264 10492
rect -7200 9668 -7184 10492
rect -5868 10492 -5772 10508
rect -6861 10440 -6139 10441
rect -6861 9720 -6860 10440
rect -6140 9720 -6139 10440
rect -6861 9719 -6139 9720
rect -7280 9652 -7184 9668
rect -5868 9668 -5852 10492
rect -5788 9668 -5772 10492
rect -4456 10492 -4360 10508
rect -5449 10440 -4727 10441
rect -5449 9720 -5448 10440
rect -4728 9720 -4727 10440
rect -5449 9719 -4727 9720
rect -5868 9652 -5772 9668
rect -4456 9668 -4440 10492
rect -4376 9668 -4360 10492
rect -3044 10492 -2948 10508
rect -4037 10440 -3315 10441
rect -4037 9720 -4036 10440
rect -3316 9720 -3315 10440
rect -4037 9719 -3315 9720
rect -4456 9652 -4360 9668
rect -3044 9668 -3028 10492
rect -2964 9668 -2948 10492
rect -1632 10492 -1536 10508
rect -2625 10440 -1903 10441
rect -2625 9720 -2624 10440
rect -1904 9720 -1903 10440
rect -2625 9719 -1903 9720
rect -3044 9652 -2948 9668
rect -1632 9668 -1616 10492
rect -1552 9668 -1536 10492
rect -220 10492 -124 10508
rect -1213 10440 -491 10441
rect -1213 9720 -1212 10440
rect -492 9720 -491 10440
rect -1213 9719 -491 9720
rect -1632 9652 -1536 9668
rect -220 9668 -204 10492
rect -140 9668 -124 10492
rect 1192 10492 1288 10508
rect 199 10440 921 10441
rect 199 9720 200 10440
rect 920 9720 921 10440
rect 199 9719 921 9720
rect -220 9652 -124 9668
rect 1192 9668 1208 10492
rect 1272 9668 1288 10492
rect 2604 10492 2700 10508
rect 1611 10440 2333 10441
rect 1611 9720 1612 10440
rect 2332 9720 2333 10440
rect 1611 9719 2333 9720
rect 1192 9652 1288 9668
rect 2604 9668 2620 10492
rect 2684 9668 2700 10492
rect 4016 10492 4112 10508
rect 3023 10440 3745 10441
rect 3023 9720 3024 10440
rect 3744 9720 3745 10440
rect 3023 9719 3745 9720
rect 2604 9652 2700 9668
rect 4016 9668 4032 10492
rect 4096 9668 4112 10492
rect 5428 10492 5524 10508
rect 4435 10440 5157 10441
rect 4435 9720 4436 10440
rect 5156 9720 5157 10440
rect 4435 9719 5157 9720
rect 4016 9652 4112 9668
rect 5428 9668 5444 10492
rect 5508 9668 5524 10492
rect 6840 10492 6936 10508
rect 5847 10440 6569 10441
rect 5847 9720 5848 10440
rect 6568 9720 6569 10440
rect 5847 9719 6569 9720
rect 5428 9652 5524 9668
rect 6840 9668 6856 10492
rect 6920 9668 6936 10492
rect 8252 10492 8348 10508
rect 7259 10440 7981 10441
rect 7259 9720 7260 10440
rect 7980 9720 7981 10440
rect 7259 9719 7981 9720
rect 6840 9652 6936 9668
rect 8252 9668 8268 10492
rect 8332 9668 8348 10492
rect 9664 10492 9760 10508
rect 8671 10440 9393 10441
rect 8671 9720 8672 10440
rect 9392 9720 9393 10440
rect 8671 9719 9393 9720
rect 8252 9652 8348 9668
rect 9664 9668 9680 10492
rect 9744 9668 9760 10492
rect 11076 10492 11172 10508
rect 10083 10440 10805 10441
rect 10083 9720 10084 10440
rect 10804 9720 10805 10440
rect 10083 9719 10805 9720
rect 9664 9652 9760 9668
rect 11076 9668 11092 10492
rect 11156 9668 11172 10492
rect 12488 10492 12584 10508
rect 11495 10440 12217 10441
rect 11495 9720 11496 10440
rect 12216 9720 12217 10440
rect 11495 9719 12217 9720
rect 11076 9652 11172 9668
rect 12488 9668 12504 10492
rect 12568 9668 12584 10492
rect 13900 10492 13996 10508
rect 12907 10440 13629 10441
rect 12907 9720 12908 10440
rect 13628 9720 13629 10440
rect 12907 9719 13629 9720
rect 12488 9652 12584 9668
rect 13900 9668 13916 10492
rect 13980 9668 13996 10492
rect 15312 10492 15408 10508
rect 14319 10440 15041 10441
rect 14319 9720 14320 10440
rect 15040 9720 15041 10440
rect 14319 9719 15041 9720
rect 13900 9652 13996 9668
rect 15312 9668 15328 10492
rect 15392 9668 15408 10492
rect 16724 10492 16820 10508
rect 15731 10440 16453 10441
rect 15731 9720 15732 10440
rect 16452 9720 16453 10440
rect 15731 9719 16453 9720
rect 15312 9652 15408 9668
rect 16724 9668 16740 10492
rect 16804 9668 16820 10492
rect 18136 10492 18232 10508
rect 17143 10440 17865 10441
rect 17143 9720 17144 10440
rect 17864 9720 17865 10440
rect 17143 9719 17865 9720
rect 16724 9652 16820 9668
rect 18136 9668 18152 10492
rect 18216 9668 18232 10492
rect 19548 10492 19644 10508
rect 18555 10440 19277 10441
rect 18555 9720 18556 10440
rect 19276 9720 19277 10440
rect 18555 9719 19277 9720
rect 18136 9652 18232 9668
rect 19548 9668 19564 10492
rect 19628 9668 19644 10492
rect 20960 10492 21056 10508
rect 19967 10440 20689 10441
rect 19967 9720 19968 10440
rect 20688 9720 20689 10440
rect 19967 9719 20689 9720
rect 19548 9652 19644 9668
rect 20960 9668 20976 10492
rect 21040 9668 21056 10492
rect 22372 10492 22468 10508
rect 21379 10440 22101 10441
rect 21379 9720 21380 10440
rect 22100 9720 22101 10440
rect 21379 9719 22101 9720
rect 20960 9652 21056 9668
rect 22372 9668 22388 10492
rect 22452 9668 22468 10492
rect 23784 10492 23880 10508
rect 22791 10440 23513 10441
rect 22791 9720 22792 10440
rect 23512 9720 23513 10440
rect 22791 9719 23513 9720
rect 22372 9652 22468 9668
rect 23784 9668 23800 10492
rect 23864 9668 23880 10492
rect 23784 9652 23880 9668
rect -22812 9372 -22716 9388
rect -23805 9320 -23083 9321
rect -23805 8600 -23804 9320
rect -23084 8600 -23083 9320
rect -23805 8599 -23083 8600
rect -22812 8548 -22796 9372
rect -22732 8548 -22716 9372
rect -21400 9372 -21304 9388
rect -22393 9320 -21671 9321
rect -22393 8600 -22392 9320
rect -21672 8600 -21671 9320
rect -22393 8599 -21671 8600
rect -22812 8532 -22716 8548
rect -21400 8548 -21384 9372
rect -21320 8548 -21304 9372
rect -19988 9372 -19892 9388
rect -20981 9320 -20259 9321
rect -20981 8600 -20980 9320
rect -20260 8600 -20259 9320
rect -20981 8599 -20259 8600
rect -21400 8532 -21304 8548
rect -19988 8548 -19972 9372
rect -19908 8548 -19892 9372
rect -18576 9372 -18480 9388
rect -19569 9320 -18847 9321
rect -19569 8600 -19568 9320
rect -18848 8600 -18847 9320
rect -19569 8599 -18847 8600
rect -19988 8532 -19892 8548
rect -18576 8548 -18560 9372
rect -18496 8548 -18480 9372
rect -17164 9372 -17068 9388
rect -18157 9320 -17435 9321
rect -18157 8600 -18156 9320
rect -17436 8600 -17435 9320
rect -18157 8599 -17435 8600
rect -18576 8532 -18480 8548
rect -17164 8548 -17148 9372
rect -17084 8548 -17068 9372
rect -15752 9372 -15656 9388
rect -16745 9320 -16023 9321
rect -16745 8600 -16744 9320
rect -16024 8600 -16023 9320
rect -16745 8599 -16023 8600
rect -17164 8532 -17068 8548
rect -15752 8548 -15736 9372
rect -15672 8548 -15656 9372
rect -14340 9372 -14244 9388
rect -15333 9320 -14611 9321
rect -15333 8600 -15332 9320
rect -14612 8600 -14611 9320
rect -15333 8599 -14611 8600
rect -15752 8532 -15656 8548
rect -14340 8548 -14324 9372
rect -14260 8548 -14244 9372
rect -12928 9372 -12832 9388
rect -13921 9320 -13199 9321
rect -13921 8600 -13920 9320
rect -13200 8600 -13199 9320
rect -13921 8599 -13199 8600
rect -14340 8532 -14244 8548
rect -12928 8548 -12912 9372
rect -12848 8548 -12832 9372
rect -11516 9372 -11420 9388
rect -12509 9320 -11787 9321
rect -12509 8600 -12508 9320
rect -11788 8600 -11787 9320
rect -12509 8599 -11787 8600
rect -12928 8532 -12832 8548
rect -11516 8548 -11500 9372
rect -11436 8548 -11420 9372
rect -10104 9372 -10008 9388
rect -11097 9320 -10375 9321
rect -11097 8600 -11096 9320
rect -10376 8600 -10375 9320
rect -11097 8599 -10375 8600
rect -11516 8532 -11420 8548
rect -10104 8548 -10088 9372
rect -10024 8548 -10008 9372
rect -8692 9372 -8596 9388
rect -9685 9320 -8963 9321
rect -9685 8600 -9684 9320
rect -8964 8600 -8963 9320
rect -9685 8599 -8963 8600
rect -10104 8532 -10008 8548
rect -8692 8548 -8676 9372
rect -8612 8548 -8596 9372
rect -7280 9372 -7184 9388
rect -8273 9320 -7551 9321
rect -8273 8600 -8272 9320
rect -7552 8600 -7551 9320
rect -8273 8599 -7551 8600
rect -8692 8532 -8596 8548
rect -7280 8548 -7264 9372
rect -7200 8548 -7184 9372
rect -5868 9372 -5772 9388
rect -6861 9320 -6139 9321
rect -6861 8600 -6860 9320
rect -6140 8600 -6139 9320
rect -6861 8599 -6139 8600
rect -7280 8532 -7184 8548
rect -5868 8548 -5852 9372
rect -5788 8548 -5772 9372
rect -4456 9372 -4360 9388
rect -5449 9320 -4727 9321
rect -5449 8600 -5448 9320
rect -4728 8600 -4727 9320
rect -5449 8599 -4727 8600
rect -5868 8532 -5772 8548
rect -4456 8548 -4440 9372
rect -4376 8548 -4360 9372
rect -3044 9372 -2948 9388
rect -4037 9320 -3315 9321
rect -4037 8600 -4036 9320
rect -3316 8600 -3315 9320
rect -4037 8599 -3315 8600
rect -4456 8532 -4360 8548
rect -3044 8548 -3028 9372
rect -2964 8548 -2948 9372
rect -1632 9372 -1536 9388
rect -2625 9320 -1903 9321
rect -2625 8600 -2624 9320
rect -1904 8600 -1903 9320
rect -2625 8599 -1903 8600
rect -3044 8532 -2948 8548
rect -1632 8548 -1616 9372
rect -1552 8548 -1536 9372
rect -220 9372 -124 9388
rect -1213 9320 -491 9321
rect -1213 8600 -1212 9320
rect -492 8600 -491 9320
rect -1213 8599 -491 8600
rect -1632 8532 -1536 8548
rect -220 8548 -204 9372
rect -140 8548 -124 9372
rect 1192 9372 1288 9388
rect 199 9320 921 9321
rect 199 8600 200 9320
rect 920 8600 921 9320
rect 199 8599 921 8600
rect -220 8532 -124 8548
rect 1192 8548 1208 9372
rect 1272 8548 1288 9372
rect 2604 9372 2700 9388
rect 1611 9320 2333 9321
rect 1611 8600 1612 9320
rect 2332 8600 2333 9320
rect 1611 8599 2333 8600
rect 1192 8532 1288 8548
rect 2604 8548 2620 9372
rect 2684 8548 2700 9372
rect 4016 9372 4112 9388
rect 3023 9320 3745 9321
rect 3023 8600 3024 9320
rect 3744 8600 3745 9320
rect 3023 8599 3745 8600
rect 2604 8532 2700 8548
rect 4016 8548 4032 9372
rect 4096 8548 4112 9372
rect 5428 9372 5524 9388
rect 4435 9320 5157 9321
rect 4435 8600 4436 9320
rect 5156 8600 5157 9320
rect 4435 8599 5157 8600
rect 4016 8532 4112 8548
rect 5428 8548 5444 9372
rect 5508 8548 5524 9372
rect 6840 9372 6936 9388
rect 5847 9320 6569 9321
rect 5847 8600 5848 9320
rect 6568 8600 6569 9320
rect 5847 8599 6569 8600
rect 5428 8532 5524 8548
rect 6840 8548 6856 9372
rect 6920 8548 6936 9372
rect 8252 9372 8348 9388
rect 7259 9320 7981 9321
rect 7259 8600 7260 9320
rect 7980 8600 7981 9320
rect 7259 8599 7981 8600
rect 6840 8532 6936 8548
rect 8252 8548 8268 9372
rect 8332 8548 8348 9372
rect 9664 9372 9760 9388
rect 8671 9320 9393 9321
rect 8671 8600 8672 9320
rect 9392 8600 9393 9320
rect 8671 8599 9393 8600
rect 8252 8532 8348 8548
rect 9664 8548 9680 9372
rect 9744 8548 9760 9372
rect 11076 9372 11172 9388
rect 10083 9320 10805 9321
rect 10083 8600 10084 9320
rect 10804 8600 10805 9320
rect 10083 8599 10805 8600
rect 9664 8532 9760 8548
rect 11076 8548 11092 9372
rect 11156 8548 11172 9372
rect 12488 9372 12584 9388
rect 11495 9320 12217 9321
rect 11495 8600 11496 9320
rect 12216 8600 12217 9320
rect 11495 8599 12217 8600
rect 11076 8532 11172 8548
rect 12488 8548 12504 9372
rect 12568 8548 12584 9372
rect 13900 9372 13996 9388
rect 12907 9320 13629 9321
rect 12907 8600 12908 9320
rect 13628 8600 13629 9320
rect 12907 8599 13629 8600
rect 12488 8532 12584 8548
rect 13900 8548 13916 9372
rect 13980 8548 13996 9372
rect 15312 9372 15408 9388
rect 14319 9320 15041 9321
rect 14319 8600 14320 9320
rect 15040 8600 15041 9320
rect 14319 8599 15041 8600
rect 13900 8532 13996 8548
rect 15312 8548 15328 9372
rect 15392 8548 15408 9372
rect 16724 9372 16820 9388
rect 15731 9320 16453 9321
rect 15731 8600 15732 9320
rect 16452 8600 16453 9320
rect 15731 8599 16453 8600
rect 15312 8532 15408 8548
rect 16724 8548 16740 9372
rect 16804 8548 16820 9372
rect 18136 9372 18232 9388
rect 17143 9320 17865 9321
rect 17143 8600 17144 9320
rect 17864 8600 17865 9320
rect 17143 8599 17865 8600
rect 16724 8532 16820 8548
rect 18136 8548 18152 9372
rect 18216 8548 18232 9372
rect 19548 9372 19644 9388
rect 18555 9320 19277 9321
rect 18555 8600 18556 9320
rect 19276 8600 19277 9320
rect 18555 8599 19277 8600
rect 18136 8532 18232 8548
rect 19548 8548 19564 9372
rect 19628 8548 19644 9372
rect 20960 9372 21056 9388
rect 19967 9320 20689 9321
rect 19967 8600 19968 9320
rect 20688 8600 20689 9320
rect 19967 8599 20689 8600
rect 19548 8532 19644 8548
rect 20960 8548 20976 9372
rect 21040 8548 21056 9372
rect 22372 9372 22468 9388
rect 21379 9320 22101 9321
rect 21379 8600 21380 9320
rect 22100 8600 22101 9320
rect 21379 8599 22101 8600
rect 20960 8532 21056 8548
rect 22372 8548 22388 9372
rect 22452 8548 22468 9372
rect 23784 9372 23880 9388
rect 22791 9320 23513 9321
rect 22791 8600 22792 9320
rect 23512 8600 23513 9320
rect 22791 8599 23513 8600
rect 22372 8532 22468 8548
rect 23784 8548 23800 9372
rect 23864 8548 23880 9372
rect 23784 8532 23880 8548
rect -22812 8252 -22716 8268
rect -23805 8200 -23083 8201
rect -23805 7480 -23804 8200
rect -23084 7480 -23083 8200
rect -23805 7479 -23083 7480
rect -22812 7428 -22796 8252
rect -22732 7428 -22716 8252
rect -21400 8252 -21304 8268
rect -22393 8200 -21671 8201
rect -22393 7480 -22392 8200
rect -21672 7480 -21671 8200
rect -22393 7479 -21671 7480
rect -22812 7412 -22716 7428
rect -21400 7428 -21384 8252
rect -21320 7428 -21304 8252
rect -19988 8252 -19892 8268
rect -20981 8200 -20259 8201
rect -20981 7480 -20980 8200
rect -20260 7480 -20259 8200
rect -20981 7479 -20259 7480
rect -21400 7412 -21304 7428
rect -19988 7428 -19972 8252
rect -19908 7428 -19892 8252
rect -18576 8252 -18480 8268
rect -19569 8200 -18847 8201
rect -19569 7480 -19568 8200
rect -18848 7480 -18847 8200
rect -19569 7479 -18847 7480
rect -19988 7412 -19892 7428
rect -18576 7428 -18560 8252
rect -18496 7428 -18480 8252
rect -17164 8252 -17068 8268
rect -18157 8200 -17435 8201
rect -18157 7480 -18156 8200
rect -17436 7480 -17435 8200
rect -18157 7479 -17435 7480
rect -18576 7412 -18480 7428
rect -17164 7428 -17148 8252
rect -17084 7428 -17068 8252
rect -15752 8252 -15656 8268
rect -16745 8200 -16023 8201
rect -16745 7480 -16744 8200
rect -16024 7480 -16023 8200
rect -16745 7479 -16023 7480
rect -17164 7412 -17068 7428
rect -15752 7428 -15736 8252
rect -15672 7428 -15656 8252
rect -14340 8252 -14244 8268
rect -15333 8200 -14611 8201
rect -15333 7480 -15332 8200
rect -14612 7480 -14611 8200
rect -15333 7479 -14611 7480
rect -15752 7412 -15656 7428
rect -14340 7428 -14324 8252
rect -14260 7428 -14244 8252
rect -12928 8252 -12832 8268
rect -13921 8200 -13199 8201
rect -13921 7480 -13920 8200
rect -13200 7480 -13199 8200
rect -13921 7479 -13199 7480
rect -14340 7412 -14244 7428
rect -12928 7428 -12912 8252
rect -12848 7428 -12832 8252
rect -11516 8252 -11420 8268
rect -12509 8200 -11787 8201
rect -12509 7480 -12508 8200
rect -11788 7480 -11787 8200
rect -12509 7479 -11787 7480
rect -12928 7412 -12832 7428
rect -11516 7428 -11500 8252
rect -11436 7428 -11420 8252
rect -10104 8252 -10008 8268
rect -11097 8200 -10375 8201
rect -11097 7480 -11096 8200
rect -10376 7480 -10375 8200
rect -11097 7479 -10375 7480
rect -11516 7412 -11420 7428
rect -10104 7428 -10088 8252
rect -10024 7428 -10008 8252
rect -8692 8252 -8596 8268
rect -9685 8200 -8963 8201
rect -9685 7480 -9684 8200
rect -8964 7480 -8963 8200
rect -9685 7479 -8963 7480
rect -10104 7412 -10008 7428
rect -8692 7428 -8676 8252
rect -8612 7428 -8596 8252
rect -7280 8252 -7184 8268
rect -8273 8200 -7551 8201
rect -8273 7480 -8272 8200
rect -7552 7480 -7551 8200
rect -8273 7479 -7551 7480
rect -8692 7412 -8596 7428
rect -7280 7428 -7264 8252
rect -7200 7428 -7184 8252
rect -5868 8252 -5772 8268
rect -6861 8200 -6139 8201
rect -6861 7480 -6860 8200
rect -6140 7480 -6139 8200
rect -6861 7479 -6139 7480
rect -7280 7412 -7184 7428
rect -5868 7428 -5852 8252
rect -5788 7428 -5772 8252
rect -4456 8252 -4360 8268
rect -5449 8200 -4727 8201
rect -5449 7480 -5448 8200
rect -4728 7480 -4727 8200
rect -5449 7479 -4727 7480
rect -5868 7412 -5772 7428
rect -4456 7428 -4440 8252
rect -4376 7428 -4360 8252
rect -3044 8252 -2948 8268
rect -4037 8200 -3315 8201
rect -4037 7480 -4036 8200
rect -3316 7480 -3315 8200
rect -4037 7479 -3315 7480
rect -4456 7412 -4360 7428
rect -3044 7428 -3028 8252
rect -2964 7428 -2948 8252
rect -1632 8252 -1536 8268
rect -2625 8200 -1903 8201
rect -2625 7480 -2624 8200
rect -1904 7480 -1903 8200
rect -2625 7479 -1903 7480
rect -3044 7412 -2948 7428
rect -1632 7428 -1616 8252
rect -1552 7428 -1536 8252
rect -220 8252 -124 8268
rect -1213 8200 -491 8201
rect -1213 7480 -1212 8200
rect -492 7480 -491 8200
rect -1213 7479 -491 7480
rect -1632 7412 -1536 7428
rect -220 7428 -204 8252
rect -140 7428 -124 8252
rect 1192 8252 1288 8268
rect 199 8200 921 8201
rect 199 7480 200 8200
rect 920 7480 921 8200
rect 199 7479 921 7480
rect -220 7412 -124 7428
rect 1192 7428 1208 8252
rect 1272 7428 1288 8252
rect 2604 8252 2700 8268
rect 1611 8200 2333 8201
rect 1611 7480 1612 8200
rect 2332 7480 2333 8200
rect 1611 7479 2333 7480
rect 1192 7412 1288 7428
rect 2604 7428 2620 8252
rect 2684 7428 2700 8252
rect 4016 8252 4112 8268
rect 3023 8200 3745 8201
rect 3023 7480 3024 8200
rect 3744 7480 3745 8200
rect 3023 7479 3745 7480
rect 2604 7412 2700 7428
rect 4016 7428 4032 8252
rect 4096 7428 4112 8252
rect 5428 8252 5524 8268
rect 4435 8200 5157 8201
rect 4435 7480 4436 8200
rect 5156 7480 5157 8200
rect 4435 7479 5157 7480
rect 4016 7412 4112 7428
rect 5428 7428 5444 8252
rect 5508 7428 5524 8252
rect 6840 8252 6936 8268
rect 5847 8200 6569 8201
rect 5847 7480 5848 8200
rect 6568 7480 6569 8200
rect 5847 7479 6569 7480
rect 5428 7412 5524 7428
rect 6840 7428 6856 8252
rect 6920 7428 6936 8252
rect 8252 8252 8348 8268
rect 7259 8200 7981 8201
rect 7259 7480 7260 8200
rect 7980 7480 7981 8200
rect 7259 7479 7981 7480
rect 6840 7412 6936 7428
rect 8252 7428 8268 8252
rect 8332 7428 8348 8252
rect 9664 8252 9760 8268
rect 8671 8200 9393 8201
rect 8671 7480 8672 8200
rect 9392 7480 9393 8200
rect 8671 7479 9393 7480
rect 8252 7412 8348 7428
rect 9664 7428 9680 8252
rect 9744 7428 9760 8252
rect 11076 8252 11172 8268
rect 10083 8200 10805 8201
rect 10083 7480 10084 8200
rect 10804 7480 10805 8200
rect 10083 7479 10805 7480
rect 9664 7412 9760 7428
rect 11076 7428 11092 8252
rect 11156 7428 11172 8252
rect 12488 8252 12584 8268
rect 11495 8200 12217 8201
rect 11495 7480 11496 8200
rect 12216 7480 12217 8200
rect 11495 7479 12217 7480
rect 11076 7412 11172 7428
rect 12488 7428 12504 8252
rect 12568 7428 12584 8252
rect 13900 8252 13996 8268
rect 12907 8200 13629 8201
rect 12907 7480 12908 8200
rect 13628 7480 13629 8200
rect 12907 7479 13629 7480
rect 12488 7412 12584 7428
rect 13900 7428 13916 8252
rect 13980 7428 13996 8252
rect 15312 8252 15408 8268
rect 14319 8200 15041 8201
rect 14319 7480 14320 8200
rect 15040 7480 15041 8200
rect 14319 7479 15041 7480
rect 13900 7412 13996 7428
rect 15312 7428 15328 8252
rect 15392 7428 15408 8252
rect 16724 8252 16820 8268
rect 15731 8200 16453 8201
rect 15731 7480 15732 8200
rect 16452 7480 16453 8200
rect 15731 7479 16453 7480
rect 15312 7412 15408 7428
rect 16724 7428 16740 8252
rect 16804 7428 16820 8252
rect 18136 8252 18232 8268
rect 17143 8200 17865 8201
rect 17143 7480 17144 8200
rect 17864 7480 17865 8200
rect 17143 7479 17865 7480
rect 16724 7412 16820 7428
rect 18136 7428 18152 8252
rect 18216 7428 18232 8252
rect 19548 8252 19644 8268
rect 18555 8200 19277 8201
rect 18555 7480 18556 8200
rect 19276 7480 19277 8200
rect 18555 7479 19277 7480
rect 18136 7412 18232 7428
rect 19548 7428 19564 8252
rect 19628 7428 19644 8252
rect 20960 8252 21056 8268
rect 19967 8200 20689 8201
rect 19967 7480 19968 8200
rect 20688 7480 20689 8200
rect 19967 7479 20689 7480
rect 19548 7412 19644 7428
rect 20960 7428 20976 8252
rect 21040 7428 21056 8252
rect 22372 8252 22468 8268
rect 21379 8200 22101 8201
rect 21379 7480 21380 8200
rect 22100 7480 22101 8200
rect 21379 7479 22101 7480
rect 20960 7412 21056 7428
rect 22372 7428 22388 8252
rect 22452 7428 22468 8252
rect 23784 8252 23880 8268
rect 22791 8200 23513 8201
rect 22791 7480 22792 8200
rect 23512 7480 23513 8200
rect 22791 7479 23513 7480
rect 22372 7412 22468 7428
rect 23784 7428 23800 8252
rect 23864 7428 23880 8252
rect 23784 7412 23880 7428
rect -22812 7132 -22716 7148
rect -23805 7080 -23083 7081
rect -23805 6360 -23804 7080
rect -23084 6360 -23083 7080
rect -23805 6359 -23083 6360
rect -22812 6308 -22796 7132
rect -22732 6308 -22716 7132
rect -21400 7132 -21304 7148
rect -22393 7080 -21671 7081
rect -22393 6360 -22392 7080
rect -21672 6360 -21671 7080
rect -22393 6359 -21671 6360
rect -22812 6292 -22716 6308
rect -21400 6308 -21384 7132
rect -21320 6308 -21304 7132
rect -19988 7132 -19892 7148
rect -20981 7080 -20259 7081
rect -20981 6360 -20980 7080
rect -20260 6360 -20259 7080
rect -20981 6359 -20259 6360
rect -21400 6292 -21304 6308
rect -19988 6308 -19972 7132
rect -19908 6308 -19892 7132
rect -18576 7132 -18480 7148
rect -19569 7080 -18847 7081
rect -19569 6360 -19568 7080
rect -18848 6360 -18847 7080
rect -19569 6359 -18847 6360
rect -19988 6292 -19892 6308
rect -18576 6308 -18560 7132
rect -18496 6308 -18480 7132
rect -17164 7132 -17068 7148
rect -18157 7080 -17435 7081
rect -18157 6360 -18156 7080
rect -17436 6360 -17435 7080
rect -18157 6359 -17435 6360
rect -18576 6292 -18480 6308
rect -17164 6308 -17148 7132
rect -17084 6308 -17068 7132
rect -15752 7132 -15656 7148
rect -16745 7080 -16023 7081
rect -16745 6360 -16744 7080
rect -16024 6360 -16023 7080
rect -16745 6359 -16023 6360
rect -17164 6292 -17068 6308
rect -15752 6308 -15736 7132
rect -15672 6308 -15656 7132
rect -14340 7132 -14244 7148
rect -15333 7080 -14611 7081
rect -15333 6360 -15332 7080
rect -14612 6360 -14611 7080
rect -15333 6359 -14611 6360
rect -15752 6292 -15656 6308
rect -14340 6308 -14324 7132
rect -14260 6308 -14244 7132
rect -12928 7132 -12832 7148
rect -13921 7080 -13199 7081
rect -13921 6360 -13920 7080
rect -13200 6360 -13199 7080
rect -13921 6359 -13199 6360
rect -14340 6292 -14244 6308
rect -12928 6308 -12912 7132
rect -12848 6308 -12832 7132
rect -11516 7132 -11420 7148
rect -12509 7080 -11787 7081
rect -12509 6360 -12508 7080
rect -11788 6360 -11787 7080
rect -12509 6359 -11787 6360
rect -12928 6292 -12832 6308
rect -11516 6308 -11500 7132
rect -11436 6308 -11420 7132
rect -10104 7132 -10008 7148
rect -11097 7080 -10375 7081
rect -11097 6360 -11096 7080
rect -10376 6360 -10375 7080
rect -11097 6359 -10375 6360
rect -11516 6292 -11420 6308
rect -10104 6308 -10088 7132
rect -10024 6308 -10008 7132
rect -8692 7132 -8596 7148
rect -9685 7080 -8963 7081
rect -9685 6360 -9684 7080
rect -8964 6360 -8963 7080
rect -9685 6359 -8963 6360
rect -10104 6292 -10008 6308
rect -8692 6308 -8676 7132
rect -8612 6308 -8596 7132
rect -7280 7132 -7184 7148
rect -8273 7080 -7551 7081
rect -8273 6360 -8272 7080
rect -7552 6360 -7551 7080
rect -8273 6359 -7551 6360
rect -8692 6292 -8596 6308
rect -7280 6308 -7264 7132
rect -7200 6308 -7184 7132
rect -5868 7132 -5772 7148
rect -6861 7080 -6139 7081
rect -6861 6360 -6860 7080
rect -6140 6360 -6139 7080
rect -6861 6359 -6139 6360
rect -7280 6292 -7184 6308
rect -5868 6308 -5852 7132
rect -5788 6308 -5772 7132
rect -4456 7132 -4360 7148
rect -5449 7080 -4727 7081
rect -5449 6360 -5448 7080
rect -4728 6360 -4727 7080
rect -5449 6359 -4727 6360
rect -5868 6292 -5772 6308
rect -4456 6308 -4440 7132
rect -4376 6308 -4360 7132
rect -3044 7132 -2948 7148
rect -4037 7080 -3315 7081
rect -4037 6360 -4036 7080
rect -3316 6360 -3315 7080
rect -4037 6359 -3315 6360
rect -4456 6292 -4360 6308
rect -3044 6308 -3028 7132
rect -2964 6308 -2948 7132
rect -1632 7132 -1536 7148
rect -2625 7080 -1903 7081
rect -2625 6360 -2624 7080
rect -1904 6360 -1903 7080
rect -2625 6359 -1903 6360
rect -3044 6292 -2948 6308
rect -1632 6308 -1616 7132
rect -1552 6308 -1536 7132
rect -220 7132 -124 7148
rect -1213 7080 -491 7081
rect -1213 6360 -1212 7080
rect -492 6360 -491 7080
rect -1213 6359 -491 6360
rect -1632 6292 -1536 6308
rect -220 6308 -204 7132
rect -140 6308 -124 7132
rect 1192 7132 1288 7148
rect 199 7080 921 7081
rect 199 6360 200 7080
rect 920 6360 921 7080
rect 199 6359 921 6360
rect -220 6292 -124 6308
rect 1192 6308 1208 7132
rect 1272 6308 1288 7132
rect 2604 7132 2700 7148
rect 1611 7080 2333 7081
rect 1611 6360 1612 7080
rect 2332 6360 2333 7080
rect 1611 6359 2333 6360
rect 1192 6292 1288 6308
rect 2604 6308 2620 7132
rect 2684 6308 2700 7132
rect 4016 7132 4112 7148
rect 3023 7080 3745 7081
rect 3023 6360 3024 7080
rect 3744 6360 3745 7080
rect 3023 6359 3745 6360
rect 2604 6292 2700 6308
rect 4016 6308 4032 7132
rect 4096 6308 4112 7132
rect 5428 7132 5524 7148
rect 4435 7080 5157 7081
rect 4435 6360 4436 7080
rect 5156 6360 5157 7080
rect 4435 6359 5157 6360
rect 4016 6292 4112 6308
rect 5428 6308 5444 7132
rect 5508 6308 5524 7132
rect 6840 7132 6936 7148
rect 5847 7080 6569 7081
rect 5847 6360 5848 7080
rect 6568 6360 6569 7080
rect 5847 6359 6569 6360
rect 5428 6292 5524 6308
rect 6840 6308 6856 7132
rect 6920 6308 6936 7132
rect 8252 7132 8348 7148
rect 7259 7080 7981 7081
rect 7259 6360 7260 7080
rect 7980 6360 7981 7080
rect 7259 6359 7981 6360
rect 6840 6292 6936 6308
rect 8252 6308 8268 7132
rect 8332 6308 8348 7132
rect 9664 7132 9760 7148
rect 8671 7080 9393 7081
rect 8671 6360 8672 7080
rect 9392 6360 9393 7080
rect 8671 6359 9393 6360
rect 8252 6292 8348 6308
rect 9664 6308 9680 7132
rect 9744 6308 9760 7132
rect 11076 7132 11172 7148
rect 10083 7080 10805 7081
rect 10083 6360 10084 7080
rect 10804 6360 10805 7080
rect 10083 6359 10805 6360
rect 9664 6292 9760 6308
rect 11076 6308 11092 7132
rect 11156 6308 11172 7132
rect 12488 7132 12584 7148
rect 11495 7080 12217 7081
rect 11495 6360 11496 7080
rect 12216 6360 12217 7080
rect 11495 6359 12217 6360
rect 11076 6292 11172 6308
rect 12488 6308 12504 7132
rect 12568 6308 12584 7132
rect 13900 7132 13996 7148
rect 12907 7080 13629 7081
rect 12907 6360 12908 7080
rect 13628 6360 13629 7080
rect 12907 6359 13629 6360
rect 12488 6292 12584 6308
rect 13900 6308 13916 7132
rect 13980 6308 13996 7132
rect 15312 7132 15408 7148
rect 14319 7080 15041 7081
rect 14319 6360 14320 7080
rect 15040 6360 15041 7080
rect 14319 6359 15041 6360
rect 13900 6292 13996 6308
rect 15312 6308 15328 7132
rect 15392 6308 15408 7132
rect 16724 7132 16820 7148
rect 15731 7080 16453 7081
rect 15731 6360 15732 7080
rect 16452 6360 16453 7080
rect 15731 6359 16453 6360
rect 15312 6292 15408 6308
rect 16724 6308 16740 7132
rect 16804 6308 16820 7132
rect 18136 7132 18232 7148
rect 17143 7080 17865 7081
rect 17143 6360 17144 7080
rect 17864 6360 17865 7080
rect 17143 6359 17865 6360
rect 16724 6292 16820 6308
rect 18136 6308 18152 7132
rect 18216 6308 18232 7132
rect 19548 7132 19644 7148
rect 18555 7080 19277 7081
rect 18555 6360 18556 7080
rect 19276 6360 19277 7080
rect 18555 6359 19277 6360
rect 18136 6292 18232 6308
rect 19548 6308 19564 7132
rect 19628 6308 19644 7132
rect 20960 7132 21056 7148
rect 19967 7080 20689 7081
rect 19967 6360 19968 7080
rect 20688 6360 20689 7080
rect 19967 6359 20689 6360
rect 19548 6292 19644 6308
rect 20960 6308 20976 7132
rect 21040 6308 21056 7132
rect 22372 7132 22468 7148
rect 21379 7080 22101 7081
rect 21379 6360 21380 7080
rect 22100 6360 22101 7080
rect 21379 6359 22101 6360
rect 20960 6292 21056 6308
rect 22372 6308 22388 7132
rect 22452 6308 22468 7132
rect 23784 7132 23880 7148
rect 22791 7080 23513 7081
rect 22791 6360 22792 7080
rect 23512 6360 23513 7080
rect 22791 6359 23513 6360
rect 22372 6292 22468 6308
rect 23784 6308 23800 7132
rect 23864 6308 23880 7132
rect 23784 6292 23880 6308
rect -22812 6012 -22716 6028
rect -23805 5960 -23083 5961
rect -23805 5240 -23804 5960
rect -23084 5240 -23083 5960
rect -23805 5239 -23083 5240
rect -22812 5188 -22796 6012
rect -22732 5188 -22716 6012
rect -21400 6012 -21304 6028
rect -22393 5960 -21671 5961
rect -22393 5240 -22392 5960
rect -21672 5240 -21671 5960
rect -22393 5239 -21671 5240
rect -22812 5172 -22716 5188
rect -21400 5188 -21384 6012
rect -21320 5188 -21304 6012
rect -19988 6012 -19892 6028
rect -20981 5960 -20259 5961
rect -20981 5240 -20980 5960
rect -20260 5240 -20259 5960
rect -20981 5239 -20259 5240
rect -21400 5172 -21304 5188
rect -19988 5188 -19972 6012
rect -19908 5188 -19892 6012
rect -18576 6012 -18480 6028
rect -19569 5960 -18847 5961
rect -19569 5240 -19568 5960
rect -18848 5240 -18847 5960
rect -19569 5239 -18847 5240
rect -19988 5172 -19892 5188
rect -18576 5188 -18560 6012
rect -18496 5188 -18480 6012
rect -17164 6012 -17068 6028
rect -18157 5960 -17435 5961
rect -18157 5240 -18156 5960
rect -17436 5240 -17435 5960
rect -18157 5239 -17435 5240
rect -18576 5172 -18480 5188
rect -17164 5188 -17148 6012
rect -17084 5188 -17068 6012
rect -15752 6012 -15656 6028
rect -16745 5960 -16023 5961
rect -16745 5240 -16744 5960
rect -16024 5240 -16023 5960
rect -16745 5239 -16023 5240
rect -17164 5172 -17068 5188
rect -15752 5188 -15736 6012
rect -15672 5188 -15656 6012
rect -14340 6012 -14244 6028
rect -15333 5960 -14611 5961
rect -15333 5240 -15332 5960
rect -14612 5240 -14611 5960
rect -15333 5239 -14611 5240
rect -15752 5172 -15656 5188
rect -14340 5188 -14324 6012
rect -14260 5188 -14244 6012
rect -12928 6012 -12832 6028
rect -13921 5960 -13199 5961
rect -13921 5240 -13920 5960
rect -13200 5240 -13199 5960
rect -13921 5239 -13199 5240
rect -14340 5172 -14244 5188
rect -12928 5188 -12912 6012
rect -12848 5188 -12832 6012
rect -11516 6012 -11420 6028
rect -12509 5960 -11787 5961
rect -12509 5240 -12508 5960
rect -11788 5240 -11787 5960
rect -12509 5239 -11787 5240
rect -12928 5172 -12832 5188
rect -11516 5188 -11500 6012
rect -11436 5188 -11420 6012
rect -10104 6012 -10008 6028
rect -11097 5960 -10375 5961
rect -11097 5240 -11096 5960
rect -10376 5240 -10375 5960
rect -11097 5239 -10375 5240
rect -11516 5172 -11420 5188
rect -10104 5188 -10088 6012
rect -10024 5188 -10008 6012
rect -8692 6012 -8596 6028
rect -9685 5960 -8963 5961
rect -9685 5240 -9684 5960
rect -8964 5240 -8963 5960
rect -9685 5239 -8963 5240
rect -10104 5172 -10008 5188
rect -8692 5188 -8676 6012
rect -8612 5188 -8596 6012
rect -7280 6012 -7184 6028
rect -8273 5960 -7551 5961
rect -8273 5240 -8272 5960
rect -7552 5240 -7551 5960
rect -8273 5239 -7551 5240
rect -8692 5172 -8596 5188
rect -7280 5188 -7264 6012
rect -7200 5188 -7184 6012
rect -5868 6012 -5772 6028
rect -6861 5960 -6139 5961
rect -6861 5240 -6860 5960
rect -6140 5240 -6139 5960
rect -6861 5239 -6139 5240
rect -7280 5172 -7184 5188
rect -5868 5188 -5852 6012
rect -5788 5188 -5772 6012
rect -4456 6012 -4360 6028
rect -5449 5960 -4727 5961
rect -5449 5240 -5448 5960
rect -4728 5240 -4727 5960
rect -5449 5239 -4727 5240
rect -5868 5172 -5772 5188
rect -4456 5188 -4440 6012
rect -4376 5188 -4360 6012
rect -3044 6012 -2948 6028
rect -4037 5960 -3315 5961
rect -4037 5240 -4036 5960
rect -3316 5240 -3315 5960
rect -4037 5239 -3315 5240
rect -4456 5172 -4360 5188
rect -3044 5188 -3028 6012
rect -2964 5188 -2948 6012
rect -1632 6012 -1536 6028
rect -2625 5960 -1903 5961
rect -2625 5240 -2624 5960
rect -1904 5240 -1903 5960
rect -2625 5239 -1903 5240
rect -3044 5172 -2948 5188
rect -1632 5188 -1616 6012
rect -1552 5188 -1536 6012
rect -220 6012 -124 6028
rect -1213 5960 -491 5961
rect -1213 5240 -1212 5960
rect -492 5240 -491 5960
rect -1213 5239 -491 5240
rect -1632 5172 -1536 5188
rect -220 5188 -204 6012
rect -140 5188 -124 6012
rect 1192 6012 1288 6028
rect 199 5960 921 5961
rect 199 5240 200 5960
rect 920 5240 921 5960
rect 199 5239 921 5240
rect -220 5172 -124 5188
rect 1192 5188 1208 6012
rect 1272 5188 1288 6012
rect 2604 6012 2700 6028
rect 1611 5960 2333 5961
rect 1611 5240 1612 5960
rect 2332 5240 2333 5960
rect 1611 5239 2333 5240
rect 1192 5172 1288 5188
rect 2604 5188 2620 6012
rect 2684 5188 2700 6012
rect 4016 6012 4112 6028
rect 3023 5960 3745 5961
rect 3023 5240 3024 5960
rect 3744 5240 3745 5960
rect 3023 5239 3745 5240
rect 2604 5172 2700 5188
rect 4016 5188 4032 6012
rect 4096 5188 4112 6012
rect 5428 6012 5524 6028
rect 4435 5960 5157 5961
rect 4435 5240 4436 5960
rect 5156 5240 5157 5960
rect 4435 5239 5157 5240
rect 4016 5172 4112 5188
rect 5428 5188 5444 6012
rect 5508 5188 5524 6012
rect 6840 6012 6936 6028
rect 5847 5960 6569 5961
rect 5847 5240 5848 5960
rect 6568 5240 6569 5960
rect 5847 5239 6569 5240
rect 5428 5172 5524 5188
rect 6840 5188 6856 6012
rect 6920 5188 6936 6012
rect 8252 6012 8348 6028
rect 7259 5960 7981 5961
rect 7259 5240 7260 5960
rect 7980 5240 7981 5960
rect 7259 5239 7981 5240
rect 6840 5172 6936 5188
rect 8252 5188 8268 6012
rect 8332 5188 8348 6012
rect 9664 6012 9760 6028
rect 8671 5960 9393 5961
rect 8671 5240 8672 5960
rect 9392 5240 9393 5960
rect 8671 5239 9393 5240
rect 8252 5172 8348 5188
rect 9664 5188 9680 6012
rect 9744 5188 9760 6012
rect 11076 6012 11172 6028
rect 10083 5960 10805 5961
rect 10083 5240 10084 5960
rect 10804 5240 10805 5960
rect 10083 5239 10805 5240
rect 9664 5172 9760 5188
rect 11076 5188 11092 6012
rect 11156 5188 11172 6012
rect 12488 6012 12584 6028
rect 11495 5960 12217 5961
rect 11495 5240 11496 5960
rect 12216 5240 12217 5960
rect 11495 5239 12217 5240
rect 11076 5172 11172 5188
rect 12488 5188 12504 6012
rect 12568 5188 12584 6012
rect 13900 6012 13996 6028
rect 12907 5960 13629 5961
rect 12907 5240 12908 5960
rect 13628 5240 13629 5960
rect 12907 5239 13629 5240
rect 12488 5172 12584 5188
rect 13900 5188 13916 6012
rect 13980 5188 13996 6012
rect 15312 6012 15408 6028
rect 14319 5960 15041 5961
rect 14319 5240 14320 5960
rect 15040 5240 15041 5960
rect 14319 5239 15041 5240
rect 13900 5172 13996 5188
rect 15312 5188 15328 6012
rect 15392 5188 15408 6012
rect 16724 6012 16820 6028
rect 15731 5960 16453 5961
rect 15731 5240 15732 5960
rect 16452 5240 16453 5960
rect 15731 5239 16453 5240
rect 15312 5172 15408 5188
rect 16724 5188 16740 6012
rect 16804 5188 16820 6012
rect 18136 6012 18232 6028
rect 17143 5960 17865 5961
rect 17143 5240 17144 5960
rect 17864 5240 17865 5960
rect 17143 5239 17865 5240
rect 16724 5172 16820 5188
rect 18136 5188 18152 6012
rect 18216 5188 18232 6012
rect 19548 6012 19644 6028
rect 18555 5960 19277 5961
rect 18555 5240 18556 5960
rect 19276 5240 19277 5960
rect 18555 5239 19277 5240
rect 18136 5172 18232 5188
rect 19548 5188 19564 6012
rect 19628 5188 19644 6012
rect 20960 6012 21056 6028
rect 19967 5960 20689 5961
rect 19967 5240 19968 5960
rect 20688 5240 20689 5960
rect 19967 5239 20689 5240
rect 19548 5172 19644 5188
rect 20960 5188 20976 6012
rect 21040 5188 21056 6012
rect 22372 6012 22468 6028
rect 21379 5960 22101 5961
rect 21379 5240 21380 5960
rect 22100 5240 22101 5960
rect 21379 5239 22101 5240
rect 20960 5172 21056 5188
rect 22372 5188 22388 6012
rect 22452 5188 22468 6012
rect 23784 6012 23880 6028
rect 22791 5960 23513 5961
rect 22791 5240 22792 5960
rect 23512 5240 23513 5960
rect 22791 5239 23513 5240
rect 22372 5172 22468 5188
rect 23784 5188 23800 6012
rect 23864 5188 23880 6012
rect 23784 5172 23880 5188
rect -22812 4892 -22716 4908
rect -23805 4840 -23083 4841
rect -23805 4120 -23804 4840
rect -23084 4120 -23083 4840
rect -23805 4119 -23083 4120
rect -22812 4068 -22796 4892
rect -22732 4068 -22716 4892
rect -21400 4892 -21304 4908
rect -22393 4840 -21671 4841
rect -22393 4120 -22392 4840
rect -21672 4120 -21671 4840
rect -22393 4119 -21671 4120
rect -22812 4052 -22716 4068
rect -21400 4068 -21384 4892
rect -21320 4068 -21304 4892
rect -19988 4892 -19892 4908
rect -20981 4840 -20259 4841
rect -20981 4120 -20980 4840
rect -20260 4120 -20259 4840
rect -20981 4119 -20259 4120
rect -21400 4052 -21304 4068
rect -19988 4068 -19972 4892
rect -19908 4068 -19892 4892
rect -18576 4892 -18480 4908
rect -19569 4840 -18847 4841
rect -19569 4120 -19568 4840
rect -18848 4120 -18847 4840
rect -19569 4119 -18847 4120
rect -19988 4052 -19892 4068
rect -18576 4068 -18560 4892
rect -18496 4068 -18480 4892
rect -17164 4892 -17068 4908
rect -18157 4840 -17435 4841
rect -18157 4120 -18156 4840
rect -17436 4120 -17435 4840
rect -18157 4119 -17435 4120
rect -18576 4052 -18480 4068
rect -17164 4068 -17148 4892
rect -17084 4068 -17068 4892
rect -15752 4892 -15656 4908
rect -16745 4840 -16023 4841
rect -16745 4120 -16744 4840
rect -16024 4120 -16023 4840
rect -16745 4119 -16023 4120
rect -17164 4052 -17068 4068
rect -15752 4068 -15736 4892
rect -15672 4068 -15656 4892
rect -14340 4892 -14244 4908
rect -15333 4840 -14611 4841
rect -15333 4120 -15332 4840
rect -14612 4120 -14611 4840
rect -15333 4119 -14611 4120
rect -15752 4052 -15656 4068
rect -14340 4068 -14324 4892
rect -14260 4068 -14244 4892
rect -12928 4892 -12832 4908
rect -13921 4840 -13199 4841
rect -13921 4120 -13920 4840
rect -13200 4120 -13199 4840
rect -13921 4119 -13199 4120
rect -14340 4052 -14244 4068
rect -12928 4068 -12912 4892
rect -12848 4068 -12832 4892
rect -11516 4892 -11420 4908
rect -12509 4840 -11787 4841
rect -12509 4120 -12508 4840
rect -11788 4120 -11787 4840
rect -12509 4119 -11787 4120
rect -12928 4052 -12832 4068
rect -11516 4068 -11500 4892
rect -11436 4068 -11420 4892
rect -10104 4892 -10008 4908
rect -11097 4840 -10375 4841
rect -11097 4120 -11096 4840
rect -10376 4120 -10375 4840
rect -11097 4119 -10375 4120
rect -11516 4052 -11420 4068
rect -10104 4068 -10088 4892
rect -10024 4068 -10008 4892
rect -8692 4892 -8596 4908
rect -9685 4840 -8963 4841
rect -9685 4120 -9684 4840
rect -8964 4120 -8963 4840
rect -9685 4119 -8963 4120
rect -10104 4052 -10008 4068
rect -8692 4068 -8676 4892
rect -8612 4068 -8596 4892
rect -7280 4892 -7184 4908
rect -8273 4840 -7551 4841
rect -8273 4120 -8272 4840
rect -7552 4120 -7551 4840
rect -8273 4119 -7551 4120
rect -8692 4052 -8596 4068
rect -7280 4068 -7264 4892
rect -7200 4068 -7184 4892
rect -5868 4892 -5772 4908
rect -6861 4840 -6139 4841
rect -6861 4120 -6860 4840
rect -6140 4120 -6139 4840
rect -6861 4119 -6139 4120
rect -7280 4052 -7184 4068
rect -5868 4068 -5852 4892
rect -5788 4068 -5772 4892
rect -4456 4892 -4360 4908
rect -5449 4840 -4727 4841
rect -5449 4120 -5448 4840
rect -4728 4120 -4727 4840
rect -5449 4119 -4727 4120
rect -5868 4052 -5772 4068
rect -4456 4068 -4440 4892
rect -4376 4068 -4360 4892
rect -3044 4892 -2948 4908
rect -4037 4840 -3315 4841
rect -4037 4120 -4036 4840
rect -3316 4120 -3315 4840
rect -4037 4119 -3315 4120
rect -4456 4052 -4360 4068
rect -3044 4068 -3028 4892
rect -2964 4068 -2948 4892
rect -1632 4892 -1536 4908
rect -2625 4840 -1903 4841
rect -2625 4120 -2624 4840
rect -1904 4120 -1903 4840
rect -2625 4119 -1903 4120
rect -3044 4052 -2948 4068
rect -1632 4068 -1616 4892
rect -1552 4068 -1536 4892
rect -220 4892 -124 4908
rect -1213 4840 -491 4841
rect -1213 4120 -1212 4840
rect -492 4120 -491 4840
rect -1213 4119 -491 4120
rect -1632 4052 -1536 4068
rect -220 4068 -204 4892
rect -140 4068 -124 4892
rect 1192 4892 1288 4908
rect 199 4840 921 4841
rect 199 4120 200 4840
rect 920 4120 921 4840
rect 199 4119 921 4120
rect -220 4052 -124 4068
rect 1192 4068 1208 4892
rect 1272 4068 1288 4892
rect 2604 4892 2700 4908
rect 1611 4840 2333 4841
rect 1611 4120 1612 4840
rect 2332 4120 2333 4840
rect 1611 4119 2333 4120
rect 1192 4052 1288 4068
rect 2604 4068 2620 4892
rect 2684 4068 2700 4892
rect 4016 4892 4112 4908
rect 3023 4840 3745 4841
rect 3023 4120 3024 4840
rect 3744 4120 3745 4840
rect 3023 4119 3745 4120
rect 2604 4052 2700 4068
rect 4016 4068 4032 4892
rect 4096 4068 4112 4892
rect 5428 4892 5524 4908
rect 4435 4840 5157 4841
rect 4435 4120 4436 4840
rect 5156 4120 5157 4840
rect 4435 4119 5157 4120
rect 4016 4052 4112 4068
rect 5428 4068 5444 4892
rect 5508 4068 5524 4892
rect 6840 4892 6936 4908
rect 5847 4840 6569 4841
rect 5847 4120 5848 4840
rect 6568 4120 6569 4840
rect 5847 4119 6569 4120
rect 5428 4052 5524 4068
rect 6840 4068 6856 4892
rect 6920 4068 6936 4892
rect 8252 4892 8348 4908
rect 7259 4840 7981 4841
rect 7259 4120 7260 4840
rect 7980 4120 7981 4840
rect 7259 4119 7981 4120
rect 6840 4052 6936 4068
rect 8252 4068 8268 4892
rect 8332 4068 8348 4892
rect 9664 4892 9760 4908
rect 8671 4840 9393 4841
rect 8671 4120 8672 4840
rect 9392 4120 9393 4840
rect 8671 4119 9393 4120
rect 8252 4052 8348 4068
rect 9664 4068 9680 4892
rect 9744 4068 9760 4892
rect 11076 4892 11172 4908
rect 10083 4840 10805 4841
rect 10083 4120 10084 4840
rect 10804 4120 10805 4840
rect 10083 4119 10805 4120
rect 9664 4052 9760 4068
rect 11076 4068 11092 4892
rect 11156 4068 11172 4892
rect 12488 4892 12584 4908
rect 11495 4840 12217 4841
rect 11495 4120 11496 4840
rect 12216 4120 12217 4840
rect 11495 4119 12217 4120
rect 11076 4052 11172 4068
rect 12488 4068 12504 4892
rect 12568 4068 12584 4892
rect 13900 4892 13996 4908
rect 12907 4840 13629 4841
rect 12907 4120 12908 4840
rect 13628 4120 13629 4840
rect 12907 4119 13629 4120
rect 12488 4052 12584 4068
rect 13900 4068 13916 4892
rect 13980 4068 13996 4892
rect 15312 4892 15408 4908
rect 14319 4840 15041 4841
rect 14319 4120 14320 4840
rect 15040 4120 15041 4840
rect 14319 4119 15041 4120
rect 13900 4052 13996 4068
rect 15312 4068 15328 4892
rect 15392 4068 15408 4892
rect 16724 4892 16820 4908
rect 15731 4840 16453 4841
rect 15731 4120 15732 4840
rect 16452 4120 16453 4840
rect 15731 4119 16453 4120
rect 15312 4052 15408 4068
rect 16724 4068 16740 4892
rect 16804 4068 16820 4892
rect 18136 4892 18232 4908
rect 17143 4840 17865 4841
rect 17143 4120 17144 4840
rect 17864 4120 17865 4840
rect 17143 4119 17865 4120
rect 16724 4052 16820 4068
rect 18136 4068 18152 4892
rect 18216 4068 18232 4892
rect 19548 4892 19644 4908
rect 18555 4840 19277 4841
rect 18555 4120 18556 4840
rect 19276 4120 19277 4840
rect 18555 4119 19277 4120
rect 18136 4052 18232 4068
rect 19548 4068 19564 4892
rect 19628 4068 19644 4892
rect 20960 4892 21056 4908
rect 19967 4840 20689 4841
rect 19967 4120 19968 4840
rect 20688 4120 20689 4840
rect 19967 4119 20689 4120
rect 19548 4052 19644 4068
rect 20960 4068 20976 4892
rect 21040 4068 21056 4892
rect 22372 4892 22468 4908
rect 21379 4840 22101 4841
rect 21379 4120 21380 4840
rect 22100 4120 22101 4840
rect 21379 4119 22101 4120
rect 20960 4052 21056 4068
rect 22372 4068 22388 4892
rect 22452 4068 22468 4892
rect 23784 4892 23880 4908
rect 22791 4840 23513 4841
rect 22791 4120 22792 4840
rect 23512 4120 23513 4840
rect 22791 4119 23513 4120
rect 22372 4052 22468 4068
rect 23784 4068 23800 4892
rect 23864 4068 23880 4892
rect 23784 4052 23880 4068
rect -22812 3772 -22716 3788
rect -23805 3720 -23083 3721
rect -23805 3000 -23804 3720
rect -23084 3000 -23083 3720
rect -23805 2999 -23083 3000
rect -22812 2948 -22796 3772
rect -22732 2948 -22716 3772
rect -21400 3772 -21304 3788
rect -22393 3720 -21671 3721
rect -22393 3000 -22392 3720
rect -21672 3000 -21671 3720
rect -22393 2999 -21671 3000
rect -22812 2932 -22716 2948
rect -21400 2948 -21384 3772
rect -21320 2948 -21304 3772
rect -19988 3772 -19892 3788
rect -20981 3720 -20259 3721
rect -20981 3000 -20980 3720
rect -20260 3000 -20259 3720
rect -20981 2999 -20259 3000
rect -21400 2932 -21304 2948
rect -19988 2948 -19972 3772
rect -19908 2948 -19892 3772
rect -18576 3772 -18480 3788
rect -19569 3720 -18847 3721
rect -19569 3000 -19568 3720
rect -18848 3000 -18847 3720
rect -19569 2999 -18847 3000
rect -19988 2932 -19892 2948
rect -18576 2948 -18560 3772
rect -18496 2948 -18480 3772
rect -17164 3772 -17068 3788
rect -18157 3720 -17435 3721
rect -18157 3000 -18156 3720
rect -17436 3000 -17435 3720
rect -18157 2999 -17435 3000
rect -18576 2932 -18480 2948
rect -17164 2948 -17148 3772
rect -17084 2948 -17068 3772
rect -15752 3772 -15656 3788
rect -16745 3720 -16023 3721
rect -16745 3000 -16744 3720
rect -16024 3000 -16023 3720
rect -16745 2999 -16023 3000
rect -17164 2932 -17068 2948
rect -15752 2948 -15736 3772
rect -15672 2948 -15656 3772
rect -14340 3772 -14244 3788
rect -15333 3720 -14611 3721
rect -15333 3000 -15332 3720
rect -14612 3000 -14611 3720
rect -15333 2999 -14611 3000
rect -15752 2932 -15656 2948
rect -14340 2948 -14324 3772
rect -14260 2948 -14244 3772
rect -12928 3772 -12832 3788
rect -13921 3720 -13199 3721
rect -13921 3000 -13920 3720
rect -13200 3000 -13199 3720
rect -13921 2999 -13199 3000
rect -14340 2932 -14244 2948
rect -12928 2948 -12912 3772
rect -12848 2948 -12832 3772
rect -11516 3772 -11420 3788
rect -12509 3720 -11787 3721
rect -12509 3000 -12508 3720
rect -11788 3000 -11787 3720
rect -12509 2999 -11787 3000
rect -12928 2932 -12832 2948
rect -11516 2948 -11500 3772
rect -11436 2948 -11420 3772
rect -10104 3772 -10008 3788
rect -11097 3720 -10375 3721
rect -11097 3000 -11096 3720
rect -10376 3000 -10375 3720
rect -11097 2999 -10375 3000
rect -11516 2932 -11420 2948
rect -10104 2948 -10088 3772
rect -10024 2948 -10008 3772
rect -8692 3772 -8596 3788
rect -9685 3720 -8963 3721
rect -9685 3000 -9684 3720
rect -8964 3000 -8963 3720
rect -9685 2999 -8963 3000
rect -10104 2932 -10008 2948
rect -8692 2948 -8676 3772
rect -8612 2948 -8596 3772
rect -7280 3772 -7184 3788
rect -8273 3720 -7551 3721
rect -8273 3000 -8272 3720
rect -7552 3000 -7551 3720
rect -8273 2999 -7551 3000
rect -8692 2932 -8596 2948
rect -7280 2948 -7264 3772
rect -7200 2948 -7184 3772
rect -5868 3772 -5772 3788
rect -6861 3720 -6139 3721
rect -6861 3000 -6860 3720
rect -6140 3000 -6139 3720
rect -6861 2999 -6139 3000
rect -7280 2932 -7184 2948
rect -5868 2948 -5852 3772
rect -5788 2948 -5772 3772
rect -4456 3772 -4360 3788
rect -5449 3720 -4727 3721
rect -5449 3000 -5448 3720
rect -4728 3000 -4727 3720
rect -5449 2999 -4727 3000
rect -5868 2932 -5772 2948
rect -4456 2948 -4440 3772
rect -4376 2948 -4360 3772
rect -3044 3772 -2948 3788
rect -4037 3720 -3315 3721
rect -4037 3000 -4036 3720
rect -3316 3000 -3315 3720
rect -4037 2999 -3315 3000
rect -4456 2932 -4360 2948
rect -3044 2948 -3028 3772
rect -2964 2948 -2948 3772
rect -1632 3772 -1536 3788
rect -2625 3720 -1903 3721
rect -2625 3000 -2624 3720
rect -1904 3000 -1903 3720
rect -2625 2999 -1903 3000
rect -3044 2932 -2948 2948
rect -1632 2948 -1616 3772
rect -1552 2948 -1536 3772
rect -220 3772 -124 3788
rect -1213 3720 -491 3721
rect -1213 3000 -1212 3720
rect -492 3000 -491 3720
rect -1213 2999 -491 3000
rect -1632 2932 -1536 2948
rect -220 2948 -204 3772
rect -140 2948 -124 3772
rect 1192 3772 1288 3788
rect 199 3720 921 3721
rect 199 3000 200 3720
rect 920 3000 921 3720
rect 199 2999 921 3000
rect -220 2932 -124 2948
rect 1192 2948 1208 3772
rect 1272 2948 1288 3772
rect 2604 3772 2700 3788
rect 1611 3720 2333 3721
rect 1611 3000 1612 3720
rect 2332 3000 2333 3720
rect 1611 2999 2333 3000
rect 1192 2932 1288 2948
rect 2604 2948 2620 3772
rect 2684 2948 2700 3772
rect 4016 3772 4112 3788
rect 3023 3720 3745 3721
rect 3023 3000 3024 3720
rect 3744 3000 3745 3720
rect 3023 2999 3745 3000
rect 2604 2932 2700 2948
rect 4016 2948 4032 3772
rect 4096 2948 4112 3772
rect 5428 3772 5524 3788
rect 4435 3720 5157 3721
rect 4435 3000 4436 3720
rect 5156 3000 5157 3720
rect 4435 2999 5157 3000
rect 4016 2932 4112 2948
rect 5428 2948 5444 3772
rect 5508 2948 5524 3772
rect 6840 3772 6936 3788
rect 5847 3720 6569 3721
rect 5847 3000 5848 3720
rect 6568 3000 6569 3720
rect 5847 2999 6569 3000
rect 5428 2932 5524 2948
rect 6840 2948 6856 3772
rect 6920 2948 6936 3772
rect 8252 3772 8348 3788
rect 7259 3720 7981 3721
rect 7259 3000 7260 3720
rect 7980 3000 7981 3720
rect 7259 2999 7981 3000
rect 6840 2932 6936 2948
rect 8252 2948 8268 3772
rect 8332 2948 8348 3772
rect 9664 3772 9760 3788
rect 8671 3720 9393 3721
rect 8671 3000 8672 3720
rect 9392 3000 9393 3720
rect 8671 2999 9393 3000
rect 8252 2932 8348 2948
rect 9664 2948 9680 3772
rect 9744 2948 9760 3772
rect 11076 3772 11172 3788
rect 10083 3720 10805 3721
rect 10083 3000 10084 3720
rect 10804 3000 10805 3720
rect 10083 2999 10805 3000
rect 9664 2932 9760 2948
rect 11076 2948 11092 3772
rect 11156 2948 11172 3772
rect 12488 3772 12584 3788
rect 11495 3720 12217 3721
rect 11495 3000 11496 3720
rect 12216 3000 12217 3720
rect 11495 2999 12217 3000
rect 11076 2932 11172 2948
rect 12488 2948 12504 3772
rect 12568 2948 12584 3772
rect 13900 3772 13996 3788
rect 12907 3720 13629 3721
rect 12907 3000 12908 3720
rect 13628 3000 13629 3720
rect 12907 2999 13629 3000
rect 12488 2932 12584 2948
rect 13900 2948 13916 3772
rect 13980 2948 13996 3772
rect 15312 3772 15408 3788
rect 14319 3720 15041 3721
rect 14319 3000 14320 3720
rect 15040 3000 15041 3720
rect 14319 2999 15041 3000
rect 13900 2932 13996 2948
rect 15312 2948 15328 3772
rect 15392 2948 15408 3772
rect 16724 3772 16820 3788
rect 15731 3720 16453 3721
rect 15731 3000 15732 3720
rect 16452 3000 16453 3720
rect 15731 2999 16453 3000
rect 15312 2932 15408 2948
rect 16724 2948 16740 3772
rect 16804 2948 16820 3772
rect 18136 3772 18232 3788
rect 17143 3720 17865 3721
rect 17143 3000 17144 3720
rect 17864 3000 17865 3720
rect 17143 2999 17865 3000
rect 16724 2932 16820 2948
rect 18136 2948 18152 3772
rect 18216 2948 18232 3772
rect 19548 3772 19644 3788
rect 18555 3720 19277 3721
rect 18555 3000 18556 3720
rect 19276 3000 19277 3720
rect 18555 2999 19277 3000
rect 18136 2932 18232 2948
rect 19548 2948 19564 3772
rect 19628 2948 19644 3772
rect 20960 3772 21056 3788
rect 19967 3720 20689 3721
rect 19967 3000 19968 3720
rect 20688 3000 20689 3720
rect 19967 2999 20689 3000
rect 19548 2932 19644 2948
rect 20960 2948 20976 3772
rect 21040 2948 21056 3772
rect 22372 3772 22468 3788
rect 21379 3720 22101 3721
rect 21379 3000 21380 3720
rect 22100 3000 22101 3720
rect 21379 2999 22101 3000
rect 20960 2932 21056 2948
rect 22372 2948 22388 3772
rect 22452 2948 22468 3772
rect 23784 3772 23880 3788
rect 22791 3720 23513 3721
rect 22791 3000 22792 3720
rect 23512 3000 23513 3720
rect 22791 2999 23513 3000
rect 22372 2932 22468 2948
rect 23784 2948 23800 3772
rect 23864 2948 23880 3772
rect 23784 2932 23880 2948
rect -22812 2652 -22716 2668
rect -23805 2600 -23083 2601
rect -23805 1880 -23804 2600
rect -23084 1880 -23083 2600
rect -23805 1879 -23083 1880
rect -22812 1828 -22796 2652
rect -22732 1828 -22716 2652
rect -21400 2652 -21304 2668
rect -22393 2600 -21671 2601
rect -22393 1880 -22392 2600
rect -21672 1880 -21671 2600
rect -22393 1879 -21671 1880
rect -22812 1812 -22716 1828
rect -21400 1828 -21384 2652
rect -21320 1828 -21304 2652
rect -19988 2652 -19892 2668
rect -20981 2600 -20259 2601
rect -20981 1880 -20980 2600
rect -20260 1880 -20259 2600
rect -20981 1879 -20259 1880
rect -21400 1812 -21304 1828
rect -19988 1828 -19972 2652
rect -19908 1828 -19892 2652
rect -18576 2652 -18480 2668
rect -19569 2600 -18847 2601
rect -19569 1880 -19568 2600
rect -18848 1880 -18847 2600
rect -19569 1879 -18847 1880
rect -19988 1812 -19892 1828
rect -18576 1828 -18560 2652
rect -18496 1828 -18480 2652
rect -17164 2652 -17068 2668
rect -18157 2600 -17435 2601
rect -18157 1880 -18156 2600
rect -17436 1880 -17435 2600
rect -18157 1879 -17435 1880
rect -18576 1812 -18480 1828
rect -17164 1828 -17148 2652
rect -17084 1828 -17068 2652
rect -15752 2652 -15656 2668
rect -16745 2600 -16023 2601
rect -16745 1880 -16744 2600
rect -16024 1880 -16023 2600
rect -16745 1879 -16023 1880
rect -17164 1812 -17068 1828
rect -15752 1828 -15736 2652
rect -15672 1828 -15656 2652
rect -14340 2652 -14244 2668
rect -15333 2600 -14611 2601
rect -15333 1880 -15332 2600
rect -14612 1880 -14611 2600
rect -15333 1879 -14611 1880
rect -15752 1812 -15656 1828
rect -14340 1828 -14324 2652
rect -14260 1828 -14244 2652
rect -12928 2652 -12832 2668
rect -13921 2600 -13199 2601
rect -13921 1880 -13920 2600
rect -13200 1880 -13199 2600
rect -13921 1879 -13199 1880
rect -14340 1812 -14244 1828
rect -12928 1828 -12912 2652
rect -12848 1828 -12832 2652
rect -11516 2652 -11420 2668
rect -12509 2600 -11787 2601
rect -12509 1880 -12508 2600
rect -11788 1880 -11787 2600
rect -12509 1879 -11787 1880
rect -12928 1812 -12832 1828
rect -11516 1828 -11500 2652
rect -11436 1828 -11420 2652
rect -10104 2652 -10008 2668
rect -11097 2600 -10375 2601
rect -11097 1880 -11096 2600
rect -10376 1880 -10375 2600
rect -11097 1879 -10375 1880
rect -11516 1812 -11420 1828
rect -10104 1828 -10088 2652
rect -10024 1828 -10008 2652
rect -8692 2652 -8596 2668
rect -9685 2600 -8963 2601
rect -9685 1880 -9684 2600
rect -8964 1880 -8963 2600
rect -9685 1879 -8963 1880
rect -10104 1812 -10008 1828
rect -8692 1828 -8676 2652
rect -8612 1828 -8596 2652
rect -7280 2652 -7184 2668
rect -8273 2600 -7551 2601
rect -8273 1880 -8272 2600
rect -7552 1880 -7551 2600
rect -8273 1879 -7551 1880
rect -8692 1812 -8596 1828
rect -7280 1828 -7264 2652
rect -7200 1828 -7184 2652
rect -5868 2652 -5772 2668
rect -6861 2600 -6139 2601
rect -6861 1880 -6860 2600
rect -6140 1880 -6139 2600
rect -6861 1879 -6139 1880
rect -7280 1812 -7184 1828
rect -5868 1828 -5852 2652
rect -5788 1828 -5772 2652
rect -4456 2652 -4360 2668
rect -5449 2600 -4727 2601
rect -5449 1880 -5448 2600
rect -4728 1880 -4727 2600
rect -5449 1879 -4727 1880
rect -5868 1812 -5772 1828
rect -4456 1828 -4440 2652
rect -4376 1828 -4360 2652
rect -3044 2652 -2948 2668
rect -4037 2600 -3315 2601
rect -4037 1880 -4036 2600
rect -3316 1880 -3315 2600
rect -4037 1879 -3315 1880
rect -4456 1812 -4360 1828
rect -3044 1828 -3028 2652
rect -2964 1828 -2948 2652
rect -1632 2652 -1536 2668
rect -2625 2600 -1903 2601
rect -2625 1880 -2624 2600
rect -1904 1880 -1903 2600
rect -2625 1879 -1903 1880
rect -3044 1812 -2948 1828
rect -1632 1828 -1616 2652
rect -1552 1828 -1536 2652
rect -220 2652 -124 2668
rect -1213 2600 -491 2601
rect -1213 1880 -1212 2600
rect -492 1880 -491 2600
rect -1213 1879 -491 1880
rect -1632 1812 -1536 1828
rect -220 1828 -204 2652
rect -140 1828 -124 2652
rect 1192 2652 1288 2668
rect 199 2600 921 2601
rect 199 1880 200 2600
rect 920 1880 921 2600
rect 199 1879 921 1880
rect -220 1812 -124 1828
rect 1192 1828 1208 2652
rect 1272 1828 1288 2652
rect 2604 2652 2700 2668
rect 1611 2600 2333 2601
rect 1611 1880 1612 2600
rect 2332 1880 2333 2600
rect 1611 1879 2333 1880
rect 1192 1812 1288 1828
rect 2604 1828 2620 2652
rect 2684 1828 2700 2652
rect 4016 2652 4112 2668
rect 3023 2600 3745 2601
rect 3023 1880 3024 2600
rect 3744 1880 3745 2600
rect 3023 1879 3745 1880
rect 2604 1812 2700 1828
rect 4016 1828 4032 2652
rect 4096 1828 4112 2652
rect 5428 2652 5524 2668
rect 4435 2600 5157 2601
rect 4435 1880 4436 2600
rect 5156 1880 5157 2600
rect 4435 1879 5157 1880
rect 4016 1812 4112 1828
rect 5428 1828 5444 2652
rect 5508 1828 5524 2652
rect 6840 2652 6936 2668
rect 5847 2600 6569 2601
rect 5847 1880 5848 2600
rect 6568 1880 6569 2600
rect 5847 1879 6569 1880
rect 5428 1812 5524 1828
rect 6840 1828 6856 2652
rect 6920 1828 6936 2652
rect 8252 2652 8348 2668
rect 7259 2600 7981 2601
rect 7259 1880 7260 2600
rect 7980 1880 7981 2600
rect 7259 1879 7981 1880
rect 6840 1812 6936 1828
rect 8252 1828 8268 2652
rect 8332 1828 8348 2652
rect 9664 2652 9760 2668
rect 8671 2600 9393 2601
rect 8671 1880 8672 2600
rect 9392 1880 9393 2600
rect 8671 1879 9393 1880
rect 8252 1812 8348 1828
rect 9664 1828 9680 2652
rect 9744 1828 9760 2652
rect 11076 2652 11172 2668
rect 10083 2600 10805 2601
rect 10083 1880 10084 2600
rect 10804 1880 10805 2600
rect 10083 1879 10805 1880
rect 9664 1812 9760 1828
rect 11076 1828 11092 2652
rect 11156 1828 11172 2652
rect 12488 2652 12584 2668
rect 11495 2600 12217 2601
rect 11495 1880 11496 2600
rect 12216 1880 12217 2600
rect 11495 1879 12217 1880
rect 11076 1812 11172 1828
rect 12488 1828 12504 2652
rect 12568 1828 12584 2652
rect 13900 2652 13996 2668
rect 12907 2600 13629 2601
rect 12907 1880 12908 2600
rect 13628 1880 13629 2600
rect 12907 1879 13629 1880
rect 12488 1812 12584 1828
rect 13900 1828 13916 2652
rect 13980 1828 13996 2652
rect 15312 2652 15408 2668
rect 14319 2600 15041 2601
rect 14319 1880 14320 2600
rect 15040 1880 15041 2600
rect 14319 1879 15041 1880
rect 13900 1812 13996 1828
rect 15312 1828 15328 2652
rect 15392 1828 15408 2652
rect 16724 2652 16820 2668
rect 15731 2600 16453 2601
rect 15731 1880 15732 2600
rect 16452 1880 16453 2600
rect 15731 1879 16453 1880
rect 15312 1812 15408 1828
rect 16724 1828 16740 2652
rect 16804 1828 16820 2652
rect 18136 2652 18232 2668
rect 17143 2600 17865 2601
rect 17143 1880 17144 2600
rect 17864 1880 17865 2600
rect 17143 1879 17865 1880
rect 16724 1812 16820 1828
rect 18136 1828 18152 2652
rect 18216 1828 18232 2652
rect 19548 2652 19644 2668
rect 18555 2600 19277 2601
rect 18555 1880 18556 2600
rect 19276 1880 19277 2600
rect 18555 1879 19277 1880
rect 18136 1812 18232 1828
rect 19548 1828 19564 2652
rect 19628 1828 19644 2652
rect 20960 2652 21056 2668
rect 19967 2600 20689 2601
rect 19967 1880 19968 2600
rect 20688 1880 20689 2600
rect 19967 1879 20689 1880
rect 19548 1812 19644 1828
rect 20960 1828 20976 2652
rect 21040 1828 21056 2652
rect 22372 2652 22468 2668
rect 21379 2600 22101 2601
rect 21379 1880 21380 2600
rect 22100 1880 22101 2600
rect 21379 1879 22101 1880
rect 20960 1812 21056 1828
rect 22372 1828 22388 2652
rect 22452 1828 22468 2652
rect 23784 2652 23880 2668
rect 22791 2600 23513 2601
rect 22791 1880 22792 2600
rect 23512 1880 23513 2600
rect 22791 1879 23513 1880
rect 22372 1812 22468 1828
rect 23784 1828 23800 2652
rect 23864 1828 23880 2652
rect 23784 1812 23880 1828
rect -22812 1532 -22716 1548
rect -23805 1480 -23083 1481
rect -23805 760 -23804 1480
rect -23084 760 -23083 1480
rect -23805 759 -23083 760
rect -22812 708 -22796 1532
rect -22732 708 -22716 1532
rect -21400 1532 -21304 1548
rect -22393 1480 -21671 1481
rect -22393 760 -22392 1480
rect -21672 760 -21671 1480
rect -22393 759 -21671 760
rect -22812 692 -22716 708
rect -21400 708 -21384 1532
rect -21320 708 -21304 1532
rect -19988 1532 -19892 1548
rect -20981 1480 -20259 1481
rect -20981 760 -20980 1480
rect -20260 760 -20259 1480
rect -20981 759 -20259 760
rect -21400 692 -21304 708
rect -19988 708 -19972 1532
rect -19908 708 -19892 1532
rect -18576 1532 -18480 1548
rect -19569 1480 -18847 1481
rect -19569 760 -19568 1480
rect -18848 760 -18847 1480
rect -19569 759 -18847 760
rect -19988 692 -19892 708
rect -18576 708 -18560 1532
rect -18496 708 -18480 1532
rect -17164 1532 -17068 1548
rect -18157 1480 -17435 1481
rect -18157 760 -18156 1480
rect -17436 760 -17435 1480
rect -18157 759 -17435 760
rect -18576 692 -18480 708
rect -17164 708 -17148 1532
rect -17084 708 -17068 1532
rect -15752 1532 -15656 1548
rect -16745 1480 -16023 1481
rect -16745 760 -16744 1480
rect -16024 760 -16023 1480
rect -16745 759 -16023 760
rect -17164 692 -17068 708
rect -15752 708 -15736 1532
rect -15672 708 -15656 1532
rect -14340 1532 -14244 1548
rect -15333 1480 -14611 1481
rect -15333 760 -15332 1480
rect -14612 760 -14611 1480
rect -15333 759 -14611 760
rect -15752 692 -15656 708
rect -14340 708 -14324 1532
rect -14260 708 -14244 1532
rect -12928 1532 -12832 1548
rect -13921 1480 -13199 1481
rect -13921 760 -13920 1480
rect -13200 760 -13199 1480
rect -13921 759 -13199 760
rect -14340 692 -14244 708
rect -12928 708 -12912 1532
rect -12848 708 -12832 1532
rect -11516 1532 -11420 1548
rect -12509 1480 -11787 1481
rect -12509 760 -12508 1480
rect -11788 760 -11787 1480
rect -12509 759 -11787 760
rect -12928 692 -12832 708
rect -11516 708 -11500 1532
rect -11436 708 -11420 1532
rect -10104 1532 -10008 1548
rect -11097 1480 -10375 1481
rect -11097 760 -11096 1480
rect -10376 760 -10375 1480
rect -11097 759 -10375 760
rect -11516 692 -11420 708
rect -10104 708 -10088 1532
rect -10024 708 -10008 1532
rect -8692 1532 -8596 1548
rect -9685 1480 -8963 1481
rect -9685 760 -9684 1480
rect -8964 760 -8963 1480
rect -9685 759 -8963 760
rect -10104 692 -10008 708
rect -8692 708 -8676 1532
rect -8612 708 -8596 1532
rect -7280 1532 -7184 1548
rect -8273 1480 -7551 1481
rect -8273 760 -8272 1480
rect -7552 760 -7551 1480
rect -8273 759 -7551 760
rect -8692 692 -8596 708
rect -7280 708 -7264 1532
rect -7200 708 -7184 1532
rect -5868 1532 -5772 1548
rect -6861 1480 -6139 1481
rect -6861 760 -6860 1480
rect -6140 760 -6139 1480
rect -6861 759 -6139 760
rect -7280 692 -7184 708
rect -5868 708 -5852 1532
rect -5788 708 -5772 1532
rect -4456 1532 -4360 1548
rect -5449 1480 -4727 1481
rect -5449 760 -5448 1480
rect -4728 760 -4727 1480
rect -5449 759 -4727 760
rect -5868 692 -5772 708
rect -4456 708 -4440 1532
rect -4376 708 -4360 1532
rect -3044 1532 -2948 1548
rect -4037 1480 -3315 1481
rect -4037 760 -4036 1480
rect -3316 760 -3315 1480
rect -4037 759 -3315 760
rect -4456 692 -4360 708
rect -3044 708 -3028 1532
rect -2964 708 -2948 1532
rect -1632 1532 -1536 1548
rect -2625 1480 -1903 1481
rect -2625 760 -2624 1480
rect -1904 760 -1903 1480
rect -2625 759 -1903 760
rect -3044 692 -2948 708
rect -1632 708 -1616 1532
rect -1552 708 -1536 1532
rect -220 1532 -124 1548
rect -1213 1480 -491 1481
rect -1213 760 -1212 1480
rect -492 760 -491 1480
rect -1213 759 -491 760
rect -1632 692 -1536 708
rect -220 708 -204 1532
rect -140 708 -124 1532
rect 1192 1532 1288 1548
rect 199 1480 921 1481
rect 199 760 200 1480
rect 920 760 921 1480
rect 199 759 921 760
rect -220 692 -124 708
rect 1192 708 1208 1532
rect 1272 708 1288 1532
rect 2604 1532 2700 1548
rect 1611 1480 2333 1481
rect 1611 760 1612 1480
rect 2332 760 2333 1480
rect 1611 759 2333 760
rect 1192 692 1288 708
rect 2604 708 2620 1532
rect 2684 708 2700 1532
rect 4016 1532 4112 1548
rect 3023 1480 3745 1481
rect 3023 760 3024 1480
rect 3744 760 3745 1480
rect 3023 759 3745 760
rect 2604 692 2700 708
rect 4016 708 4032 1532
rect 4096 708 4112 1532
rect 5428 1532 5524 1548
rect 4435 1480 5157 1481
rect 4435 760 4436 1480
rect 5156 760 5157 1480
rect 4435 759 5157 760
rect 4016 692 4112 708
rect 5428 708 5444 1532
rect 5508 708 5524 1532
rect 6840 1532 6936 1548
rect 5847 1480 6569 1481
rect 5847 760 5848 1480
rect 6568 760 6569 1480
rect 5847 759 6569 760
rect 5428 692 5524 708
rect 6840 708 6856 1532
rect 6920 708 6936 1532
rect 8252 1532 8348 1548
rect 7259 1480 7981 1481
rect 7259 760 7260 1480
rect 7980 760 7981 1480
rect 7259 759 7981 760
rect 6840 692 6936 708
rect 8252 708 8268 1532
rect 8332 708 8348 1532
rect 9664 1532 9760 1548
rect 8671 1480 9393 1481
rect 8671 760 8672 1480
rect 9392 760 9393 1480
rect 8671 759 9393 760
rect 8252 692 8348 708
rect 9664 708 9680 1532
rect 9744 708 9760 1532
rect 11076 1532 11172 1548
rect 10083 1480 10805 1481
rect 10083 760 10084 1480
rect 10804 760 10805 1480
rect 10083 759 10805 760
rect 9664 692 9760 708
rect 11076 708 11092 1532
rect 11156 708 11172 1532
rect 12488 1532 12584 1548
rect 11495 1480 12217 1481
rect 11495 760 11496 1480
rect 12216 760 12217 1480
rect 11495 759 12217 760
rect 11076 692 11172 708
rect 12488 708 12504 1532
rect 12568 708 12584 1532
rect 13900 1532 13996 1548
rect 12907 1480 13629 1481
rect 12907 760 12908 1480
rect 13628 760 13629 1480
rect 12907 759 13629 760
rect 12488 692 12584 708
rect 13900 708 13916 1532
rect 13980 708 13996 1532
rect 15312 1532 15408 1548
rect 14319 1480 15041 1481
rect 14319 760 14320 1480
rect 15040 760 15041 1480
rect 14319 759 15041 760
rect 13900 692 13996 708
rect 15312 708 15328 1532
rect 15392 708 15408 1532
rect 16724 1532 16820 1548
rect 15731 1480 16453 1481
rect 15731 760 15732 1480
rect 16452 760 16453 1480
rect 15731 759 16453 760
rect 15312 692 15408 708
rect 16724 708 16740 1532
rect 16804 708 16820 1532
rect 18136 1532 18232 1548
rect 17143 1480 17865 1481
rect 17143 760 17144 1480
rect 17864 760 17865 1480
rect 17143 759 17865 760
rect 16724 692 16820 708
rect 18136 708 18152 1532
rect 18216 708 18232 1532
rect 19548 1532 19644 1548
rect 18555 1480 19277 1481
rect 18555 760 18556 1480
rect 19276 760 19277 1480
rect 18555 759 19277 760
rect 18136 692 18232 708
rect 19548 708 19564 1532
rect 19628 708 19644 1532
rect 20960 1532 21056 1548
rect 19967 1480 20689 1481
rect 19967 760 19968 1480
rect 20688 760 20689 1480
rect 19967 759 20689 760
rect 19548 692 19644 708
rect 20960 708 20976 1532
rect 21040 708 21056 1532
rect 22372 1532 22468 1548
rect 21379 1480 22101 1481
rect 21379 760 21380 1480
rect 22100 760 22101 1480
rect 21379 759 22101 760
rect 20960 692 21056 708
rect 22372 708 22388 1532
rect 22452 708 22468 1532
rect 23784 1532 23880 1548
rect 22791 1480 23513 1481
rect 22791 760 22792 1480
rect 23512 760 23513 1480
rect 22791 759 23513 760
rect 22372 692 22468 708
rect 23784 708 23800 1532
rect 23864 708 23880 1532
rect 23784 692 23880 708
rect -22812 412 -22716 428
rect -23805 360 -23083 361
rect -23805 -360 -23804 360
rect -23084 -360 -23083 360
rect -23805 -361 -23083 -360
rect -22812 -412 -22796 412
rect -22732 -412 -22716 412
rect -21400 412 -21304 428
rect -22393 360 -21671 361
rect -22393 -360 -22392 360
rect -21672 -360 -21671 360
rect -22393 -361 -21671 -360
rect -22812 -428 -22716 -412
rect -21400 -412 -21384 412
rect -21320 -412 -21304 412
rect -19988 412 -19892 428
rect -20981 360 -20259 361
rect -20981 -360 -20980 360
rect -20260 -360 -20259 360
rect -20981 -361 -20259 -360
rect -21400 -428 -21304 -412
rect -19988 -412 -19972 412
rect -19908 -412 -19892 412
rect -18576 412 -18480 428
rect -19569 360 -18847 361
rect -19569 -360 -19568 360
rect -18848 -360 -18847 360
rect -19569 -361 -18847 -360
rect -19988 -428 -19892 -412
rect -18576 -412 -18560 412
rect -18496 -412 -18480 412
rect -17164 412 -17068 428
rect -18157 360 -17435 361
rect -18157 -360 -18156 360
rect -17436 -360 -17435 360
rect -18157 -361 -17435 -360
rect -18576 -428 -18480 -412
rect -17164 -412 -17148 412
rect -17084 -412 -17068 412
rect -15752 412 -15656 428
rect -16745 360 -16023 361
rect -16745 -360 -16744 360
rect -16024 -360 -16023 360
rect -16745 -361 -16023 -360
rect -17164 -428 -17068 -412
rect -15752 -412 -15736 412
rect -15672 -412 -15656 412
rect -14340 412 -14244 428
rect -15333 360 -14611 361
rect -15333 -360 -15332 360
rect -14612 -360 -14611 360
rect -15333 -361 -14611 -360
rect -15752 -428 -15656 -412
rect -14340 -412 -14324 412
rect -14260 -412 -14244 412
rect -12928 412 -12832 428
rect -13921 360 -13199 361
rect -13921 -360 -13920 360
rect -13200 -360 -13199 360
rect -13921 -361 -13199 -360
rect -14340 -428 -14244 -412
rect -12928 -412 -12912 412
rect -12848 -412 -12832 412
rect -11516 412 -11420 428
rect -12509 360 -11787 361
rect -12509 -360 -12508 360
rect -11788 -360 -11787 360
rect -12509 -361 -11787 -360
rect -12928 -428 -12832 -412
rect -11516 -412 -11500 412
rect -11436 -412 -11420 412
rect -10104 412 -10008 428
rect -11097 360 -10375 361
rect -11097 -360 -11096 360
rect -10376 -360 -10375 360
rect -11097 -361 -10375 -360
rect -11516 -428 -11420 -412
rect -10104 -412 -10088 412
rect -10024 -412 -10008 412
rect -8692 412 -8596 428
rect -9685 360 -8963 361
rect -9685 -360 -9684 360
rect -8964 -360 -8963 360
rect -9685 -361 -8963 -360
rect -10104 -428 -10008 -412
rect -8692 -412 -8676 412
rect -8612 -412 -8596 412
rect -7280 412 -7184 428
rect -8273 360 -7551 361
rect -8273 -360 -8272 360
rect -7552 -360 -7551 360
rect -8273 -361 -7551 -360
rect -8692 -428 -8596 -412
rect -7280 -412 -7264 412
rect -7200 -412 -7184 412
rect -5868 412 -5772 428
rect -6861 360 -6139 361
rect -6861 -360 -6860 360
rect -6140 -360 -6139 360
rect -6861 -361 -6139 -360
rect -7280 -428 -7184 -412
rect -5868 -412 -5852 412
rect -5788 -412 -5772 412
rect -4456 412 -4360 428
rect -5449 360 -4727 361
rect -5449 -360 -5448 360
rect -4728 -360 -4727 360
rect -5449 -361 -4727 -360
rect -5868 -428 -5772 -412
rect -4456 -412 -4440 412
rect -4376 -412 -4360 412
rect -3044 412 -2948 428
rect -4037 360 -3315 361
rect -4037 -360 -4036 360
rect -3316 -360 -3315 360
rect -4037 -361 -3315 -360
rect -4456 -428 -4360 -412
rect -3044 -412 -3028 412
rect -2964 -412 -2948 412
rect -1632 412 -1536 428
rect -2625 360 -1903 361
rect -2625 -360 -2624 360
rect -1904 -360 -1903 360
rect -2625 -361 -1903 -360
rect -3044 -428 -2948 -412
rect -1632 -412 -1616 412
rect -1552 -412 -1536 412
rect -220 412 -124 428
rect -1213 360 -491 361
rect -1213 -360 -1212 360
rect -492 -360 -491 360
rect -1213 -361 -491 -360
rect -1632 -428 -1536 -412
rect -220 -412 -204 412
rect -140 -412 -124 412
rect 1192 412 1288 428
rect 199 360 921 361
rect 199 -360 200 360
rect 920 -360 921 360
rect 199 -361 921 -360
rect -220 -428 -124 -412
rect 1192 -412 1208 412
rect 1272 -412 1288 412
rect 2604 412 2700 428
rect 1611 360 2333 361
rect 1611 -360 1612 360
rect 2332 -360 2333 360
rect 1611 -361 2333 -360
rect 1192 -428 1288 -412
rect 2604 -412 2620 412
rect 2684 -412 2700 412
rect 4016 412 4112 428
rect 3023 360 3745 361
rect 3023 -360 3024 360
rect 3744 -360 3745 360
rect 3023 -361 3745 -360
rect 2604 -428 2700 -412
rect 4016 -412 4032 412
rect 4096 -412 4112 412
rect 5428 412 5524 428
rect 4435 360 5157 361
rect 4435 -360 4436 360
rect 5156 -360 5157 360
rect 4435 -361 5157 -360
rect 4016 -428 4112 -412
rect 5428 -412 5444 412
rect 5508 -412 5524 412
rect 6840 412 6936 428
rect 5847 360 6569 361
rect 5847 -360 5848 360
rect 6568 -360 6569 360
rect 5847 -361 6569 -360
rect 5428 -428 5524 -412
rect 6840 -412 6856 412
rect 6920 -412 6936 412
rect 8252 412 8348 428
rect 7259 360 7981 361
rect 7259 -360 7260 360
rect 7980 -360 7981 360
rect 7259 -361 7981 -360
rect 6840 -428 6936 -412
rect 8252 -412 8268 412
rect 8332 -412 8348 412
rect 9664 412 9760 428
rect 8671 360 9393 361
rect 8671 -360 8672 360
rect 9392 -360 9393 360
rect 8671 -361 9393 -360
rect 8252 -428 8348 -412
rect 9664 -412 9680 412
rect 9744 -412 9760 412
rect 11076 412 11172 428
rect 10083 360 10805 361
rect 10083 -360 10084 360
rect 10804 -360 10805 360
rect 10083 -361 10805 -360
rect 9664 -428 9760 -412
rect 11076 -412 11092 412
rect 11156 -412 11172 412
rect 12488 412 12584 428
rect 11495 360 12217 361
rect 11495 -360 11496 360
rect 12216 -360 12217 360
rect 11495 -361 12217 -360
rect 11076 -428 11172 -412
rect 12488 -412 12504 412
rect 12568 -412 12584 412
rect 13900 412 13996 428
rect 12907 360 13629 361
rect 12907 -360 12908 360
rect 13628 -360 13629 360
rect 12907 -361 13629 -360
rect 12488 -428 12584 -412
rect 13900 -412 13916 412
rect 13980 -412 13996 412
rect 15312 412 15408 428
rect 14319 360 15041 361
rect 14319 -360 14320 360
rect 15040 -360 15041 360
rect 14319 -361 15041 -360
rect 13900 -428 13996 -412
rect 15312 -412 15328 412
rect 15392 -412 15408 412
rect 16724 412 16820 428
rect 15731 360 16453 361
rect 15731 -360 15732 360
rect 16452 -360 16453 360
rect 15731 -361 16453 -360
rect 15312 -428 15408 -412
rect 16724 -412 16740 412
rect 16804 -412 16820 412
rect 18136 412 18232 428
rect 17143 360 17865 361
rect 17143 -360 17144 360
rect 17864 -360 17865 360
rect 17143 -361 17865 -360
rect 16724 -428 16820 -412
rect 18136 -412 18152 412
rect 18216 -412 18232 412
rect 19548 412 19644 428
rect 18555 360 19277 361
rect 18555 -360 18556 360
rect 19276 -360 19277 360
rect 18555 -361 19277 -360
rect 18136 -428 18232 -412
rect 19548 -412 19564 412
rect 19628 -412 19644 412
rect 20960 412 21056 428
rect 19967 360 20689 361
rect 19967 -360 19968 360
rect 20688 -360 20689 360
rect 19967 -361 20689 -360
rect 19548 -428 19644 -412
rect 20960 -412 20976 412
rect 21040 -412 21056 412
rect 22372 412 22468 428
rect 21379 360 22101 361
rect 21379 -360 21380 360
rect 22100 -360 22101 360
rect 21379 -361 22101 -360
rect 20960 -428 21056 -412
rect 22372 -412 22388 412
rect 22452 -412 22468 412
rect 23784 412 23880 428
rect 22791 360 23513 361
rect 22791 -360 22792 360
rect 23512 -360 23513 360
rect 22791 -361 23513 -360
rect 22372 -428 22468 -412
rect 23784 -412 23800 412
rect 23864 -412 23880 412
rect 23784 -428 23880 -412
rect -22812 -708 -22716 -692
rect -23805 -760 -23083 -759
rect -23805 -1480 -23804 -760
rect -23084 -1480 -23083 -760
rect -23805 -1481 -23083 -1480
rect -22812 -1532 -22796 -708
rect -22732 -1532 -22716 -708
rect -21400 -708 -21304 -692
rect -22393 -760 -21671 -759
rect -22393 -1480 -22392 -760
rect -21672 -1480 -21671 -760
rect -22393 -1481 -21671 -1480
rect -22812 -1548 -22716 -1532
rect -21400 -1532 -21384 -708
rect -21320 -1532 -21304 -708
rect -19988 -708 -19892 -692
rect -20981 -760 -20259 -759
rect -20981 -1480 -20980 -760
rect -20260 -1480 -20259 -760
rect -20981 -1481 -20259 -1480
rect -21400 -1548 -21304 -1532
rect -19988 -1532 -19972 -708
rect -19908 -1532 -19892 -708
rect -18576 -708 -18480 -692
rect -19569 -760 -18847 -759
rect -19569 -1480 -19568 -760
rect -18848 -1480 -18847 -760
rect -19569 -1481 -18847 -1480
rect -19988 -1548 -19892 -1532
rect -18576 -1532 -18560 -708
rect -18496 -1532 -18480 -708
rect -17164 -708 -17068 -692
rect -18157 -760 -17435 -759
rect -18157 -1480 -18156 -760
rect -17436 -1480 -17435 -760
rect -18157 -1481 -17435 -1480
rect -18576 -1548 -18480 -1532
rect -17164 -1532 -17148 -708
rect -17084 -1532 -17068 -708
rect -15752 -708 -15656 -692
rect -16745 -760 -16023 -759
rect -16745 -1480 -16744 -760
rect -16024 -1480 -16023 -760
rect -16745 -1481 -16023 -1480
rect -17164 -1548 -17068 -1532
rect -15752 -1532 -15736 -708
rect -15672 -1532 -15656 -708
rect -14340 -708 -14244 -692
rect -15333 -760 -14611 -759
rect -15333 -1480 -15332 -760
rect -14612 -1480 -14611 -760
rect -15333 -1481 -14611 -1480
rect -15752 -1548 -15656 -1532
rect -14340 -1532 -14324 -708
rect -14260 -1532 -14244 -708
rect -12928 -708 -12832 -692
rect -13921 -760 -13199 -759
rect -13921 -1480 -13920 -760
rect -13200 -1480 -13199 -760
rect -13921 -1481 -13199 -1480
rect -14340 -1548 -14244 -1532
rect -12928 -1532 -12912 -708
rect -12848 -1532 -12832 -708
rect -11516 -708 -11420 -692
rect -12509 -760 -11787 -759
rect -12509 -1480 -12508 -760
rect -11788 -1480 -11787 -760
rect -12509 -1481 -11787 -1480
rect -12928 -1548 -12832 -1532
rect -11516 -1532 -11500 -708
rect -11436 -1532 -11420 -708
rect -10104 -708 -10008 -692
rect -11097 -760 -10375 -759
rect -11097 -1480 -11096 -760
rect -10376 -1480 -10375 -760
rect -11097 -1481 -10375 -1480
rect -11516 -1548 -11420 -1532
rect -10104 -1532 -10088 -708
rect -10024 -1532 -10008 -708
rect -8692 -708 -8596 -692
rect -9685 -760 -8963 -759
rect -9685 -1480 -9684 -760
rect -8964 -1480 -8963 -760
rect -9685 -1481 -8963 -1480
rect -10104 -1548 -10008 -1532
rect -8692 -1532 -8676 -708
rect -8612 -1532 -8596 -708
rect -7280 -708 -7184 -692
rect -8273 -760 -7551 -759
rect -8273 -1480 -8272 -760
rect -7552 -1480 -7551 -760
rect -8273 -1481 -7551 -1480
rect -8692 -1548 -8596 -1532
rect -7280 -1532 -7264 -708
rect -7200 -1532 -7184 -708
rect -5868 -708 -5772 -692
rect -6861 -760 -6139 -759
rect -6861 -1480 -6860 -760
rect -6140 -1480 -6139 -760
rect -6861 -1481 -6139 -1480
rect -7280 -1548 -7184 -1532
rect -5868 -1532 -5852 -708
rect -5788 -1532 -5772 -708
rect -4456 -708 -4360 -692
rect -5449 -760 -4727 -759
rect -5449 -1480 -5448 -760
rect -4728 -1480 -4727 -760
rect -5449 -1481 -4727 -1480
rect -5868 -1548 -5772 -1532
rect -4456 -1532 -4440 -708
rect -4376 -1532 -4360 -708
rect -3044 -708 -2948 -692
rect -4037 -760 -3315 -759
rect -4037 -1480 -4036 -760
rect -3316 -1480 -3315 -760
rect -4037 -1481 -3315 -1480
rect -4456 -1548 -4360 -1532
rect -3044 -1532 -3028 -708
rect -2964 -1532 -2948 -708
rect -1632 -708 -1536 -692
rect -2625 -760 -1903 -759
rect -2625 -1480 -2624 -760
rect -1904 -1480 -1903 -760
rect -2625 -1481 -1903 -1480
rect -3044 -1548 -2948 -1532
rect -1632 -1532 -1616 -708
rect -1552 -1532 -1536 -708
rect -220 -708 -124 -692
rect -1213 -760 -491 -759
rect -1213 -1480 -1212 -760
rect -492 -1480 -491 -760
rect -1213 -1481 -491 -1480
rect -1632 -1548 -1536 -1532
rect -220 -1532 -204 -708
rect -140 -1532 -124 -708
rect 1192 -708 1288 -692
rect 199 -760 921 -759
rect 199 -1480 200 -760
rect 920 -1480 921 -760
rect 199 -1481 921 -1480
rect -220 -1548 -124 -1532
rect 1192 -1532 1208 -708
rect 1272 -1532 1288 -708
rect 2604 -708 2700 -692
rect 1611 -760 2333 -759
rect 1611 -1480 1612 -760
rect 2332 -1480 2333 -760
rect 1611 -1481 2333 -1480
rect 1192 -1548 1288 -1532
rect 2604 -1532 2620 -708
rect 2684 -1532 2700 -708
rect 4016 -708 4112 -692
rect 3023 -760 3745 -759
rect 3023 -1480 3024 -760
rect 3744 -1480 3745 -760
rect 3023 -1481 3745 -1480
rect 2604 -1548 2700 -1532
rect 4016 -1532 4032 -708
rect 4096 -1532 4112 -708
rect 5428 -708 5524 -692
rect 4435 -760 5157 -759
rect 4435 -1480 4436 -760
rect 5156 -1480 5157 -760
rect 4435 -1481 5157 -1480
rect 4016 -1548 4112 -1532
rect 5428 -1532 5444 -708
rect 5508 -1532 5524 -708
rect 6840 -708 6936 -692
rect 5847 -760 6569 -759
rect 5847 -1480 5848 -760
rect 6568 -1480 6569 -760
rect 5847 -1481 6569 -1480
rect 5428 -1548 5524 -1532
rect 6840 -1532 6856 -708
rect 6920 -1532 6936 -708
rect 8252 -708 8348 -692
rect 7259 -760 7981 -759
rect 7259 -1480 7260 -760
rect 7980 -1480 7981 -760
rect 7259 -1481 7981 -1480
rect 6840 -1548 6936 -1532
rect 8252 -1532 8268 -708
rect 8332 -1532 8348 -708
rect 9664 -708 9760 -692
rect 8671 -760 9393 -759
rect 8671 -1480 8672 -760
rect 9392 -1480 9393 -760
rect 8671 -1481 9393 -1480
rect 8252 -1548 8348 -1532
rect 9664 -1532 9680 -708
rect 9744 -1532 9760 -708
rect 11076 -708 11172 -692
rect 10083 -760 10805 -759
rect 10083 -1480 10084 -760
rect 10804 -1480 10805 -760
rect 10083 -1481 10805 -1480
rect 9664 -1548 9760 -1532
rect 11076 -1532 11092 -708
rect 11156 -1532 11172 -708
rect 12488 -708 12584 -692
rect 11495 -760 12217 -759
rect 11495 -1480 11496 -760
rect 12216 -1480 12217 -760
rect 11495 -1481 12217 -1480
rect 11076 -1548 11172 -1532
rect 12488 -1532 12504 -708
rect 12568 -1532 12584 -708
rect 13900 -708 13996 -692
rect 12907 -760 13629 -759
rect 12907 -1480 12908 -760
rect 13628 -1480 13629 -760
rect 12907 -1481 13629 -1480
rect 12488 -1548 12584 -1532
rect 13900 -1532 13916 -708
rect 13980 -1532 13996 -708
rect 15312 -708 15408 -692
rect 14319 -760 15041 -759
rect 14319 -1480 14320 -760
rect 15040 -1480 15041 -760
rect 14319 -1481 15041 -1480
rect 13900 -1548 13996 -1532
rect 15312 -1532 15328 -708
rect 15392 -1532 15408 -708
rect 16724 -708 16820 -692
rect 15731 -760 16453 -759
rect 15731 -1480 15732 -760
rect 16452 -1480 16453 -760
rect 15731 -1481 16453 -1480
rect 15312 -1548 15408 -1532
rect 16724 -1532 16740 -708
rect 16804 -1532 16820 -708
rect 18136 -708 18232 -692
rect 17143 -760 17865 -759
rect 17143 -1480 17144 -760
rect 17864 -1480 17865 -760
rect 17143 -1481 17865 -1480
rect 16724 -1548 16820 -1532
rect 18136 -1532 18152 -708
rect 18216 -1532 18232 -708
rect 19548 -708 19644 -692
rect 18555 -760 19277 -759
rect 18555 -1480 18556 -760
rect 19276 -1480 19277 -760
rect 18555 -1481 19277 -1480
rect 18136 -1548 18232 -1532
rect 19548 -1532 19564 -708
rect 19628 -1532 19644 -708
rect 20960 -708 21056 -692
rect 19967 -760 20689 -759
rect 19967 -1480 19968 -760
rect 20688 -1480 20689 -760
rect 19967 -1481 20689 -1480
rect 19548 -1548 19644 -1532
rect 20960 -1532 20976 -708
rect 21040 -1532 21056 -708
rect 22372 -708 22468 -692
rect 21379 -760 22101 -759
rect 21379 -1480 21380 -760
rect 22100 -1480 22101 -760
rect 21379 -1481 22101 -1480
rect 20960 -1548 21056 -1532
rect 22372 -1532 22388 -708
rect 22452 -1532 22468 -708
rect 23784 -708 23880 -692
rect 22791 -760 23513 -759
rect 22791 -1480 22792 -760
rect 23512 -1480 23513 -760
rect 22791 -1481 23513 -1480
rect 22372 -1548 22468 -1532
rect 23784 -1532 23800 -708
rect 23864 -1532 23880 -708
rect 23784 -1548 23880 -1532
rect -22812 -1828 -22716 -1812
rect -23805 -1880 -23083 -1879
rect -23805 -2600 -23804 -1880
rect -23084 -2600 -23083 -1880
rect -23805 -2601 -23083 -2600
rect -22812 -2652 -22796 -1828
rect -22732 -2652 -22716 -1828
rect -21400 -1828 -21304 -1812
rect -22393 -1880 -21671 -1879
rect -22393 -2600 -22392 -1880
rect -21672 -2600 -21671 -1880
rect -22393 -2601 -21671 -2600
rect -22812 -2668 -22716 -2652
rect -21400 -2652 -21384 -1828
rect -21320 -2652 -21304 -1828
rect -19988 -1828 -19892 -1812
rect -20981 -1880 -20259 -1879
rect -20981 -2600 -20980 -1880
rect -20260 -2600 -20259 -1880
rect -20981 -2601 -20259 -2600
rect -21400 -2668 -21304 -2652
rect -19988 -2652 -19972 -1828
rect -19908 -2652 -19892 -1828
rect -18576 -1828 -18480 -1812
rect -19569 -1880 -18847 -1879
rect -19569 -2600 -19568 -1880
rect -18848 -2600 -18847 -1880
rect -19569 -2601 -18847 -2600
rect -19988 -2668 -19892 -2652
rect -18576 -2652 -18560 -1828
rect -18496 -2652 -18480 -1828
rect -17164 -1828 -17068 -1812
rect -18157 -1880 -17435 -1879
rect -18157 -2600 -18156 -1880
rect -17436 -2600 -17435 -1880
rect -18157 -2601 -17435 -2600
rect -18576 -2668 -18480 -2652
rect -17164 -2652 -17148 -1828
rect -17084 -2652 -17068 -1828
rect -15752 -1828 -15656 -1812
rect -16745 -1880 -16023 -1879
rect -16745 -2600 -16744 -1880
rect -16024 -2600 -16023 -1880
rect -16745 -2601 -16023 -2600
rect -17164 -2668 -17068 -2652
rect -15752 -2652 -15736 -1828
rect -15672 -2652 -15656 -1828
rect -14340 -1828 -14244 -1812
rect -15333 -1880 -14611 -1879
rect -15333 -2600 -15332 -1880
rect -14612 -2600 -14611 -1880
rect -15333 -2601 -14611 -2600
rect -15752 -2668 -15656 -2652
rect -14340 -2652 -14324 -1828
rect -14260 -2652 -14244 -1828
rect -12928 -1828 -12832 -1812
rect -13921 -1880 -13199 -1879
rect -13921 -2600 -13920 -1880
rect -13200 -2600 -13199 -1880
rect -13921 -2601 -13199 -2600
rect -14340 -2668 -14244 -2652
rect -12928 -2652 -12912 -1828
rect -12848 -2652 -12832 -1828
rect -11516 -1828 -11420 -1812
rect -12509 -1880 -11787 -1879
rect -12509 -2600 -12508 -1880
rect -11788 -2600 -11787 -1880
rect -12509 -2601 -11787 -2600
rect -12928 -2668 -12832 -2652
rect -11516 -2652 -11500 -1828
rect -11436 -2652 -11420 -1828
rect -10104 -1828 -10008 -1812
rect -11097 -1880 -10375 -1879
rect -11097 -2600 -11096 -1880
rect -10376 -2600 -10375 -1880
rect -11097 -2601 -10375 -2600
rect -11516 -2668 -11420 -2652
rect -10104 -2652 -10088 -1828
rect -10024 -2652 -10008 -1828
rect -8692 -1828 -8596 -1812
rect -9685 -1880 -8963 -1879
rect -9685 -2600 -9684 -1880
rect -8964 -2600 -8963 -1880
rect -9685 -2601 -8963 -2600
rect -10104 -2668 -10008 -2652
rect -8692 -2652 -8676 -1828
rect -8612 -2652 -8596 -1828
rect -7280 -1828 -7184 -1812
rect -8273 -1880 -7551 -1879
rect -8273 -2600 -8272 -1880
rect -7552 -2600 -7551 -1880
rect -8273 -2601 -7551 -2600
rect -8692 -2668 -8596 -2652
rect -7280 -2652 -7264 -1828
rect -7200 -2652 -7184 -1828
rect -5868 -1828 -5772 -1812
rect -6861 -1880 -6139 -1879
rect -6861 -2600 -6860 -1880
rect -6140 -2600 -6139 -1880
rect -6861 -2601 -6139 -2600
rect -7280 -2668 -7184 -2652
rect -5868 -2652 -5852 -1828
rect -5788 -2652 -5772 -1828
rect -4456 -1828 -4360 -1812
rect -5449 -1880 -4727 -1879
rect -5449 -2600 -5448 -1880
rect -4728 -2600 -4727 -1880
rect -5449 -2601 -4727 -2600
rect -5868 -2668 -5772 -2652
rect -4456 -2652 -4440 -1828
rect -4376 -2652 -4360 -1828
rect -3044 -1828 -2948 -1812
rect -4037 -1880 -3315 -1879
rect -4037 -2600 -4036 -1880
rect -3316 -2600 -3315 -1880
rect -4037 -2601 -3315 -2600
rect -4456 -2668 -4360 -2652
rect -3044 -2652 -3028 -1828
rect -2964 -2652 -2948 -1828
rect -1632 -1828 -1536 -1812
rect -2625 -1880 -1903 -1879
rect -2625 -2600 -2624 -1880
rect -1904 -2600 -1903 -1880
rect -2625 -2601 -1903 -2600
rect -3044 -2668 -2948 -2652
rect -1632 -2652 -1616 -1828
rect -1552 -2652 -1536 -1828
rect -220 -1828 -124 -1812
rect -1213 -1880 -491 -1879
rect -1213 -2600 -1212 -1880
rect -492 -2600 -491 -1880
rect -1213 -2601 -491 -2600
rect -1632 -2668 -1536 -2652
rect -220 -2652 -204 -1828
rect -140 -2652 -124 -1828
rect 1192 -1828 1288 -1812
rect 199 -1880 921 -1879
rect 199 -2600 200 -1880
rect 920 -2600 921 -1880
rect 199 -2601 921 -2600
rect -220 -2668 -124 -2652
rect 1192 -2652 1208 -1828
rect 1272 -2652 1288 -1828
rect 2604 -1828 2700 -1812
rect 1611 -1880 2333 -1879
rect 1611 -2600 1612 -1880
rect 2332 -2600 2333 -1880
rect 1611 -2601 2333 -2600
rect 1192 -2668 1288 -2652
rect 2604 -2652 2620 -1828
rect 2684 -2652 2700 -1828
rect 4016 -1828 4112 -1812
rect 3023 -1880 3745 -1879
rect 3023 -2600 3024 -1880
rect 3744 -2600 3745 -1880
rect 3023 -2601 3745 -2600
rect 2604 -2668 2700 -2652
rect 4016 -2652 4032 -1828
rect 4096 -2652 4112 -1828
rect 5428 -1828 5524 -1812
rect 4435 -1880 5157 -1879
rect 4435 -2600 4436 -1880
rect 5156 -2600 5157 -1880
rect 4435 -2601 5157 -2600
rect 4016 -2668 4112 -2652
rect 5428 -2652 5444 -1828
rect 5508 -2652 5524 -1828
rect 6840 -1828 6936 -1812
rect 5847 -1880 6569 -1879
rect 5847 -2600 5848 -1880
rect 6568 -2600 6569 -1880
rect 5847 -2601 6569 -2600
rect 5428 -2668 5524 -2652
rect 6840 -2652 6856 -1828
rect 6920 -2652 6936 -1828
rect 8252 -1828 8348 -1812
rect 7259 -1880 7981 -1879
rect 7259 -2600 7260 -1880
rect 7980 -2600 7981 -1880
rect 7259 -2601 7981 -2600
rect 6840 -2668 6936 -2652
rect 8252 -2652 8268 -1828
rect 8332 -2652 8348 -1828
rect 9664 -1828 9760 -1812
rect 8671 -1880 9393 -1879
rect 8671 -2600 8672 -1880
rect 9392 -2600 9393 -1880
rect 8671 -2601 9393 -2600
rect 8252 -2668 8348 -2652
rect 9664 -2652 9680 -1828
rect 9744 -2652 9760 -1828
rect 11076 -1828 11172 -1812
rect 10083 -1880 10805 -1879
rect 10083 -2600 10084 -1880
rect 10804 -2600 10805 -1880
rect 10083 -2601 10805 -2600
rect 9664 -2668 9760 -2652
rect 11076 -2652 11092 -1828
rect 11156 -2652 11172 -1828
rect 12488 -1828 12584 -1812
rect 11495 -1880 12217 -1879
rect 11495 -2600 11496 -1880
rect 12216 -2600 12217 -1880
rect 11495 -2601 12217 -2600
rect 11076 -2668 11172 -2652
rect 12488 -2652 12504 -1828
rect 12568 -2652 12584 -1828
rect 13900 -1828 13996 -1812
rect 12907 -1880 13629 -1879
rect 12907 -2600 12908 -1880
rect 13628 -2600 13629 -1880
rect 12907 -2601 13629 -2600
rect 12488 -2668 12584 -2652
rect 13900 -2652 13916 -1828
rect 13980 -2652 13996 -1828
rect 15312 -1828 15408 -1812
rect 14319 -1880 15041 -1879
rect 14319 -2600 14320 -1880
rect 15040 -2600 15041 -1880
rect 14319 -2601 15041 -2600
rect 13900 -2668 13996 -2652
rect 15312 -2652 15328 -1828
rect 15392 -2652 15408 -1828
rect 16724 -1828 16820 -1812
rect 15731 -1880 16453 -1879
rect 15731 -2600 15732 -1880
rect 16452 -2600 16453 -1880
rect 15731 -2601 16453 -2600
rect 15312 -2668 15408 -2652
rect 16724 -2652 16740 -1828
rect 16804 -2652 16820 -1828
rect 18136 -1828 18232 -1812
rect 17143 -1880 17865 -1879
rect 17143 -2600 17144 -1880
rect 17864 -2600 17865 -1880
rect 17143 -2601 17865 -2600
rect 16724 -2668 16820 -2652
rect 18136 -2652 18152 -1828
rect 18216 -2652 18232 -1828
rect 19548 -1828 19644 -1812
rect 18555 -1880 19277 -1879
rect 18555 -2600 18556 -1880
rect 19276 -2600 19277 -1880
rect 18555 -2601 19277 -2600
rect 18136 -2668 18232 -2652
rect 19548 -2652 19564 -1828
rect 19628 -2652 19644 -1828
rect 20960 -1828 21056 -1812
rect 19967 -1880 20689 -1879
rect 19967 -2600 19968 -1880
rect 20688 -2600 20689 -1880
rect 19967 -2601 20689 -2600
rect 19548 -2668 19644 -2652
rect 20960 -2652 20976 -1828
rect 21040 -2652 21056 -1828
rect 22372 -1828 22468 -1812
rect 21379 -1880 22101 -1879
rect 21379 -2600 21380 -1880
rect 22100 -2600 22101 -1880
rect 21379 -2601 22101 -2600
rect 20960 -2668 21056 -2652
rect 22372 -2652 22388 -1828
rect 22452 -2652 22468 -1828
rect 23784 -1828 23880 -1812
rect 22791 -1880 23513 -1879
rect 22791 -2600 22792 -1880
rect 23512 -2600 23513 -1880
rect 22791 -2601 23513 -2600
rect 22372 -2668 22468 -2652
rect 23784 -2652 23800 -1828
rect 23864 -2652 23880 -1828
rect 23784 -2668 23880 -2652
rect -22812 -2948 -22716 -2932
rect -23805 -3000 -23083 -2999
rect -23805 -3720 -23804 -3000
rect -23084 -3720 -23083 -3000
rect -23805 -3721 -23083 -3720
rect -22812 -3772 -22796 -2948
rect -22732 -3772 -22716 -2948
rect -21400 -2948 -21304 -2932
rect -22393 -3000 -21671 -2999
rect -22393 -3720 -22392 -3000
rect -21672 -3720 -21671 -3000
rect -22393 -3721 -21671 -3720
rect -22812 -3788 -22716 -3772
rect -21400 -3772 -21384 -2948
rect -21320 -3772 -21304 -2948
rect -19988 -2948 -19892 -2932
rect -20981 -3000 -20259 -2999
rect -20981 -3720 -20980 -3000
rect -20260 -3720 -20259 -3000
rect -20981 -3721 -20259 -3720
rect -21400 -3788 -21304 -3772
rect -19988 -3772 -19972 -2948
rect -19908 -3772 -19892 -2948
rect -18576 -2948 -18480 -2932
rect -19569 -3000 -18847 -2999
rect -19569 -3720 -19568 -3000
rect -18848 -3720 -18847 -3000
rect -19569 -3721 -18847 -3720
rect -19988 -3788 -19892 -3772
rect -18576 -3772 -18560 -2948
rect -18496 -3772 -18480 -2948
rect -17164 -2948 -17068 -2932
rect -18157 -3000 -17435 -2999
rect -18157 -3720 -18156 -3000
rect -17436 -3720 -17435 -3000
rect -18157 -3721 -17435 -3720
rect -18576 -3788 -18480 -3772
rect -17164 -3772 -17148 -2948
rect -17084 -3772 -17068 -2948
rect -15752 -2948 -15656 -2932
rect -16745 -3000 -16023 -2999
rect -16745 -3720 -16744 -3000
rect -16024 -3720 -16023 -3000
rect -16745 -3721 -16023 -3720
rect -17164 -3788 -17068 -3772
rect -15752 -3772 -15736 -2948
rect -15672 -3772 -15656 -2948
rect -14340 -2948 -14244 -2932
rect -15333 -3000 -14611 -2999
rect -15333 -3720 -15332 -3000
rect -14612 -3720 -14611 -3000
rect -15333 -3721 -14611 -3720
rect -15752 -3788 -15656 -3772
rect -14340 -3772 -14324 -2948
rect -14260 -3772 -14244 -2948
rect -12928 -2948 -12832 -2932
rect -13921 -3000 -13199 -2999
rect -13921 -3720 -13920 -3000
rect -13200 -3720 -13199 -3000
rect -13921 -3721 -13199 -3720
rect -14340 -3788 -14244 -3772
rect -12928 -3772 -12912 -2948
rect -12848 -3772 -12832 -2948
rect -11516 -2948 -11420 -2932
rect -12509 -3000 -11787 -2999
rect -12509 -3720 -12508 -3000
rect -11788 -3720 -11787 -3000
rect -12509 -3721 -11787 -3720
rect -12928 -3788 -12832 -3772
rect -11516 -3772 -11500 -2948
rect -11436 -3772 -11420 -2948
rect -10104 -2948 -10008 -2932
rect -11097 -3000 -10375 -2999
rect -11097 -3720 -11096 -3000
rect -10376 -3720 -10375 -3000
rect -11097 -3721 -10375 -3720
rect -11516 -3788 -11420 -3772
rect -10104 -3772 -10088 -2948
rect -10024 -3772 -10008 -2948
rect -8692 -2948 -8596 -2932
rect -9685 -3000 -8963 -2999
rect -9685 -3720 -9684 -3000
rect -8964 -3720 -8963 -3000
rect -9685 -3721 -8963 -3720
rect -10104 -3788 -10008 -3772
rect -8692 -3772 -8676 -2948
rect -8612 -3772 -8596 -2948
rect -7280 -2948 -7184 -2932
rect -8273 -3000 -7551 -2999
rect -8273 -3720 -8272 -3000
rect -7552 -3720 -7551 -3000
rect -8273 -3721 -7551 -3720
rect -8692 -3788 -8596 -3772
rect -7280 -3772 -7264 -2948
rect -7200 -3772 -7184 -2948
rect -5868 -2948 -5772 -2932
rect -6861 -3000 -6139 -2999
rect -6861 -3720 -6860 -3000
rect -6140 -3720 -6139 -3000
rect -6861 -3721 -6139 -3720
rect -7280 -3788 -7184 -3772
rect -5868 -3772 -5852 -2948
rect -5788 -3772 -5772 -2948
rect -4456 -2948 -4360 -2932
rect -5449 -3000 -4727 -2999
rect -5449 -3720 -5448 -3000
rect -4728 -3720 -4727 -3000
rect -5449 -3721 -4727 -3720
rect -5868 -3788 -5772 -3772
rect -4456 -3772 -4440 -2948
rect -4376 -3772 -4360 -2948
rect -3044 -2948 -2948 -2932
rect -4037 -3000 -3315 -2999
rect -4037 -3720 -4036 -3000
rect -3316 -3720 -3315 -3000
rect -4037 -3721 -3315 -3720
rect -4456 -3788 -4360 -3772
rect -3044 -3772 -3028 -2948
rect -2964 -3772 -2948 -2948
rect -1632 -2948 -1536 -2932
rect -2625 -3000 -1903 -2999
rect -2625 -3720 -2624 -3000
rect -1904 -3720 -1903 -3000
rect -2625 -3721 -1903 -3720
rect -3044 -3788 -2948 -3772
rect -1632 -3772 -1616 -2948
rect -1552 -3772 -1536 -2948
rect -220 -2948 -124 -2932
rect -1213 -3000 -491 -2999
rect -1213 -3720 -1212 -3000
rect -492 -3720 -491 -3000
rect -1213 -3721 -491 -3720
rect -1632 -3788 -1536 -3772
rect -220 -3772 -204 -2948
rect -140 -3772 -124 -2948
rect 1192 -2948 1288 -2932
rect 199 -3000 921 -2999
rect 199 -3720 200 -3000
rect 920 -3720 921 -3000
rect 199 -3721 921 -3720
rect -220 -3788 -124 -3772
rect 1192 -3772 1208 -2948
rect 1272 -3772 1288 -2948
rect 2604 -2948 2700 -2932
rect 1611 -3000 2333 -2999
rect 1611 -3720 1612 -3000
rect 2332 -3720 2333 -3000
rect 1611 -3721 2333 -3720
rect 1192 -3788 1288 -3772
rect 2604 -3772 2620 -2948
rect 2684 -3772 2700 -2948
rect 4016 -2948 4112 -2932
rect 3023 -3000 3745 -2999
rect 3023 -3720 3024 -3000
rect 3744 -3720 3745 -3000
rect 3023 -3721 3745 -3720
rect 2604 -3788 2700 -3772
rect 4016 -3772 4032 -2948
rect 4096 -3772 4112 -2948
rect 5428 -2948 5524 -2932
rect 4435 -3000 5157 -2999
rect 4435 -3720 4436 -3000
rect 5156 -3720 5157 -3000
rect 4435 -3721 5157 -3720
rect 4016 -3788 4112 -3772
rect 5428 -3772 5444 -2948
rect 5508 -3772 5524 -2948
rect 6840 -2948 6936 -2932
rect 5847 -3000 6569 -2999
rect 5847 -3720 5848 -3000
rect 6568 -3720 6569 -3000
rect 5847 -3721 6569 -3720
rect 5428 -3788 5524 -3772
rect 6840 -3772 6856 -2948
rect 6920 -3772 6936 -2948
rect 8252 -2948 8348 -2932
rect 7259 -3000 7981 -2999
rect 7259 -3720 7260 -3000
rect 7980 -3720 7981 -3000
rect 7259 -3721 7981 -3720
rect 6840 -3788 6936 -3772
rect 8252 -3772 8268 -2948
rect 8332 -3772 8348 -2948
rect 9664 -2948 9760 -2932
rect 8671 -3000 9393 -2999
rect 8671 -3720 8672 -3000
rect 9392 -3720 9393 -3000
rect 8671 -3721 9393 -3720
rect 8252 -3788 8348 -3772
rect 9664 -3772 9680 -2948
rect 9744 -3772 9760 -2948
rect 11076 -2948 11172 -2932
rect 10083 -3000 10805 -2999
rect 10083 -3720 10084 -3000
rect 10804 -3720 10805 -3000
rect 10083 -3721 10805 -3720
rect 9664 -3788 9760 -3772
rect 11076 -3772 11092 -2948
rect 11156 -3772 11172 -2948
rect 12488 -2948 12584 -2932
rect 11495 -3000 12217 -2999
rect 11495 -3720 11496 -3000
rect 12216 -3720 12217 -3000
rect 11495 -3721 12217 -3720
rect 11076 -3788 11172 -3772
rect 12488 -3772 12504 -2948
rect 12568 -3772 12584 -2948
rect 13900 -2948 13996 -2932
rect 12907 -3000 13629 -2999
rect 12907 -3720 12908 -3000
rect 13628 -3720 13629 -3000
rect 12907 -3721 13629 -3720
rect 12488 -3788 12584 -3772
rect 13900 -3772 13916 -2948
rect 13980 -3772 13996 -2948
rect 15312 -2948 15408 -2932
rect 14319 -3000 15041 -2999
rect 14319 -3720 14320 -3000
rect 15040 -3720 15041 -3000
rect 14319 -3721 15041 -3720
rect 13900 -3788 13996 -3772
rect 15312 -3772 15328 -2948
rect 15392 -3772 15408 -2948
rect 16724 -2948 16820 -2932
rect 15731 -3000 16453 -2999
rect 15731 -3720 15732 -3000
rect 16452 -3720 16453 -3000
rect 15731 -3721 16453 -3720
rect 15312 -3788 15408 -3772
rect 16724 -3772 16740 -2948
rect 16804 -3772 16820 -2948
rect 18136 -2948 18232 -2932
rect 17143 -3000 17865 -2999
rect 17143 -3720 17144 -3000
rect 17864 -3720 17865 -3000
rect 17143 -3721 17865 -3720
rect 16724 -3788 16820 -3772
rect 18136 -3772 18152 -2948
rect 18216 -3772 18232 -2948
rect 19548 -2948 19644 -2932
rect 18555 -3000 19277 -2999
rect 18555 -3720 18556 -3000
rect 19276 -3720 19277 -3000
rect 18555 -3721 19277 -3720
rect 18136 -3788 18232 -3772
rect 19548 -3772 19564 -2948
rect 19628 -3772 19644 -2948
rect 20960 -2948 21056 -2932
rect 19967 -3000 20689 -2999
rect 19967 -3720 19968 -3000
rect 20688 -3720 20689 -3000
rect 19967 -3721 20689 -3720
rect 19548 -3788 19644 -3772
rect 20960 -3772 20976 -2948
rect 21040 -3772 21056 -2948
rect 22372 -2948 22468 -2932
rect 21379 -3000 22101 -2999
rect 21379 -3720 21380 -3000
rect 22100 -3720 22101 -3000
rect 21379 -3721 22101 -3720
rect 20960 -3788 21056 -3772
rect 22372 -3772 22388 -2948
rect 22452 -3772 22468 -2948
rect 23784 -2948 23880 -2932
rect 22791 -3000 23513 -2999
rect 22791 -3720 22792 -3000
rect 23512 -3720 23513 -3000
rect 22791 -3721 23513 -3720
rect 22372 -3788 22468 -3772
rect 23784 -3772 23800 -2948
rect 23864 -3772 23880 -2948
rect 23784 -3788 23880 -3772
rect -22812 -4068 -22716 -4052
rect -23805 -4120 -23083 -4119
rect -23805 -4840 -23804 -4120
rect -23084 -4840 -23083 -4120
rect -23805 -4841 -23083 -4840
rect -22812 -4892 -22796 -4068
rect -22732 -4892 -22716 -4068
rect -21400 -4068 -21304 -4052
rect -22393 -4120 -21671 -4119
rect -22393 -4840 -22392 -4120
rect -21672 -4840 -21671 -4120
rect -22393 -4841 -21671 -4840
rect -22812 -4908 -22716 -4892
rect -21400 -4892 -21384 -4068
rect -21320 -4892 -21304 -4068
rect -19988 -4068 -19892 -4052
rect -20981 -4120 -20259 -4119
rect -20981 -4840 -20980 -4120
rect -20260 -4840 -20259 -4120
rect -20981 -4841 -20259 -4840
rect -21400 -4908 -21304 -4892
rect -19988 -4892 -19972 -4068
rect -19908 -4892 -19892 -4068
rect -18576 -4068 -18480 -4052
rect -19569 -4120 -18847 -4119
rect -19569 -4840 -19568 -4120
rect -18848 -4840 -18847 -4120
rect -19569 -4841 -18847 -4840
rect -19988 -4908 -19892 -4892
rect -18576 -4892 -18560 -4068
rect -18496 -4892 -18480 -4068
rect -17164 -4068 -17068 -4052
rect -18157 -4120 -17435 -4119
rect -18157 -4840 -18156 -4120
rect -17436 -4840 -17435 -4120
rect -18157 -4841 -17435 -4840
rect -18576 -4908 -18480 -4892
rect -17164 -4892 -17148 -4068
rect -17084 -4892 -17068 -4068
rect -15752 -4068 -15656 -4052
rect -16745 -4120 -16023 -4119
rect -16745 -4840 -16744 -4120
rect -16024 -4840 -16023 -4120
rect -16745 -4841 -16023 -4840
rect -17164 -4908 -17068 -4892
rect -15752 -4892 -15736 -4068
rect -15672 -4892 -15656 -4068
rect -14340 -4068 -14244 -4052
rect -15333 -4120 -14611 -4119
rect -15333 -4840 -15332 -4120
rect -14612 -4840 -14611 -4120
rect -15333 -4841 -14611 -4840
rect -15752 -4908 -15656 -4892
rect -14340 -4892 -14324 -4068
rect -14260 -4892 -14244 -4068
rect -12928 -4068 -12832 -4052
rect -13921 -4120 -13199 -4119
rect -13921 -4840 -13920 -4120
rect -13200 -4840 -13199 -4120
rect -13921 -4841 -13199 -4840
rect -14340 -4908 -14244 -4892
rect -12928 -4892 -12912 -4068
rect -12848 -4892 -12832 -4068
rect -11516 -4068 -11420 -4052
rect -12509 -4120 -11787 -4119
rect -12509 -4840 -12508 -4120
rect -11788 -4840 -11787 -4120
rect -12509 -4841 -11787 -4840
rect -12928 -4908 -12832 -4892
rect -11516 -4892 -11500 -4068
rect -11436 -4892 -11420 -4068
rect -10104 -4068 -10008 -4052
rect -11097 -4120 -10375 -4119
rect -11097 -4840 -11096 -4120
rect -10376 -4840 -10375 -4120
rect -11097 -4841 -10375 -4840
rect -11516 -4908 -11420 -4892
rect -10104 -4892 -10088 -4068
rect -10024 -4892 -10008 -4068
rect -8692 -4068 -8596 -4052
rect -9685 -4120 -8963 -4119
rect -9685 -4840 -9684 -4120
rect -8964 -4840 -8963 -4120
rect -9685 -4841 -8963 -4840
rect -10104 -4908 -10008 -4892
rect -8692 -4892 -8676 -4068
rect -8612 -4892 -8596 -4068
rect -7280 -4068 -7184 -4052
rect -8273 -4120 -7551 -4119
rect -8273 -4840 -8272 -4120
rect -7552 -4840 -7551 -4120
rect -8273 -4841 -7551 -4840
rect -8692 -4908 -8596 -4892
rect -7280 -4892 -7264 -4068
rect -7200 -4892 -7184 -4068
rect -5868 -4068 -5772 -4052
rect -6861 -4120 -6139 -4119
rect -6861 -4840 -6860 -4120
rect -6140 -4840 -6139 -4120
rect -6861 -4841 -6139 -4840
rect -7280 -4908 -7184 -4892
rect -5868 -4892 -5852 -4068
rect -5788 -4892 -5772 -4068
rect -4456 -4068 -4360 -4052
rect -5449 -4120 -4727 -4119
rect -5449 -4840 -5448 -4120
rect -4728 -4840 -4727 -4120
rect -5449 -4841 -4727 -4840
rect -5868 -4908 -5772 -4892
rect -4456 -4892 -4440 -4068
rect -4376 -4892 -4360 -4068
rect -3044 -4068 -2948 -4052
rect -4037 -4120 -3315 -4119
rect -4037 -4840 -4036 -4120
rect -3316 -4840 -3315 -4120
rect -4037 -4841 -3315 -4840
rect -4456 -4908 -4360 -4892
rect -3044 -4892 -3028 -4068
rect -2964 -4892 -2948 -4068
rect -1632 -4068 -1536 -4052
rect -2625 -4120 -1903 -4119
rect -2625 -4840 -2624 -4120
rect -1904 -4840 -1903 -4120
rect -2625 -4841 -1903 -4840
rect -3044 -4908 -2948 -4892
rect -1632 -4892 -1616 -4068
rect -1552 -4892 -1536 -4068
rect -220 -4068 -124 -4052
rect -1213 -4120 -491 -4119
rect -1213 -4840 -1212 -4120
rect -492 -4840 -491 -4120
rect -1213 -4841 -491 -4840
rect -1632 -4908 -1536 -4892
rect -220 -4892 -204 -4068
rect -140 -4892 -124 -4068
rect 1192 -4068 1288 -4052
rect 199 -4120 921 -4119
rect 199 -4840 200 -4120
rect 920 -4840 921 -4120
rect 199 -4841 921 -4840
rect -220 -4908 -124 -4892
rect 1192 -4892 1208 -4068
rect 1272 -4892 1288 -4068
rect 2604 -4068 2700 -4052
rect 1611 -4120 2333 -4119
rect 1611 -4840 1612 -4120
rect 2332 -4840 2333 -4120
rect 1611 -4841 2333 -4840
rect 1192 -4908 1288 -4892
rect 2604 -4892 2620 -4068
rect 2684 -4892 2700 -4068
rect 4016 -4068 4112 -4052
rect 3023 -4120 3745 -4119
rect 3023 -4840 3024 -4120
rect 3744 -4840 3745 -4120
rect 3023 -4841 3745 -4840
rect 2604 -4908 2700 -4892
rect 4016 -4892 4032 -4068
rect 4096 -4892 4112 -4068
rect 5428 -4068 5524 -4052
rect 4435 -4120 5157 -4119
rect 4435 -4840 4436 -4120
rect 5156 -4840 5157 -4120
rect 4435 -4841 5157 -4840
rect 4016 -4908 4112 -4892
rect 5428 -4892 5444 -4068
rect 5508 -4892 5524 -4068
rect 6840 -4068 6936 -4052
rect 5847 -4120 6569 -4119
rect 5847 -4840 5848 -4120
rect 6568 -4840 6569 -4120
rect 5847 -4841 6569 -4840
rect 5428 -4908 5524 -4892
rect 6840 -4892 6856 -4068
rect 6920 -4892 6936 -4068
rect 8252 -4068 8348 -4052
rect 7259 -4120 7981 -4119
rect 7259 -4840 7260 -4120
rect 7980 -4840 7981 -4120
rect 7259 -4841 7981 -4840
rect 6840 -4908 6936 -4892
rect 8252 -4892 8268 -4068
rect 8332 -4892 8348 -4068
rect 9664 -4068 9760 -4052
rect 8671 -4120 9393 -4119
rect 8671 -4840 8672 -4120
rect 9392 -4840 9393 -4120
rect 8671 -4841 9393 -4840
rect 8252 -4908 8348 -4892
rect 9664 -4892 9680 -4068
rect 9744 -4892 9760 -4068
rect 11076 -4068 11172 -4052
rect 10083 -4120 10805 -4119
rect 10083 -4840 10084 -4120
rect 10804 -4840 10805 -4120
rect 10083 -4841 10805 -4840
rect 9664 -4908 9760 -4892
rect 11076 -4892 11092 -4068
rect 11156 -4892 11172 -4068
rect 12488 -4068 12584 -4052
rect 11495 -4120 12217 -4119
rect 11495 -4840 11496 -4120
rect 12216 -4840 12217 -4120
rect 11495 -4841 12217 -4840
rect 11076 -4908 11172 -4892
rect 12488 -4892 12504 -4068
rect 12568 -4892 12584 -4068
rect 13900 -4068 13996 -4052
rect 12907 -4120 13629 -4119
rect 12907 -4840 12908 -4120
rect 13628 -4840 13629 -4120
rect 12907 -4841 13629 -4840
rect 12488 -4908 12584 -4892
rect 13900 -4892 13916 -4068
rect 13980 -4892 13996 -4068
rect 15312 -4068 15408 -4052
rect 14319 -4120 15041 -4119
rect 14319 -4840 14320 -4120
rect 15040 -4840 15041 -4120
rect 14319 -4841 15041 -4840
rect 13900 -4908 13996 -4892
rect 15312 -4892 15328 -4068
rect 15392 -4892 15408 -4068
rect 16724 -4068 16820 -4052
rect 15731 -4120 16453 -4119
rect 15731 -4840 15732 -4120
rect 16452 -4840 16453 -4120
rect 15731 -4841 16453 -4840
rect 15312 -4908 15408 -4892
rect 16724 -4892 16740 -4068
rect 16804 -4892 16820 -4068
rect 18136 -4068 18232 -4052
rect 17143 -4120 17865 -4119
rect 17143 -4840 17144 -4120
rect 17864 -4840 17865 -4120
rect 17143 -4841 17865 -4840
rect 16724 -4908 16820 -4892
rect 18136 -4892 18152 -4068
rect 18216 -4892 18232 -4068
rect 19548 -4068 19644 -4052
rect 18555 -4120 19277 -4119
rect 18555 -4840 18556 -4120
rect 19276 -4840 19277 -4120
rect 18555 -4841 19277 -4840
rect 18136 -4908 18232 -4892
rect 19548 -4892 19564 -4068
rect 19628 -4892 19644 -4068
rect 20960 -4068 21056 -4052
rect 19967 -4120 20689 -4119
rect 19967 -4840 19968 -4120
rect 20688 -4840 20689 -4120
rect 19967 -4841 20689 -4840
rect 19548 -4908 19644 -4892
rect 20960 -4892 20976 -4068
rect 21040 -4892 21056 -4068
rect 22372 -4068 22468 -4052
rect 21379 -4120 22101 -4119
rect 21379 -4840 21380 -4120
rect 22100 -4840 22101 -4120
rect 21379 -4841 22101 -4840
rect 20960 -4908 21056 -4892
rect 22372 -4892 22388 -4068
rect 22452 -4892 22468 -4068
rect 23784 -4068 23880 -4052
rect 22791 -4120 23513 -4119
rect 22791 -4840 22792 -4120
rect 23512 -4840 23513 -4120
rect 22791 -4841 23513 -4840
rect 22372 -4908 22468 -4892
rect 23784 -4892 23800 -4068
rect 23864 -4892 23880 -4068
rect 23784 -4908 23880 -4892
rect -22812 -5188 -22716 -5172
rect -23805 -5240 -23083 -5239
rect -23805 -5960 -23804 -5240
rect -23084 -5960 -23083 -5240
rect -23805 -5961 -23083 -5960
rect -22812 -6012 -22796 -5188
rect -22732 -6012 -22716 -5188
rect -21400 -5188 -21304 -5172
rect -22393 -5240 -21671 -5239
rect -22393 -5960 -22392 -5240
rect -21672 -5960 -21671 -5240
rect -22393 -5961 -21671 -5960
rect -22812 -6028 -22716 -6012
rect -21400 -6012 -21384 -5188
rect -21320 -6012 -21304 -5188
rect -19988 -5188 -19892 -5172
rect -20981 -5240 -20259 -5239
rect -20981 -5960 -20980 -5240
rect -20260 -5960 -20259 -5240
rect -20981 -5961 -20259 -5960
rect -21400 -6028 -21304 -6012
rect -19988 -6012 -19972 -5188
rect -19908 -6012 -19892 -5188
rect -18576 -5188 -18480 -5172
rect -19569 -5240 -18847 -5239
rect -19569 -5960 -19568 -5240
rect -18848 -5960 -18847 -5240
rect -19569 -5961 -18847 -5960
rect -19988 -6028 -19892 -6012
rect -18576 -6012 -18560 -5188
rect -18496 -6012 -18480 -5188
rect -17164 -5188 -17068 -5172
rect -18157 -5240 -17435 -5239
rect -18157 -5960 -18156 -5240
rect -17436 -5960 -17435 -5240
rect -18157 -5961 -17435 -5960
rect -18576 -6028 -18480 -6012
rect -17164 -6012 -17148 -5188
rect -17084 -6012 -17068 -5188
rect -15752 -5188 -15656 -5172
rect -16745 -5240 -16023 -5239
rect -16745 -5960 -16744 -5240
rect -16024 -5960 -16023 -5240
rect -16745 -5961 -16023 -5960
rect -17164 -6028 -17068 -6012
rect -15752 -6012 -15736 -5188
rect -15672 -6012 -15656 -5188
rect -14340 -5188 -14244 -5172
rect -15333 -5240 -14611 -5239
rect -15333 -5960 -15332 -5240
rect -14612 -5960 -14611 -5240
rect -15333 -5961 -14611 -5960
rect -15752 -6028 -15656 -6012
rect -14340 -6012 -14324 -5188
rect -14260 -6012 -14244 -5188
rect -12928 -5188 -12832 -5172
rect -13921 -5240 -13199 -5239
rect -13921 -5960 -13920 -5240
rect -13200 -5960 -13199 -5240
rect -13921 -5961 -13199 -5960
rect -14340 -6028 -14244 -6012
rect -12928 -6012 -12912 -5188
rect -12848 -6012 -12832 -5188
rect -11516 -5188 -11420 -5172
rect -12509 -5240 -11787 -5239
rect -12509 -5960 -12508 -5240
rect -11788 -5960 -11787 -5240
rect -12509 -5961 -11787 -5960
rect -12928 -6028 -12832 -6012
rect -11516 -6012 -11500 -5188
rect -11436 -6012 -11420 -5188
rect -10104 -5188 -10008 -5172
rect -11097 -5240 -10375 -5239
rect -11097 -5960 -11096 -5240
rect -10376 -5960 -10375 -5240
rect -11097 -5961 -10375 -5960
rect -11516 -6028 -11420 -6012
rect -10104 -6012 -10088 -5188
rect -10024 -6012 -10008 -5188
rect -8692 -5188 -8596 -5172
rect -9685 -5240 -8963 -5239
rect -9685 -5960 -9684 -5240
rect -8964 -5960 -8963 -5240
rect -9685 -5961 -8963 -5960
rect -10104 -6028 -10008 -6012
rect -8692 -6012 -8676 -5188
rect -8612 -6012 -8596 -5188
rect -7280 -5188 -7184 -5172
rect -8273 -5240 -7551 -5239
rect -8273 -5960 -8272 -5240
rect -7552 -5960 -7551 -5240
rect -8273 -5961 -7551 -5960
rect -8692 -6028 -8596 -6012
rect -7280 -6012 -7264 -5188
rect -7200 -6012 -7184 -5188
rect -5868 -5188 -5772 -5172
rect -6861 -5240 -6139 -5239
rect -6861 -5960 -6860 -5240
rect -6140 -5960 -6139 -5240
rect -6861 -5961 -6139 -5960
rect -7280 -6028 -7184 -6012
rect -5868 -6012 -5852 -5188
rect -5788 -6012 -5772 -5188
rect -4456 -5188 -4360 -5172
rect -5449 -5240 -4727 -5239
rect -5449 -5960 -5448 -5240
rect -4728 -5960 -4727 -5240
rect -5449 -5961 -4727 -5960
rect -5868 -6028 -5772 -6012
rect -4456 -6012 -4440 -5188
rect -4376 -6012 -4360 -5188
rect -3044 -5188 -2948 -5172
rect -4037 -5240 -3315 -5239
rect -4037 -5960 -4036 -5240
rect -3316 -5960 -3315 -5240
rect -4037 -5961 -3315 -5960
rect -4456 -6028 -4360 -6012
rect -3044 -6012 -3028 -5188
rect -2964 -6012 -2948 -5188
rect -1632 -5188 -1536 -5172
rect -2625 -5240 -1903 -5239
rect -2625 -5960 -2624 -5240
rect -1904 -5960 -1903 -5240
rect -2625 -5961 -1903 -5960
rect -3044 -6028 -2948 -6012
rect -1632 -6012 -1616 -5188
rect -1552 -6012 -1536 -5188
rect -220 -5188 -124 -5172
rect -1213 -5240 -491 -5239
rect -1213 -5960 -1212 -5240
rect -492 -5960 -491 -5240
rect -1213 -5961 -491 -5960
rect -1632 -6028 -1536 -6012
rect -220 -6012 -204 -5188
rect -140 -6012 -124 -5188
rect 1192 -5188 1288 -5172
rect 199 -5240 921 -5239
rect 199 -5960 200 -5240
rect 920 -5960 921 -5240
rect 199 -5961 921 -5960
rect -220 -6028 -124 -6012
rect 1192 -6012 1208 -5188
rect 1272 -6012 1288 -5188
rect 2604 -5188 2700 -5172
rect 1611 -5240 2333 -5239
rect 1611 -5960 1612 -5240
rect 2332 -5960 2333 -5240
rect 1611 -5961 2333 -5960
rect 1192 -6028 1288 -6012
rect 2604 -6012 2620 -5188
rect 2684 -6012 2700 -5188
rect 4016 -5188 4112 -5172
rect 3023 -5240 3745 -5239
rect 3023 -5960 3024 -5240
rect 3744 -5960 3745 -5240
rect 3023 -5961 3745 -5960
rect 2604 -6028 2700 -6012
rect 4016 -6012 4032 -5188
rect 4096 -6012 4112 -5188
rect 5428 -5188 5524 -5172
rect 4435 -5240 5157 -5239
rect 4435 -5960 4436 -5240
rect 5156 -5960 5157 -5240
rect 4435 -5961 5157 -5960
rect 4016 -6028 4112 -6012
rect 5428 -6012 5444 -5188
rect 5508 -6012 5524 -5188
rect 6840 -5188 6936 -5172
rect 5847 -5240 6569 -5239
rect 5847 -5960 5848 -5240
rect 6568 -5960 6569 -5240
rect 5847 -5961 6569 -5960
rect 5428 -6028 5524 -6012
rect 6840 -6012 6856 -5188
rect 6920 -6012 6936 -5188
rect 8252 -5188 8348 -5172
rect 7259 -5240 7981 -5239
rect 7259 -5960 7260 -5240
rect 7980 -5960 7981 -5240
rect 7259 -5961 7981 -5960
rect 6840 -6028 6936 -6012
rect 8252 -6012 8268 -5188
rect 8332 -6012 8348 -5188
rect 9664 -5188 9760 -5172
rect 8671 -5240 9393 -5239
rect 8671 -5960 8672 -5240
rect 9392 -5960 9393 -5240
rect 8671 -5961 9393 -5960
rect 8252 -6028 8348 -6012
rect 9664 -6012 9680 -5188
rect 9744 -6012 9760 -5188
rect 11076 -5188 11172 -5172
rect 10083 -5240 10805 -5239
rect 10083 -5960 10084 -5240
rect 10804 -5960 10805 -5240
rect 10083 -5961 10805 -5960
rect 9664 -6028 9760 -6012
rect 11076 -6012 11092 -5188
rect 11156 -6012 11172 -5188
rect 12488 -5188 12584 -5172
rect 11495 -5240 12217 -5239
rect 11495 -5960 11496 -5240
rect 12216 -5960 12217 -5240
rect 11495 -5961 12217 -5960
rect 11076 -6028 11172 -6012
rect 12488 -6012 12504 -5188
rect 12568 -6012 12584 -5188
rect 13900 -5188 13996 -5172
rect 12907 -5240 13629 -5239
rect 12907 -5960 12908 -5240
rect 13628 -5960 13629 -5240
rect 12907 -5961 13629 -5960
rect 12488 -6028 12584 -6012
rect 13900 -6012 13916 -5188
rect 13980 -6012 13996 -5188
rect 15312 -5188 15408 -5172
rect 14319 -5240 15041 -5239
rect 14319 -5960 14320 -5240
rect 15040 -5960 15041 -5240
rect 14319 -5961 15041 -5960
rect 13900 -6028 13996 -6012
rect 15312 -6012 15328 -5188
rect 15392 -6012 15408 -5188
rect 16724 -5188 16820 -5172
rect 15731 -5240 16453 -5239
rect 15731 -5960 15732 -5240
rect 16452 -5960 16453 -5240
rect 15731 -5961 16453 -5960
rect 15312 -6028 15408 -6012
rect 16724 -6012 16740 -5188
rect 16804 -6012 16820 -5188
rect 18136 -5188 18232 -5172
rect 17143 -5240 17865 -5239
rect 17143 -5960 17144 -5240
rect 17864 -5960 17865 -5240
rect 17143 -5961 17865 -5960
rect 16724 -6028 16820 -6012
rect 18136 -6012 18152 -5188
rect 18216 -6012 18232 -5188
rect 19548 -5188 19644 -5172
rect 18555 -5240 19277 -5239
rect 18555 -5960 18556 -5240
rect 19276 -5960 19277 -5240
rect 18555 -5961 19277 -5960
rect 18136 -6028 18232 -6012
rect 19548 -6012 19564 -5188
rect 19628 -6012 19644 -5188
rect 20960 -5188 21056 -5172
rect 19967 -5240 20689 -5239
rect 19967 -5960 19968 -5240
rect 20688 -5960 20689 -5240
rect 19967 -5961 20689 -5960
rect 19548 -6028 19644 -6012
rect 20960 -6012 20976 -5188
rect 21040 -6012 21056 -5188
rect 22372 -5188 22468 -5172
rect 21379 -5240 22101 -5239
rect 21379 -5960 21380 -5240
rect 22100 -5960 22101 -5240
rect 21379 -5961 22101 -5960
rect 20960 -6028 21056 -6012
rect 22372 -6012 22388 -5188
rect 22452 -6012 22468 -5188
rect 23784 -5188 23880 -5172
rect 22791 -5240 23513 -5239
rect 22791 -5960 22792 -5240
rect 23512 -5960 23513 -5240
rect 22791 -5961 23513 -5960
rect 22372 -6028 22468 -6012
rect 23784 -6012 23800 -5188
rect 23864 -6012 23880 -5188
rect 23784 -6028 23880 -6012
rect -22812 -6308 -22716 -6292
rect -23805 -6360 -23083 -6359
rect -23805 -7080 -23804 -6360
rect -23084 -7080 -23083 -6360
rect -23805 -7081 -23083 -7080
rect -22812 -7132 -22796 -6308
rect -22732 -7132 -22716 -6308
rect -21400 -6308 -21304 -6292
rect -22393 -6360 -21671 -6359
rect -22393 -7080 -22392 -6360
rect -21672 -7080 -21671 -6360
rect -22393 -7081 -21671 -7080
rect -22812 -7148 -22716 -7132
rect -21400 -7132 -21384 -6308
rect -21320 -7132 -21304 -6308
rect -19988 -6308 -19892 -6292
rect -20981 -6360 -20259 -6359
rect -20981 -7080 -20980 -6360
rect -20260 -7080 -20259 -6360
rect -20981 -7081 -20259 -7080
rect -21400 -7148 -21304 -7132
rect -19988 -7132 -19972 -6308
rect -19908 -7132 -19892 -6308
rect -18576 -6308 -18480 -6292
rect -19569 -6360 -18847 -6359
rect -19569 -7080 -19568 -6360
rect -18848 -7080 -18847 -6360
rect -19569 -7081 -18847 -7080
rect -19988 -7148 -19892 -7132
rect -18576 -7132 -18560 -6308
rect -18496 -7132 -18480 -6308
rect -17164 -6308 -17068 -6292
rect -18157 -6360 -17435 -6359
rect -18157 -7080 -18156 -6360
rect -17436 -7080 -17435 -6360
rect -18157 -7081 -17435 -7080
rect -18576 -7148 -18480 -7132
rect -17164 -7132 -17148 -6308
rect -17084 -7132 -17068 -6308
rect -15752 -6308 -15656 -6292
rect -16745 -6360 -16023 -6359
rect -16745 -7080 -16744 -6360
rect -16024 -7080 -16023 -6360
rect -16745 -7081 -16023 -7080
rect -17164 -7148 -17068 -7132
rect -15752 -7132 -15736 -6308
rect -15672 -7132 -15656 -6308
rect -14340 -6308 -14244 -6292
rect -15333 -6360 -14611 -6359
rect -15333 -7080 -15332 -6360
rect -14612 -7080 -14611 -6360
rect -15333 -7081 -14611 -7080
rect -15752 -7148 -15656 -7132
rect -14340 -7132 -14324 -6308
rect -14260 -7132 -14244 -6308
rect -12928 -6308 -12832 -6292
rect -13921 -6360 -13199 -6359
rect -13921 -7080 -13920 -6360
rect -13200 -7080 -13199 -6360
rect -13921 -7081 -13199 -7080
rect -14340 -7148 -14244 -7132
rect -12928 -7132 -12912 -6308
rect -12848 -7132 -12832 -6308
rect -11516 -6308 -11420 -6292
rect -12509 -6360 -11787 -6359
rect -12509 -7080 -12508 -6360
rect -11788 -7080 -11787 -6360
rect -12509 -7081 -11787 -7080
rect -12928 -7148 -12832 -7132
rect -11516 -7132 -11500 -6308
rect -11436 -7132 -11420 -6308
rect -10104 -6308 -10008 -6292
rect -11097 -6360 -10375 -6359
rect -11097 -7080 -11096 -6360
rect -10376 -7080 -10375 -6360
rect -11097 -7081 -10375 -7080
rect -11516 -7148 -11420 -7132
rect -10104 -7132 -10088 -6308
rect -10024 -7132 -10008 -6308
rect -8692 -6308 -8596 -6292
rect -9685 -6360 -8963 -6359
rect -9685 -7080 -9684 -6360
rect -8964 -7080 -8963 -6360
rect -9685 -7081 -8963 -7080
rect -10104 -7148 -10008 -7132
rect -8692 -7132 -8676 -6308
rect -8612 -7132 -8596 -6308
rect -7280 -6308 -7184 -6292
rect -8273 -6360 -7551 -6359
rect -8273 -7080 -8272 -6360
rect -7552 -7080 -7551 -6360
rect -8273 -7081 -7551 -7080
rect -8692 -7148 -8596 -7132
rect -7280 -7132 -7264 -6308
rect -7200 -7132 -7184 -6308
rect -5868 -6308 -5772 -6292
rect -6861 -6360 -6139 -6359
rect -6861 -7080 -6860 -6360
rect -6140 -7080 -6139 -6360
rect -6861 -7081 -6139 -7080
rect -7280 -7148 -7184 -7132
rect -5868 -7132 -5852 -6308
rect -5788 -7132 -5772 -6308
rect -4456 -6308 -4360 -6292
rect -5449 -6360 -4727 -6359
rect -5449 -7080 -5448 -6360
rect -4728 -7080 -4727 -6360
rect -5449 -7081 -4727 -7080
rect -5868 -7148 -5772 -7132
rect -4456 -7132 -4440 -6308
rect -4376 -7132 -4360 -6308
rect -3044 -6308 -2948 -6292
rect -4037 -6360 -3315 -6359
rect -4037 -7080 -4036 -6360
rect -3316 -7080 -3315 -6360
rect -4037 -7081 -3315 -7080
rect -4456 -7148 -4360 -7132
rect -3044 -7132 -3028 -6308
rect -2964 -7132 -2948 -6308
rect -1632 -6308 -1536 -6292
rect -2625 -6360 -1903 -6359
rect -2625 -7080 -2624 -6360
rect -1904 -7080 -1903 -6360
rect -2625 -7081 -1903 -7080
rect -3044 -7148 -2948 -7132
rect -1632 -7132 -1616 -6308
rect -1552 -7132 -1536 -6308
rect -220 -6308 -124 -6292
rect -1213 -6360 -491 -6359
rect -1213 -7080 -1212 -6360
rect -492 -7080 -491 -6360
rect -1213 -7081 -491 -7080
rect -1632 -7148 -1536 -7132
rect -220 -7132 -204 -6308
rect -140 -7132 -124 -6308
rect 1192 -6308 1288 -6292
rect 199 -6360 921 -6359
rect 199 -7080 200 -6360
rect 920 -7080 921 -6360
rect 199 -7081 921 -7080
rect -220 -7148 -124 -7132
rect 1192 -7132 1208 -6308
rect 1272 -7132 1288 -6308
rect 2604 -6308 2700 -6292
rect 1611 -6360 2333 -6359
rect 1611 -7080 1612 -6360
rect 2332 -7080 2333 -6360
rect 1611 -7081 2333 -7080
rect 1192 -7148 1288 -7132
rect 2604 -7132 2620 -6308
rect 2684 -7132 2700 -6308
rect 4016 -6308 4112 -6292
rect 3023 -6360 3745 -6359
rect 3023 -7080 3024 -6360
rect 3744 -7080 3745 -6360
rect 3023 -7081 3745 -7080
rect 2604 -7148 2700 -7132
rect 4016 -7132 4032 -6308
rect 4096 -7132 4112 -6308
rect 5428 -6308 5524 -6292
rect 4435 -6360 5157 -6359
rect 4435 -7080 4436 -6360
rect 5156 -7080 5157 -6360
rect 4435 -7081 5157 -7080
rect 4016 -7148 4112 -7132
rect 5428 -7132 5444 -6308
rect 5508 -7132 5524 -6308
rect 6840 -6308 6936 -6292
rect 5847 -6360 6569 -6359
rect 5847 -7080 5848 -6360
rect 6568 -7080 6569 -6360
rect 5847 -7081 6569 -7080
rect 5428 -7148 5524 -7132
rect 6840 -7132 6856 -6308
rect 6920 -7132 6936 -6308
rect 8252 -6308 8348 -6292
rect 7259 -6360 7981 -6359
rect 7259 -7080 7260 -6360
rect 7980 -7080 7981 -6360
rect 7259 -7081 7981 -7080
rect 6840 -7148 6936 -7132
rect 8252 -7132 8268 -6308
rect 8332 -7132 8348 -6308
rect 9664 -6308 9760 -6292
rect 8671 -6360 9393 -6359
rect 8671 -7080 8672 -6360
rect 9392 -7080 9393 -6360
rect 8671 -7081 9393 -7080
rect 8252 -7148 8348 -7132
rect 9664 -7132 9680 -6308
rect 9744 -7132 9760 -6308
rect 11076 -6308 11172 -6292
rect 10083 -6360 10805 -6359
rect 10083 -7080 10084 -6360
rect 10804 -7080 10805 -6360
rect 10083 -7081 10805 -7080
rect 9664 -7148 9760 -7132
rect 11076 -7132 11092 -6308
rect 11156 -7132 11172 -6308
rect 12488 -6308 12584 -6292
rect 11495 -6360 12217 -6359
rect 11495 -7080 11496 -6360
rect 12216 -7080 12217 -6360
rect 11495 -7081 12217 -7080
rect 11076 -7148 11172 -7132
rect 12488 -7132 12504 -6308
rect 12568 -7132 12584 -6308
rect 13900 -6308 13996 -6292
rect 12907 -6360 13629 -6359
rect 12907 -7080 12908 -6360
rect 13628 -7080 13629 -6360
rect 12907 -7081 13629 -7080
rect 12488 -7148 12584 -7132
rect 13900 -7132 13916 -6308
rect 13980 -7132 13996 -6308
rect 15312 -6308 15408 -6292
rect 14319 -6360 15041 -6359
rect 14319 -7080 14320 -6360
rect 15040 -7080 15041 -6360
rect 14319 -7081 15041 -7080
rect 13900 -7148 13996 -7132
rect 15312 -7132 15328 -6308
rect 15392 -7132 15408 -6308
rect 16724 -6308 16820 -6292
rect 15731 -6360 16453 -6359
rect 15731 -7080 15732 -6360
rect 16452 -7080 16453 -6360
rect 15731 -7081 16453 -7080
rect 15312 -7148 15408 -7132
rect 16724 -7132 16740 -6308
rect 16804 -7132 16820 -6308
rect 18136 -6308 18232 -6292
rect 17143 -6360 17865 -6359
rect 17143 -7080 17144 -6360
rect 17864 -7080 17865 -6360
rect 17143 -7081 17865 -7080
rect 16724 -7148 16820 -7132
rect 18136 -7132 18152 -6308
rect 18216 -7132 18232 -6308
rect 19548 -6308 19644 -6292
rect 18555 -6360 19277 -6359
rect 18555 -7080 18556 -6360
rect 19276 -7080 19277 -6360
rect 18555 -7081 19277 -7080
rect 18136 -7148 18232 -7132
rect 19548 -7132 19564 -6308
rect 19628 -7132 19644 -6308
rect 20960 -6308 21056 -6292
rect 19967 -6360 20689 -6359
rect 19967 -7080 19968 -6360
rect 20688 -7080 20689 -6360
rect 19967 -7081 20689 -7080
rect 19548 -7148 19644 -7132
rect 20960 -7132 20976 -6308
rect 21040 -7132 21056 -6308
rect 22372 -6308 22468 -6292
rect 21379 -6360 22101 -6359
rect 21379 -7080 21380 -6360
rect 22100 -7080 22101 -6360
rect 21379 -7081 22101 -7080
rect 20960 -7148 21056 -7132
rect 22372 -7132 22388 -6308
rect 22452 -7132 22468 -6308
rect 23784 -6308 23880 -6292
rect 22791 -6360 23513 -6359
rect 22791 -7080 22792 -6360
rect 23512 -7080 23513 -6360
rect 22791 -7081 23513 -7080
rect 22372 -7148 22468 -7132
rect 23784 -7132 23800 -6308
rect 23864 -7132 23880 -6308
rect 23784 -7148 23880 -7132
rect -22812 -7428 -22716 -7412
rect -23805 -7480 -23083 -7479
rect -23805 -8200 -23804 -7480
rect -23084 -8200 -23083 -7480
rect -23805 -8201 -23083 -8200
rect -22812 -8252 -22796 -7428
rect -22732 -8252 -22716 -7428
rect -21400 -7428 -21304 -7412
rect -22393 -7480 -21671 -7479
rect -22393 -8200 -22392 -7480
rect -21672 -8200 -21671 -7480
rect -22393 -8201 -21671 -8200
rect -22812 -8268 -22716 -8252
rect -21400 -8252 -21384 -7428
rect -21320 -8252 -21304 -7428
rect -19988 -7428 -19892 -7412
rect -20981 -7480 -20259 -7479
rect -20981 -8200 -20980 -7480
rect -20260 -8200 -20259 -7480
rect -20981 -8201 -20259 -8200
rect -21400 -8268 -21304 -8252
rect -19988 -8252 -19972 -7428
rect -19908 -8252 -19892 -7428
rect -18576 -7428 -18480 -7412
rect -19569 -7480 -18847 -7479
rect -19569 -8200 -19568 -7480
rect -18848 -8200 -18847 -7480
rect -19569 -8201 -18847 -8200
rect -19988 -8268 -19892 -8252
rect -18576 -8252 -18560 -7428
rect -18496 -8252 -18480 -7428
rect -17164 -7428 -17068 -7412
rect -18157 -7480 -17435 -7479
rect -18157 -8200 -18156 -7480
rect -17436 -8200 -17435 -7480
rect -18157 -8201 -17435 -8200
rect -18576 -8268 -18480 -8252
rect -17164 -8252 -17148 -7428
rect -17084 -8252 -17068 -7428
rect -15752 -7428 -15656 -7412
rect -16745 -7480 -16023 -7479
rect -16745 -8200 -16744 -7480
rect -16024 -8200 -16023 -7480
rect -16745 -8201 -16023 -8200
rect -17164 -8268 -17068 -8252
rect -15752 -8252 -15736 -7428
rect -15672 -8252 -15656 -7428
rect -14340 -7428 -14244 -7412
rect -15333 -7480 -14611 -7479
rect -15333 -8200 -15332 -7480
rect -14612 -8200 -14611 -7480
rect -15333 -8201 -14611 -8200
rect -15752 -8268 -15656 -8252
rect -14340 -8252 -14324 -7428
rect -14260 -8252 -14244 -7428
rect -12928 -7428 -12832 -7412
rect -13921 -7480 -13199 -7479
rect -13921 -8200 -13920 -7480
rect -13200 -8200 -13199 -7480
rect -13921 -8201 -13199 -8200
rect -14340 -8268 -14244 -8252
rect -12928 -8252 -12912 -7428
rect -12848 -8252 -12832 -7428
rect -11516 -7428 -11420 -7412
rect -12509 -7480 -11787 -7479
rect -12509 -8200 -12508 -7480
rect -11788 -8200 -11787 -7480
rect -12509 -8201 -11787 -8200
rect -12928 -8268 -12832 -8252
rect -11516 -8252 -11500 -7428
rect -11436 -8252 -11420 -7428
rect -10104 -7428 -10008 -7412
rect -11097 -7480 -10375 -7479
rect -11097 -8200 -11096 -7480
rect -10376 -8200 -10375 -7480
rect -11097 -8201 -10375 -8200
rect -11516 -8268 -11420 -8252
rect -10104 -8252 -10088 -7428
rect -10024 -8252 -10008 -7428
rect -8692 -7428 -8596 -7412
rect -9685 -7480 -8963 -7479
rect -9685 -8200 -9684 -7480
rect -8964 -8200 -8963 -7480
rect -9685 -8201 -8963 -8200
rect -10104 -8268 -10008 -8252
rect -8692 -8252 -8676 -7428
rect -8612 -8252 -8596 -7428
rect -7280 -7428 -7184 -7412
rect -8273 -7480 -7551 -7479
rect -8273 -8200 -8272 -7480
rect -7552 -8200 -7551 -7480
rect -8273 -8201 -7551 -8200
rect -8692 -8268 -8596 -8252
rect -7280 -8252 -7264 -7428
rect -7200 -8252 -7184 -7428
rect -5868 -7428 -5772 -7412
rect -6861 -7480 -6139 -7479
rect -6861 -8200 -6860 -7480
rect -6140 -8200 -6139 -7480
rect -6861 -8201 -6139 -8200
rect -7280 -8268 -7184 -8252
rect -5868 -8252 -5852 -7428
rect -5788 -8252 -5772 -7428
rect -4456 -7428 -4360 -7412
rect -5449 -7480 -4727 -7479
rect -5449 -8200 -5448 -7480
rect -4728 -8200 -4727 -7480
rect -5449 -8201 -4727 -8200
rect -5868 -8268 -5772 -8252
rect -4456 -8252 -4440 -7428
rect -4376 -8252 -4360 -7428
rect -3044 -7428 -2948 -7412
rect -4037 -7480 -3315 -7479
rect -4037 -8200 -4036 -7480
rect -3316 -8200 -3315 -7480
rect -4037 -8201 -3315 -8200
rect -4456 -8268 -4360 -8252
rect -3044 -8252 -3028 -7428
rect -2964 -8252 -2948 -7428
rect -1632 -7428 -1536 -7412
rect -2625 -7480 -1903 -7479
rect -2625 -8200 -2624 -7480
rect -1904 -8200 -1903 -7480
rect -2625 -8201 -1903 -8200
rect -3044 -8268 -2948 -8252
rect -1632 -8252 -1616 -7428
rect -1552 -8252 -1536 -7428
rect -220 -7428 -124 -7412
rect -1213 -7480 -491 -7479
rect -1213 -8200 -1212 -7480
rect -492 -8200 -491 -7480
rect -1213 -8201 -491 -8200
rect -1632 -8268 -1536 -8252
rect -220 -8252 -204 -7428
rect -140 -8252 -124 -7428
rect 1192 -7428 1288 -7412
rect 199 -7480 921 -7479
rect 199 -8200 200 -7480
rect 920 -8200 921 -7480
rect 199 -8201 921 -8200
rect -220 -8268 -124 -8252
rect 1192 -8252 1208 -7428
rect 1272 -8252 1288 -7428
rect 2604 -7428 2700 -7412
rect 1611 -7480 2333 -7479
rect 1611 -8200 1612 -7480
rect 2332 -8200 2333 -7480
rect 1611 -8201 2333 -8200
rect 1192 -8268 1288 -8252
rect 2604 -8252 2620 -7428
rect 2684 -8252 2700 -7428
rect 4016 -7428 4112 -7412
rect 3023 -7480 3745 -7479
rect 3023 -8200 3024 -7480
rect 3744 -8200 3745 -7480
rect 3023 -8201 3745 -8200
rect 2604 -8268 2700 -8252
rect 4016 -8252 4032 -7428
rect 4096 -8252 4112 -7428
rect 5428 -7428 5524 -7412
rect 4435 -7480 5157 -7479
rect 4435 -8200 4436 -7480
rect 5156 -8200 5157 -7480
rect 4435 -8201 5157 -8200
rect 4016 -8268 4112 -8252
rect 5428 -8252 5444 -7428
rect 5508 -8252 5524 -7428
rect 6840 -7428 6936 -7412
rect 5847 -7480 6569 -7479
rect 5847 -8200 5848 -7480
rect 6568 -8200 6569 -7480
rect 5847 -8201 6569 -8200
rect 5428 -8268 5524 -8252
rect 6840 -8252 6856 -7428
rect 6920 -8252 6936 -7428
rect 8252 -7428 8348 -7412
rect 7259 -7480 7981 -7479
rect 7259 -8200 7260 -7480
rect 7980 -8200 7981 -7480
rect 7259 -8201 7981 -8200
rect 6840 -8268 6936 -8252
rect 8252 -8252 8268 -7428
rect 8332 -8252 8348 -7428
rect 9664 -7428 9760 -7412
rect 8671 -7480 9393 -7479
rect 8671 -8200 8672 -7480
rect 9392 -8200 9393 -7480
rect 8671 -8201 9393 -8200
rect 8252 -8268 8348 -8252
rect 9664 -8252 9680 -7428
rect 9744 -8252 9760 -7428
rect 11076 -7428 11172 -7412
rect 10083 -7480 10805 -7479
rect 10083 -8200 10084 -7480
rect 10804 -8200 10805 -7480
rect 10083 -8201 10805 -8200
rect 9664 -8268 9760 -8252
rect 11076 -8252 11092 -7428
rect 11156 -8252 11172 -7428
rect 12488 -7428 12584 -7412
rect 11495 -7480 12217 -7479
rect 11495 -8200 11496 -7480
rect 12216 -8200 12217 -7480
rect 11495 -8201 12217 -8200
rect 11076 -8268 11172 -8252
rect 12488 -8252 12504 -7428
rect 12568 -8252 12584 -7428
rect 13900 -7428 13996 -7412
rect 12907 -7480 13629 -7479
rect 12907 -8200 12908 -7480
rect 13628 -8200 13629 -7480
rect 12907 -8201 13629 -8200
rect 12488 -8268 12584 -8252
rect 13900 -8252 13916 -7428
rect 13980 -8252 13996 -7428
rect 15312 -7428 15408 -7412
rect 14319 -7480 15041 -7479
rect 14319 -8200 14320 -7480
rect 15040 -8200 15041 -7480
rect 14319 -8201 15041 -8200
rect 13900 -8268 13996 -8252
rect 15312 -8252 15328 -7428
rect 15392 -8252 15408 -7428
rect 16724 -7428 16820 -7412
rect 15731 -7480 16453 -7479
rect 15731 -8200 15732 -7480
rect 16452 -8200 16453 -7480
rect 15731 -8201 16453 -8200
rect 15312 -8268 15408 -8252
rect 16724 -8252 16740 -7428
rect 16804 -8252 16820 -7428
rect 18136 -7428 18232 -7412
rect 17143 -7480 17865 -7479
rect 17143 -8200 17144 -7480
rect 17864 -8200 17865 -7480
rect 17143 -8201 17865 -8200
rect 16724 -8268 16820 -8252
rect 18136 -8252 18152 -7428
rect 18216 -8252 18232 -7428
rect 19548 -7428 19644 -7412
rect 18555 -7480 19277 -7479
rect 18555 -8200 18556 -7480
rect 19276 -8200 19277 -7480
rect 18555 -8201 19277 -8200
rect 18136 -8268 18232 -8252
rect 19548 -8252 19564 -7428
rect 19628 -8252 19644 -7428
rect 20960 -7428 21056 -7412
rect 19967 -7480 20689 -7479
rect 19967 -8200 19968 -7480
rect 20688 -8200 20689 -7480
rect 19967 -8201 20689 -8200
rect 19548 -8268 19644 -8252
rect 20960 -8252 20976 -7428
rect 21040 -8252 21056 -7428
rect 22372 -7428 22468 -7412
rect 21379 -7480 22101 -7479
rect 21379 -8200 21380 -7480
rect 22100 -8200 22101 -7480
rect 21379 -8201 22101 -8200
rect 20960 -8268 21056 -8252
rect 22372 -8252 22388 -7428
rect 22452 -8252 22468 -7428
rect 23784 -7428 23880 -7412
rect 22791 -7480 23513 -7479
rect 22791 -8200 22792 -7480
rect 23512 -8200 23513 -7480
rect 22791 -8201 23513 -8200
rect 22372 -8268 22468 -8252
rect 23784 -8252 23800 -7428
rect 23864 -8252 23880 -7428
rect 23784 -8268 23880 -8252
rect -22812 -8548 -22716 -8532
rect -23805 -8600 -23083 -8599
rect -23805 -9320 -23804 -8600
rect -23084 -9320 -23083 -8600
rect -23805 -9321 -23083 -9320
rect -22812 -9372 -22796 -8548
rect -22732 -9372 -22716 -8548
rect -21400 -8548 -21304 -8532
rect -22393 -8600 -21671 -8599
rect -22393 -9320 -22392 -8600
rect -21672 -9320 -21671 -8600
rect -22393 -9321 -21671 -9320
rect -22812 -9388 -22716 -9372
rect -21400 -9372 -21384 -8548
rect -21320 -9372 -21304 -8548
rect -19988 -8548 -19892 -8532
rect -20981 -8600 -20259 -8599
rect -20981 -9320 -20980 -8600
rect -20260 -9320 -20259 -8600
rect -20981 -9321 -20259 -9320
rect -21400 -9388 -21304 -9372
rect -19988 -9372 -19972 -8548
rect -19908 -9372 -19892 -8548
rect -18576 -8548 -18480 -8532
rect -19569 -8600 -18847 -8599
rect -19569 -9320 -19568 -8600
rect -18848 -9320 -18847 -8600
rect -19569 -9321 -18847 -9320
rect -19988 -9388 -19892 -9372
rect -18576 -9372 -18560 -8548
rect -18496 -9372 -18480 -8548
rect -17164 -8548 -17068 -8532
rect -18157 -8600 -17435 -8599
rect -18157 -9320 -18156 -8600
rect -17436 -9320 -17435 -8600
rect -18157 -9321 -17435 -9320
rect -18576 -9388 -18480 -9372
rect -17164 -9372 -17148 -8548
rect -17084 -9372 -17068 -8548
rect -15752 -8548 -15656 -8532
rect -16745 -8600 -16023 -8599
rect -16745 -9320 -16744 -8600
rect -16024 -9320 -16023 -8600
rect -16745 -9321 -16023 -9320
rect -17164 -9388 -17068 -9372
rect -15752 -9372 -15736 -8548
rect -15672 -9372 -15656 -8548
rect -14340 -8548 -14244 -8532
rect -15333 -8600 -14611 -8599
rect -15333 -9320 -15332 -8600
rect -14612 -9320 -14611 -8600
rect -15333 -9321 -14611 -9320
rect -15752 -9388 -15656 -9372
rect -14340 -9372 -14324 -8548
rect -14260 -9372 -14244 -8548
rect -12928 -8548 -12832 -8532
rect -13921 -8600 -13199 -8599
rect -13921 -9320 -13920 -8600
rect -13200 -9320 -13199 -8600
rect -13921 -9321 -13199 -9320
rect -14340 -9388 -14244 -9372
rect -12928 -9372 -12912 -8548
rect -12848 -9372 -12832 -8548
rect -11516 -8548 -11420 -8532
rect -12509 -8600 -11787 -8599
rect -12509 -9320 -12508 -8600
rect -11788 -9320 -11787 -8600
rect -12509 -9321 -11787 -9320
rect -12928 -9388 -12832 -9372
rect -11516 -9372 -11500 -8548
rect -11436 -9372 -11420 -8548
rect -10104 -8548 -10008 -8532
rect -11097 -8600 -10375 -8599
rect -11097 -9320 -11096 -8600
rect -10376 -9320 -10375 -8600
rect -11097 -9321 -10375 -9320
rect -11516 -9388 -11420 -9372
rect -10104 -9372 -10088 -8548
rect -10024 -9372 -10008 -8548
rect -8692 -8548 -8596 -8532
rect -9685 -8600 -8963 -8599
rect -9685 -9320 -9684 -8600
rect -8964 -9320 -8963 -8600
rect -9685 -9321 -8963 -9320
rect -10104 -9388 -10008 -9372
rect -8692 -9372 -8676 -8548
rect -8612 -9372 -8596 -8548
rect -7280 -8548 -7184 -8532
rect -8273 -8600 -7551 -8599
rect -8273 -9320 -8272 -8600
rect -7552 -9320 -7551 -8600
rect -8273 -9321 -7551 -9320
rect -8692 -9388 -8596 -9372
rect -7280 -9372 -7264 -8548
rect -7200 -9372 -7184 -8548
rect -5868 -8548 -5772 -8532
rect -6861 -8600 -6139 -8599
rect -6861 -9320 -6860 -8600
rect -6140 -9320 -6139 -8600
rect -6861 -9321 -6139 -9320
rect -7280 -9388 -7184 -9372
rect -5868 -9372 -5852 -8548
rect -5788 -9372 -5772 -8548
rect -4456 -8548 -4360 -8532
rect -5449 -8600 -4727 -8599
rect -5449 -9320 -5448 -8600
rect -4728 -9320 -4727 -8600
rect -5449 -9321 -4727 -9320
rect -5868 -9388 -5772 -9372
rect -4456 -9372 -4440 -8548
rect -4376 -9372 -4360 -8548
rect -3044 -8548 -2948 -8532
rect -4037 -8600 -3315 -8599
rect -4037 -9320 -4036 -8600
rect -3316 -9320 -3315 -8600
rect -4037 -9321 -3315 -9320
rect -4456 -9388 -4360 -9372
rect -3044 -9372 -3028 -8548
rect -2964 -9372 -2948 -8548
rect -1632 -8548 -1536 -8532
rect -2625 -8600 -1903 -8599
rect -2625 -9320 -2624 -8600
rect -1904 -9320 -1903 -8600
rect -2625 -9321 -1903 -9320
rect -3044 -9388 -2948 -9372
rect -1632 -9372 -1616 -8548
rect -1552 -9372 -1536 -8548
rect -220 -8548 -124 -8532
rect -1213 -8600 -491 -8599
rect -1213 -9320 -1212 -8600
rect -492 -9320 -491 -8600
rect -1213 -9321 -491 -9320
rect -1632 -9388 -1536 -9372
rect -220 -9372 -204 -8548
rect -140 -9372 -124 -8548
rect 1192 -8548 1288 -8532
rect 199 -8600 921 -8599
rect 199 -9320 200 -8600
rect 920 -9320 921 -8600
rect 199 -9321 921 -9320
rect -220 -9388 -124 -9372
rect 1192 -9372 1208 -8548
rect 1272 -9372 1288 -8548
rect 2604 -8548 2700 -8532
rect 1611 -8600 2333 -8599
rect 1611 -9320 1612 -8600
rect 2332 -9320 2333 -8600
rect 1611 -9321 2333 -9320
rect 1192 -9388 1288 -9372
rect 2604 -9372 2620 -8548
rect 2684 -9372 2700 -8548
rect 4016 -8548 4112 -8532
rect 3023 -8600 3745 -8599
rect 3023 -9320 3024 -8600
rect 3744 -9320 3745 -8600
rect 3023 -9321 3745 -9320
rect 2604 -9388 2700 -9372
rect 4016 -9372 4032 -8548
rect 4096 -9372 4112 -8548
rect 5428 -8548 5524 -8532
rect 4435 -8600 5157 -8599
rect 4435 -9320 4436 -8600
rect 5156 -9320 5157 -8600
rect 4435 -9321 5157 -9320
rect 4016 -9388 4112 -9372
rect 5428 -9372 5444 -8548
rect 5508 -9372 5524 -8548
rect 6840 -8548 6936 -8532
rect 5847 -8600 6569 -8599
rect 5847 -9320 5848 -8600
rect 6568 -9320 6569 -8600
rect 5847 -9321 6569 -9320
rect 5428 -9388 5524 -9372
rect 6840 -9372 6856 -8548
rect 6920 -9372 6936 -8548
rect 8252 -8548 8348 -8532
rect 7259 -8600 7981 -8599
rect 7259 -9320 7260 -8600
rect 7980 -9320 7981 -8600
rect 7259 -9321 7981 -9320
rect 6840 -9388 6936 -9372
rect 8252 -9372 8268 -8548
rect 8332 -9372 8348 -8548
rect 9664 -8548 9760 -8532
rect 8671 -8600 9393 -8599
rect 8671 -9320 8672 -8600
rect 9392 -9320 9393 -8600
rect 8671 -9321 9393 -9320
rect 8252 -9388 8348 -9372
rect 9664 -9372 9680 -8548
rect 9744 -9372 9760 -8548
rect 11076 -8548 11172 -8532
rect 10083 -8600 10805 -8599
rect 10083 -9320 10084 -8600
rect 10804 -9320 10805 -8600
rect 10083 -9321 10805 -9320
rect 9664 -9388 9760 -9372
rect 11076 -9372 11092 -8548
rect 11156 -9372 11172 -8548
rect 12488 -8548 12584 -8532
rect 11495 -8600 12217 -8599
rect 11495 -9320 11496 -8600
rect 12216 -9320 12217 -8600
rect 11495 -9321 12217 -9320
rect 11076 -9388 11172 -9372
rect 12488 -9372 12504 -8548
rect 12568 -9372 12584 -8548
rect 13900 -8548 13996 -8532
rect 12907 -8600 13629 -8599
rect 12907 -9320 12908 -8600
rect 13628 -9320 13629 -8600
rect 12907 -9321 13629 -9320
rect 12488 -9388 12584 -9372
rect 13900 -9372 13916 -8548
rect 13980 -9372 13996 -8548
rect 15312 -8548 15408 -8532
rect 14319 -8600 15041 -8599
rect 14319 -9320 14320 -8600
rect 15040 -9320 15041 -8600
rect 14319 -9321 15041 -9320
rect 13900 -9388 13996 -9372
rect 15312 -9372 15328 -8548
rect 15392 -9372 15408 -8548
rect 16724 -8548 16820 -8532
rect 15731 -8600 16453 -8599
rect 15731 -9320 15732 -8600
rect 16452 -9320 16453 -8600
rect 15731 -9321 16453 -9320
rect 15312 -9388 15408 -9372
rect 16724 -9372 16740 -8548
rect 16804 -9372 16820 -8548
rect 18136 -8548 18232 -8532
rect 17143 -8600 17865 -8599
rect 17143 -9320 17144 -8600
rect 17864 -9320 17865 -8600
rect 17143 -9321 17865 -9320
rect 16724 -9388 16820 -9372
rect 18136 -9372 18152 -8548
rect 18216 -9372 18232 -8548
rect 19548 -8548 19644 -8532
rect 18555 -8600 19277 -8599
rect 18555 -9320 18556 -8600
rect 19276 -9320 19277 -8600
rect 18555 -9321 19277 -9320
rect 18136 -9388 18232 -9372
rect 19548 -9372 19564 -8548
rect 19628 -9372 19644 -8548
rect 20960 -8548 21056 -8532
rect 19967 -8600 20689 -8599
rect 19967 -9320 19968 -8600
rect 20688 -9320 20689 -8600
rect 19967 -9321 20689 -9320
rect 19548 -9388 19644 -9372
rect 20960 -9372 20976 -8548
rect 21040 -9372 21056 -8548
rect 22372 -8548 22468 -8532
rect 21379 -8600 22101 -8599
rect 21379 -9320 21380 -8600
rect 22100 -9320 22101 -8600
rect 21379 -9321 22101 -9320
rect 20960 -9388 21056 -9372
rect 22372 -9372 22388 -8548
rect 22452 -9372 22468 -8548
rect 23784 -8548 23880 -8532
rect 22791 -8600 23513 -8599
rect 22791 -9320 22792 -8600
rect 23512 -9320 23513 -8600
rect 22791 -9321 23513 -9320
rect 22372 -9388 22468 -9372
rect 23784 -9372 23800 -8548
rect 23864 -9372 23880 -8548
rect 23784 -9388 23880 -9372
rect -22812 -9668 -22716 -9652
rect -23805 -9720 -23083 -9719
rect -23805 -10440 -23804 -9720
rect -23084 -10440 -23083 -9720
rect -23805 -10441 -23083 -10440
rect -22812 -10492 -22796 -9668
rect -22732 -10492 -22716 -9668
rect -21400 -9668 -21304 -9652
rect -22393 -9720 -21671 -9719
rect -22393 -10440 -22392 -9720
rect -21672 -10440 -21671 -9720
rect -22393 -10441 -21671 -10440
rect -22812 -10508 -22716 -10492
rect -21400 -10492 -21384 -9668
rect -21320 -10492 -21304 -9668
rect -19988 -9668 -19892 -9652
rect -20981 -9720 -20259 -9719
rect -20981 -10440 -20980 -9720
rect -20260 -10440 -20259 -9720
rect -20981 -10441 -20259 -10440
rect -21400 -10508 -21304 -10492
rect -19988 -10492 -19972 -9668
rect -19908 -10492 -19892 -9668
rect -18576 -9668 -18480 -9652
rect -19569 -9720 -18847 -9719
rect -19569 -10440 -19568 -9720
rect -18848 -10440 -18847 -9720
rect -19569 -10441 -18847 -10440
rect -19988 -10508 -19892 -10492
rect -18576 -10492 -18560 -9668
rect -18496 -10492 -18480 -9668
rect -17164 -9668 -17068 -9652
rect -18157 -9720 -17435 -9719
rect -18157 -10440 -18156 -9720
rect -17436 -10440 -17435 -9720
rect -18157 -10441 -17435 -10440
rect -18576 -10508 -18480 -10492
rect -17164 -10492 -17148 -9668
rect -17084 -10492 -17068 -9668
rect -15752 -9668 -15656 -9652
rect -16745 -9720 -16023 -9719
rect -16745 -10440 -16744 -9720
rect -16024 -10440 -16023 -9720
rect -16745 -10441 -16023 -10440
rect -17164 -10508 -17068 -10492
rect -15752 -10492 -15736 -9668
rect -15672 -10492 -15656 -9668
rect -14340 -9668 -14244 -9652
rect -15333 -9720 -14611 -9719
rect -15333 -10440 -15332 -9720
rect -14612 -10440 -14611 -9720
rect -15333 -10441 -14611 -10440
rect -15752 -10508 -15656 -10492
rect -14340 -10492 -14324 -9668
rect -14260 -10492 -14244 -9668
rect -12928 -9668 -12832 -9652
rect -13921 -9720 -13199 -9719
rect -13921 -10440 -13920 -9720
rect -13200 -10440 -13199 -9720
rect -13921 -10441 -13199 -10440
rect -14340 -10508 -14244 -10492
rect -12928 -10492 -12912 -9668
rect -12848 -10492 -12832 -9668
rect -11516 -9668 -11420 -9652
rect -12509 -9720 -11787 -9719
rect -12509 -10440 -12508 -9720
rect -11788 -10440 -11787 -9720
rect -12509 -10441 -11787 -10440
rect -12928 -10508 -12832 -10492
rect -11516 -10492 -11500 -9668
rect -11436 -10492 -11420 -9668
rect -10104 -9668 -10008 -9652
rect -11097 -9720 -10375 -9719
rect -11097 -10440 -11096 -9720
rect -10376 -10440 -10375 -9720
rect -11097 -10441 -10375 -10440
rect -11516 -10508 -11420 -10492
rect -10104 -10492 -10088 -9668
rect -10024 -10492 -10008 -9668
rect -8692 -9668 -8596 -9652
rect -9685 -9720 -8963 -9719
rect -9685 -10440 -9684 -9720
rect -8964 -10440 -8963 -9720
rect -9685 -10441 -8963 -10440
rect -10104 -10508 -10008 -10492
rect -8692 -10492 -8676 -9668
rect -8612 -10492 -8596 -9668
rect -7280 -9668 -7184 -9652
rect -8273 -9720 -7551 -9719
rect -8273 -10440 -8272 -9720
rect -7552 -10440 -7551 -9720
rect -8273 -10441 -7551 -10440
rect -8692 -10508 -8596 -10492
rect -7280 -10492 -7264 -9668
rect -7200 -10492 -7184 -9668
rect -5868 -9668 -5772 -9652
rect -6861 -9720 -6139 -9719
rect -6861 -10440 -6860 -9720
rect -6140 -10440 -6139 -9720
rect -6861 -10441 -6139 -10440
rect -7280 -10508 -7184 -10492
rect -5868 -10492 -5852 -9668
rect -5788 -10492 -5772 -9668
rect -4456 -9668 -4360 -9652
rect -5449 -9720 -4727 -9719
rect -5449 -10440 -5448 -9720
rect -4728 -10440 -4727 -9720
rect -5449 -10441 -4727 -10440
rect -5868 -10508 -5772 -10492
rect -4456 -10492 -4440 -9668
rect -4376 -10492 -4360 -9668
rect -3044 -9668 -2948 -9652
rect -4037 -9720 -3315 -9719
rect -4037 -10440 -4036 -9720
rect -3316 -10440 -3315 -9720
rect -4037 -10441 -3315 -10440
rect -4456 -10508 -4360 -10492
rect -3044 -10492 -3028 -9668
rect -2964 -10492 -2948 -9668
rect -1632 -9668 -1536 -9652
rect -2625 -9720 -1903 -9719
rect -2625 -10440 -2624 -9720
rect -1904 -10440 -1903 -9720
rect -2625 -10441 -1903 -10440
rect -3044 -10508 -2948 -10492
rect -1632 -10492 -1616 -9668
rect -1552 -10492 -1536 -9668
rect -220 -9668 -124 -9652
rect -1213 -9720 -491 -9719
rect -1213 -10440 -1212 -9720
rect -492 -10440 -491 -9720
rect -1213 -10441 -491 -10440
rect -1632 -10508 -1536 -10492
rect -220 -10492 -204 -9668
rect -140 -10492 -124 -9668
rect 1192 -9668 1288 -9652
rect 199 -9720 921 -9719
rect 199 -10440 200 -9720
rect 920 -10440 921 -9720
rect 199 -10441 921 -10440
rect -220 -10508 -124 -10492
rect 1192 -10492 1208 -9668
rect 1272 -10492 1288 -9668
rect 2604 -9668 2700 -9652
rect 1611 -9720 2333 -9719
rect 1611 -10440 1612 -9720
rect 2332 -10440 2333 -9720
rect 1611 -10441 2333 -10440
rect 1192 -10508 1288 -10492
rect 2604 -10492 2620 -9668
rect 2684 -10492 2700 -9668
rect 4016 -9668 4112 -9652
rect 3023 -9720 3745 -9719
rect 3023 -10440 3024 -9720
rect 3744 -10440 3745 -9720
rect 3023 -10441 3745 -10440
rect 2604 -10508 2700 -10492
rect 4016 -10492 4032 -9668
rect 4096 -10492 4112 -9668
rect 5428 -9668 5524 -9652
rect 4435 -9720 5157 -9719
rect 4435 -10440 4436 -9720
rect 5156 -10440 5157 -9720
rect 4435 -10441 5157 -10440
rect 4016 -10508 4112 -10492
rect 5428 -10492 5444 -9668
rect 5508 -10492 5524 -9668
rect 6840 -9668 6936 -9652
rect 5847 -9720 6569 -9719
rect 5847 -10440 5848 -9720
rect 6568 -10440 6569 -9720
rect 5847 -10441 6569 -10440
rect 5428 -10508 5524 -10492
rect 6840 -10492 6856 -9668
rect 6920 -10492 6936 -9668
rect 8252 -9668 8348 -9652
rect 7259 -9720 7981 -9719
rect 7259 -10440 7260 -9720
rect 7980 -10440 7981 -9720
rect 7259 -10441 7981 -10440
rect 6840 -10508 6936 -10492
rect 8252 -10492 8268 -9668
rect 8332 -10492 8348 -9668
rect 9664 -9668 9760 -9652
rect 8671 -9720 9393 -9719
rect 8671 -10440 8672 -9720
rect 9392 -10440 9393 -9720
rect 8671 -10441 9393 -10440
rect 8252 -10508 8348 -10492
rect 9664 -10492 9680 -9668
rect 9744 -10492 9760 -9668
rect 11076 -9668 11172 -9652
rect 10083 -9720 10805 -9719
rect 10083 -10440 10084 -9720
rect 10804 -10440 10805 -9720
rect 10083 -10441 10805 -10440
rect 9664 -10508 9760 -10492
rect 11076 -10492 11092 -9668
rect 11156 -10492 11172 -9668
rect 12488 -9668 12584 -9652
rect 11495 -9720 12217 -9719
rect 11495 -10440 11496 -9720
rect 12216 -10440 12217 -9720
rect 11495 -10441 12217 -10440
rect 11076 -10508 11172 -10492
rect 12488 -10492 12504 -9668
rect 12568 -10492 12584 -9668
rect 13900 -9668 13996 -9652
rect 12907 -9720 13629 -9719
rect 12907 -10440 12908 -9720
rect 13628 -10440 13629 -9720
rect 12907 -10441 13629 -10440
rect 12488 -10508 12584 -10492
rect 13900 -10492 13916 -9668
rect 13980 -10492 13996 -9668
rect 15312 -9668 15408 -9652
rect 14319 -9720 15041 -9719
rect 14319 -10440 14320 -9720
rect 15040 -10440 15041 -9720
rect 14319 -10441 15041 -10440
rect 13900 -10508 13996 -10492
rect 15312 -10492 15328 -9668
rect 15392 -10492 15408 -9668
rect 16724 -9668 16820 -9652
rect 15731 -9720 16453 -9719
rect 15731 -10440 15732 -9720
rect 16452 -10440 16453 -9720
rect 15731 -10441 16453 -10440
rect 15312 -10508 15408 -10492
rect 16724 -10492 16740 -9668
rect 16804 -10492 16820 -9668
rect 18136 -9668 18232 -9652
rect 17143 -9720 17865 -9719
rect 17143 -10440 17144 -9720
rect 17864 -10440 17865 -9720
rect 17143 -10441 17865 -10440
rect 16724 -10508 16820 -10492
rect 18136 -10492 18152 -9668
rect 18216 -10492 18232 -9668
rect 19548 -9668 19644 -9652
rect 18555 -9720 19277 -9719
rect 18555 -10440 18556 -9720
rect 19276 -10440 19277 -9720
rect 18555 -10441 19277 -10440
rect 18136 -10508 18232 -10492
rect 19548 -10492 19564 -9668
rect 19628 -10492 19644 -9668
rect 20960 -9668 21056 -9652
rect 19967 -9720 20689 -9719
rect 19967 -10440 19968 -9720
rect 20688 -10440 20689 -9720
rect 19967 -10441 20689 -10440
rect 19548 -10508 19644 -10492
rect 20960 -10492 20976 -9668
rect 21040 -10492 21056 -9668
rect 22372 -9668 22468 -9652
rect 21379 -9720 22101 -9719
rect 21379 -10440 21380 -9720
rect 22100 -10440 22101 -9720
rect 21379 -10441 22101 -10440
rect 20960 -10508 21056 -10492
rect 22372 -10492 22388 -9668
rect 22452 -10492 22468 -9668
rect 23784 -9668 23880 -9652
rect 22791 -9720 23513 -9719
rect 22791 -10440 22792 -9720
rect 23512 -10440 23513 -9720
rect 22791 -10441 23513 -10440
rect 22372 -10508 22468 -10492
rect 23784 -10492 23800 -9668
rect 23864 -10492 23880 -9668
rect 23784 -10508 23880 -10492
rect -22812 -10788 -22716 -10772
rect -23805 -10840 -23083 -10839
rect -23805 -11560 -23804 -10840
rect -23084 -11560 -23083 -10840
rect -23805 -11561 -23083 -11560
rect -22812 -11612 -22796 -10788
rect -22732 -11612 -22716 -10788
rect -21400 -10788 -21304 -10772
rect -22393 -10840 -21671 -10839
rect -22393 -11560 -22392 -10840
rect -21672 -11560 -21671 -10840
rect -22393 -11561 -21671 -11560
rect -22812 -11628 -22716 -11612
rect -21400 -11612 -21384 -10788
rect -21320 -11612 -21304 -10788
rect -19988 -10788 -19892 -10772
rect -20981 -10840 -20259 -10839
rect -20981 -11560 -20980 -10840
rect -20260 -11560 -20259 -10840
rect -20981 -11561 -20259 -11560
rect -21400 -11628 -21304 -11612
rect -19988 -11612 -19972 -10788
rect -19908 -11612 -19892 -10788
rect -18576 -10788 -18480 -10772
rect -19569 -10840 -18847 -10839
rect -19569 -11560 -19568 -10840
rect -18848 -11560 -18847 -10840
rect -19569 -11561 -18847 -11560
rect -19988 -11628 -19892 -11612
rect -18576 -11612 -18560 -10788
rect -18496 -11612 -18480 -10788
rect -17164 -10788 -17068 -10772
rect -18157 -10840 -17435 -10839
rect -18157 -11560 -18156 -10840
rect -17436 -11560 -17435 -10840
rect -18157 -11561 -17435 -11560
rect -18576 -11628 -18480 -11612
rect -17164 -11612 -17148 -10788
rect -17084 -11612 -17068 -10788
rect -15752 -10788 -15656 -10772
rect -16745 -10840 -16023 -10839
rect -16745 -11560 -16744 -10840
rect -16024 -11560 -16023 -10840
rect -16745 -11561 -16023 -11560
rect -17164 -11628 -17068 -11612
rect -15752 -11612 -15736 -10788
rect -15672 -11612 -15656 -10788
rect -14340 -10788 -14244 -10772
rect -15333 -10840 -14611 -10839
rect -15333 -11560 -15332 -10840
rect -14612 -11560 -14611 -10840
rect -15333 -11561 -14611 -11560
rect -15752 -11628 -15656 -11612
rect -14340 -11612 -14324 -10788
rect -14260 -11612 -14244 -10788
rect -12928 -10788 -12832 -10772
rect -13921 -10840 -13199 -10839
rect -13921 -11560 -13920 -10840
rect -13200 -11560 -13199 -10840
rect -13921 -11561 -13199 -11560
rect -14340 -11628 -14244 -11612
rect -12928 -11612 -12912 -10788
rect -12848 -11612 -12832 -10788
rect -11516 -10788 -11420 -10772
rect -12509 -10840 -11787 -10839
rect -12509 -11560 -12508 -10840
rect -11788 -11560 -11787 -10840
rect -12509 -11561 -11787 -11560
rect -12928 -11628 -12832 -11612
rect -11516 -11612 -11500 -10788
rect -11436 -11612 -11420 -10788
rect -10104 -10788 -10008 -10772
rect -11097 -10840 -10375 -10839
rect -11097 -11560 -11096 -10840
rect -10376 -11560 -10375 -10840
rect -11097 -11561 -10375 -11560
rect -11516 -11628 -11420 -11612
rect -10104 -11612 -10088 -10788
rect -10024 -11612 -10008 -10788
rect -8692 -10788 -8596 -10772
rect -9685 -10840 -8963 -10839
rect -9685 -11560 -9684 -10840
rect -8964 -11560 -8963 -10840
rect -9685 -11561 -8963 -11560
rect -10104 -11628 -10008 -11612
rect -8692 -11612 -8676 -10788
rect -8612 -11612 -8596 -10788
rect -7280 -10788 -7184 -10772
rect -8273 -10840 -7551 -10839
rect -8273 -11560 -8272 -10840
rect -7552 -11560 -7551 -10840
rect -8273 -11561 -7551 -11560
rect -8692 -11628 -8596 -11612
rect -7280 -11612 -7264 -10788
rect -7200 -11612 -7184 -10788
rect -5868 -10788 -5772 -10772
rect -6861 -10840 -6139 -10839
rect -6861 -11560 -6860 -10840
rect -6140 -11560 -6139 -10840
rect -6861 -11561 -6139 -11560
rect -7280 -11628 -7184 -11612
rect -5868 -11612 -5852 -10788
rect -5788 -11612 -5772 -10788
rect -4456 -10788 -4360 -10772
rect -5449 -10840 -4727 -10839
rect -5449 -11560 -5448 -10840
rect -4728 -11560 -4727 -10840
rect -5449 -11561 -4727 -11560
rect -5868 -11628 -5772 -11612
rect -4456 -11612 -4440 -10788
rect -4376 -11612 -4360 -10788
rect -3044 -10788 -2948 -10772
rect -4037 -10840 -3315 -10839
rect -4037 -11560 -4036 -10840
rect -3316 -11560 -3315 -10840
rect -4037 -11561 -3315 -11560
rect -4456 -11628 -4360 -11612
rect -3044 -11612 -3028 -10788
rect -2964 -11612 -2948 -10788
rect -1632 -10788 -1536 -10772
rect -2625 -10840 -1903 -10839
rect -2625 -11560 -2624 -10840
rect -1904 -11560 -1903 -10840
rect -2625 -11561 -1903 -11560
rect -3044 -11628 -2948 -11612
rect -1632 -11612 -1616 -10788
rect -1552 -11612 -1536 -10788
rect -220 -10788 -124 -10772
rect -1213 -10840 -491 -10839
rect -1213 -11560 -1212 -10840
rect -492 -11560 -491 -10840
rect -1213 -11561 -491 -11560
rect -1632 -11628 -1536 -11612
rect -220 -11612 -204 -10788
rect -140 -11612 -124 -10788
rect 1192 -10788 1288 -10772
rect 199 -10840 921 -10839
rect 199 -11560 200 -10840
rect 920 -11560 921 -10840
rect 199 -11561 921 -11560
rect -220 -11628 -124 -11612
rect 1192 -11612 1208 -10788
rect 1272 -11612 1288 -10788
rect 2604 -10788 2700 -10772
rect 1611 -10840 2333 -10839
rect 1611 -11560 1612 -10840
rect 2332 -11560 2333 -10840
rect 1611 -11561 2333 -11560
rect 1192 -11628 1288 -11612
rect 2604 -11612 2620 -10788
rect 2684 -11612 2700 -10788
rect 4016 -10788 4112 -10772
rect 3023 -10840 3745 -10839
rect 3023 -11560 3024 -10840
rect 3744 -11560 3745 -10840
rect 3023 -11561 3745 -11560
rect 2604 -11628 2700 -11612
rect 4016 -11612 4032 -10788
rect 4096 -11612 4112 -10788
rect 5428 -10788 5524 -10772
rect 4435 -10840 5157 -10839
rect 4435 -11560 4436 -10840
rect 5156 -11560 5157 -10840
rect 4435 -11561 5157 -11560
rect 4016 -11628 4112 -11612
rect 5428 -11612 5444 -10788
rect 5508 -11612 5524 -10788
rect 6840 -10788 6936 -10772
rect 5847 -10840 6569 -10839
rect 5847 -11560 5848 -10840
rect 6568 -11560 6569 -10840
rect 5847 -11561 6569 -11560
rect 5428 -11628 5524 -11612
rect 6840 -11612 6856 -10788
rect 6920 -11612 6936 -10788
rect 8252 -10788 8348 -10772
rect 7259 -10840 7981 -10839
rect 7259 -11560 7260 -10840
rect 7980 -11560 7981 -10840
rect 7259 -11561 7981 -11560
rect 6840 -11628 6936 -11612
rect 8252 -11612 8268 -10788
rect 8332 -11612 8348 -10788
rect 9664 -10788 9760 -10772
rect 8671 -10840 9393 -10839
rect 8671 -11560 8672 -10840
rect 9392 -11560 9393 -10840
rect 8671 -11561 9393 -11560
rect 8252 -11628 8348 -11612
rect 9664 -11612 9680 -10788
rect 9744 -11612 9760 -10788
rect 11076 -10788 11172 -10772
rect 10083 -10840 10805 -10839
rect 10083 -11560 10084 -10840
rect 10804 -11560 10805 -10840
rect 10083 -11561 10805 -11560
rect 9664 -11628 9760 -11612
rect 11076 -11612 11092 -10788
rect 11156 -11612 11172 -10788
rect 12488 -10788 12584 -10772
rect 11495 -10840 12217 -10839
rect 11495 -11560 11496 -10840
rect 12216 -11560 12217 -10840
rect 11495 -11561 12217 -11560
rect 11076 -11628 11172 -11612
rect 12488 -11612 12504 -10788
rect 12568 -11612 12584 -10788
rect 13900 -10788 13996 -10772
rect 12907 -10840 13629 -10839
rect 12907 -11560 12908 -10840
rect 13628 -11560 13629 -10840
rect 12907 -11561 13629 -11560
rect 12488 -11628 12584 -11612
rect 13900 -11612 13916 -10788
rect 13980 -11612 13996 -10788
rect 15312 -10788 15408 -10772
rect 14319 -10840 15041 -10839
rect 14319 -11560 14320 -10840
rect 15040 -11560 15041 -10840
rect 14319 -11561 15041 -11560
rect 13900 -11628 13996 -11612
rect 15312 -11612 15328 -10788
rect 15392 -11612 15408 -10788
rect 16724 -10788 16820 -10772
rect 15731 -10840 16453 -10839
rect 15731 -11560 15732 -10840
rect 16452 -11560 16453 -10840
rect 15731 -11561 16453 -11560
rect 15312 -11628 15408 -11612
rect 16724 -11612 16740 -10788
rect 16804 -11612 16820 -10788
rect 18136 -10788 18232 -10772
rect 17143 -10840 17865 -10839
rect 17143 -11560 17144 -10840
rect 17864 -11560 17865 -10840
rect 17143 -11561 17865 -11560
rect 16724 -11628 16820 -11612
rect 18136 -11612 18152 -10788
rect 18216 -11612 18232 -10788
rect 19548 -10788 19644 -10772
rect 18555 -10840 19277 -10839
rect 18555 -11560 18556 -10840
rect 19276 -11560 19277 -10840
rect 18555 -11561 19277 -11560
rect 18136 -11628 18232 -11612
rect 19548 -11612 19564 -10788
rect 19628 -11612 19644 -10788
rect 20960 -10788 21056 -10772
rect 19967 -10840 20689 -10839
rect 19967 -11560 19968 -10840
rect 20688 -11560 20689 -10840
rect 19967 -11561 20689 -11560
rect 19548 -11628 19644 -11612
rect 20960 -11612 20976 -10788
rect 21040 -11612 21056 -10788
rect 22372 -10788 22468 -10772
rect 21379 -10840 22101 -10839
rect 21379 -11560 21380 -10840
rect 22100 -11560 22101 -10840
rect 21379 -11561 22101 -11560
rect 20960 -11628 21056 -11612
rect 22372 -11612 22388 -10788
rect 22452 -11612 22468 -10788
rect 23784 -10788 23880 -10772
rect 22791 -10840 23513 -10839
rect 22791 -11560 22792 -10840
rect 23512 -11560 23513 -10840
rect 22791 -11561 23513 -11560
rect 22372 -11628 22468 -11612
rect 23784 -11612 23800 -10788
rect 23864 -11612 23880 -10788
rect 23784 -11628 23880 -11612
rect -22812 -11908 -22716 -11892
rect -23805 -11960 -23083 -11959
rect -23805 -12680 -23804 -11960
rect -23084 -12680 -23083 -11960
rect -23805 -12681 -23083 -12680
rect -22812 -12732 -22796 -11908
rect -22732 -12732 -22716 -11908
rect -21400 -11908 -21304 -11892
rect -22393 -11960 -21671 -11959
rect -22393 -12680 -22392 -11960
rect -21672 -12680 -21671 -11960
rect -22393 -12681 -21671 -12680
rect -22812 -12748 -22716 -12732
rect -21400 -12732 -21384 -11908
rect -21320 -12732 -21304 -11908
rect -19988 -11908 -19892 -11892
rect -20981 -11960 -20259 -11959
rect -20981 -12680 -20980 -11960
rect -20260 -12680 -20259 -11960
rect -20981 -12681 -20259 -12680
rect -21400 -12748 -21304 -12732
rect -19988 -12732 -19972 -11908
rect -19908 -12732 -19892 -11908
rect -18576 -11908 -18480 -11892
rect -19569 -11960 -18847 -11959
rect -19569 -12680 -19568 -11960
rect -18848 -12680 -18847 -11960
rect -19569 -12681 -18847 -12680
rect -19988 -12748 -19892 -12732
rect -18576 -12732 -18560 -11908
rect -18496 -12732 -18480 -11908
rect -17164 -11908 -17068 -11892
rect -18157 -11960 -17435 -11959
rect -18157 -12680 -18156 -11960
rect -17436 -12680 -17435 -11960
rect -18157 -12681 -17435 -12680
rect -18576 -12748 -18480 -12732
rect -17164 -12732 -17148 -11908
rect -17084 -12732 -17068 -11908
rect -15752 -11908 -15656 -11892
rect -16745 -11960 -16023 -11959
rect -16745 -12680 -16744 -11960
rect -16024 -12680 -16023 -11960
rect -16745 -12681 -16023 -12680
rect -17164 -12748 -17068 -12732
rect -15752 -12732 -15736 -11908
rect -15672 -12732 -15656 -11908
rect -14340 -11908 -14244 -11892
rect -15333 -11960 -14611 -11959
rect -15333 -12680 -15332 -11960
rect -14612 -12680 -14611 -11960
rect -15333 -12681 -14611 -12680
rect -15752 -12748 -15656 -12732
rect -14340 -12732 -14324 -11908
rect -14260 -12732 -14244 -11908
rect -12928 -11908 -12832 -11892
rect -13921 -11960 -13199 -11959
rect -13921 -12680 -13920 -11960
rect -13200 -12680 -13199 -11960
rect -13921 -12681 -13199 -12680
rect -14340 -12748 -14244 -12732
rect -12928 -12732 -12912 -11908
rect -12848 -12732 -12832 -11908
rect -11516 -11908 -11420 -11892
rect -12509 -11960 -11787 -11959
rect -12509 -12680 -12508 -11960
rect -11788 -12680 -11787 -11960
rect -12509 -12681 -11787 -12680
rect -12928 -12748 -12832 -12732
rect -11516 -12732 -11500 -11908
rect -11436 -12732 -11420 -11908
rect -10104 -11908 -10008 -11892
rect -11097 -11960 -10375 -11959
rect -11097 -12680 -11096 -11960
rect -10376 -12680 -10375 -11960
rect -11097 -12681 -10375 -12680
rect -11516 -12748 -11420 -12732
rect -10104 -12732 -10088 -11908
rect -10024 -12732 -10008 -11908
rect -8692 -11908 -8596 -11892
rect -9685 -11960 -8963 -11959
rect -9685 -12680 -9684 -11960
rect -8964 -12680 -8963 -11960
rect -9685 -12681 -8963 -12680
rect -10104 -12748 -10008 -12732
rect -8692 -12732 -8676 -11908
rect -8612 -12732 -8596 -11908
rect -7280 -11908 -7184 -11892
rect -8273 -11960 -7551 -11959
rect -8273 -12680 -8272 -11960
rect -7552 -12680 -7551 -11960
rect -8273 -12681 -7551 -12680
rect -8692 -12748 -8596 -12732
rect -7280 -12732 -7264 -11908
rect -7200 -12732 -7184 -11908
rect -5868 -11908 -5772 -11892
rect -6861 -11960 -6139 -11959
rect -6861 -12680 -6860 -11960
rect -6140 -12680 -6139 -11960
rect -6861 -12681 -6139 -12680
rect -7280 -12748 -7184 -12732
rect -5868 -12732 -5852 -11908
rect -5788 -12732 -5772 -11908
rect -4456 -11908 -4360 -11892
rect -5449 -11960 -4727 -11959
rect -5449 -12680 -5448 -11960
rect -4728 -12680 -4727 -11960
rect -5449 -12681 -4727 -12680
rect -5868 -12748 -5772 -12732
rect -4456 -12732 -4440 -11908
rect -4376 -12732 -4360 -11908
rect -3044 -11908 -2948 -11892
rect -4037 -11960 -3315 -11959
rect -4037 -12680 -4036 -11960
rect -3316 -12680 -3315 -11960
rect -4037 -12681 -3315 -12680
rect -4456 -12748 -4360 -12732
rect -3044 -12732 -3028 -11908
rect -2964 -12732 -2948 -11908
rect -1632 -11908 -1536 -11892
rect -2625 -11960 -1903 -11959
rect -2625 -12680 -2624 -11960
rect -1904 -12680 -1903 -11960
rect -2625 -12681 -1903 -12680
rect -3044 -12748 -2948 -12732
rect -1632 -12732 -1616 -11908
rect -1552 -12732 -1536 -11908
rect -220 -11908 -124 -11892
rect -1213 -11960 -491 -11959
rect -1213 -12680 -1212 -11960
rect -492 -12680 -491 -11960
rect -1213 -12681 -491 -12680
rect -1632 -12748 -1536 -12732
rect -220 -12732 -204 -11908
rect -140 -12732 -124 -11908
rect 1192 -11908 1288 -11892
rect 199 -11960 921 -11959
rect 199 -12680 200 -11960
rect 920 -12680 921 -11960
rect 199 -12681 921 -12680
rect -220 -12748 -124 -12732
rect 1192 -12732 1208 -11908
rect 1272 -12732 1288 -11908
rect 2604 -11908 2700 -11892
rect 1611 -11960 2333 -11959
rect 1611 -12680 1612 -11960
rect 2332 -12680 2333 -11960
rect 1611 -12681 2333 -12680
rect 1192 -12748 1288 -12732
rect 2604 -12732 2620 -11908
rect 2684 -12732 2700 -11908
rect 4016 -11908 4112 -11892
rect 3023 -11960 3745 -11959
rect 3023 -12680 3024 -11960
rect 3744 -12680 3745 -11960
rect 3023 -12681 3745 -12680
rect 2604 -12748 2700 -12732
rect 4016 -12732 4032 -11908
rect 4096 -12732 4112 -11908
rect 5428 -11908 5524 -11892
rect 4435 -11960 5157 -11959
rect 4435 -12680 4436 -11960
rect 5156 -12680 5157 -11960
rect 4435 -12681 5157 -12680
rect 4016 -12748 4112 -12732
rect 5428 -12732 5444 -11908
rect 5508 -12732 5524 -11908
rect 6840 -11908 6936 -11892
rect 5847 -11960 6569 -11959
rect 5847 -12680 5848 -11960
rect 6568 -12680 6569 -11960
rect 5847 -12681 6569 -12680
rect 5428 -12748 5524 -12732
rect 6840 -12732 6856 -11908
rect 6920 -12732 6936 -11908
rect 8252 -11908 8348 -11892
rect 7259 -11960 7981 -11959
rect 7259 -12680 7260 -11960
rect 7980 -12680 7981 -11960
rect 7259 -12681 7981 -12680
rect 6840 -12748 6936 -12732
rect 8252 -12732 8268 -11908
rect 8332 -12732 8348 -11908
rect 9664 -11908 9760 -11892
rect 8671 -11960 9393 -11959
rect 8671 -12680 8672 -11960
rect 9392 -12680 9393 -11960
rect 8671 -12681 9393 -12680
rect 8252 -12748 8348 -12732
rect 9664 -12732 9680 -11908
rect 9744 -12732 9760 -11908
rect 11076 -11908 11172 -11892
rect 10083 -11960 10805 -11959
rect 10083 -12680 10084 -11960
rect 10804 -12680 10805 -11960
rect 10083 -12681 10805 -12680
rect 9664 -12748 9760 -12732
rect 11076 -12732 11092 -11908
rect 11156 -12732 11172 -11908
rect 12488 -11908 12584 -11892
rect 11495 -11960 12217 -11959
rect 11495 -12680 11496 -11960
rect 12216 -12680 12217 -11960
rect 11495 -12681 12217 -12680
rect 11076 -12748 11172 -12732
rect 12488 -12732 12504 -11908
rect 12568 -12732 12584 -11908
rect 13900 -11908 13996 -11892
rect 12907 -11960 13629 -11959
rect 12907 -12680 12908 -11960
rect 13628 -12680 13629 -11960
rect 12907 -12681 13629 -12680
rect 12488 -12748 12584 -12732
rect 13900 -12732 13916 -11908
rect 13980 -12732 13996 -11908
rect 15312 -11908 15408 -11892
rect 14319 -11960 15041 -11959
rect 14319 -12680 14320 -11960
rect 15040 -12680 15041 -11960
rect 14319 -12681 15041 -12680
rect 13900 -12748 13996 -12732
rect 15312 -12732 15328 -11908
rect 15392 -12732 15408 -11908
rect 16724 -11908 16820 -11892
rect 15731 -11960 16453 -11959
rect 15731 -12680 15732 -11960
rect 16452 -12680 16453 -11960
rect 15731 -12681 16453 -12680
rect 15312 -12748 15408 -12732
rect 16724 -12732 16740 -11908
rect 16804 -12732 16820 -11908
rect 18136 -11908 18232 -11892
rect 17143 -11960 17865 -11959
rect 17143 -12680 17144 -11960
rect 17864 -12680 17865 -11960
rect 17143 -12681 17865 -12680
rect 16724 -12748 16820 -12732
rect 18136 -12732 18152 -11908
rect 18216 -12732 18232 -11908
rect 19548 -11908 19644 -11892
rect 18555 -11960 19277 -11959
rect 18555 -12680 18556 -11960
rect 19276 -12680 19277 -11960
rect 18555 -12681 19277 -12680
rect 18136 -12748 18232 -12732
rect 19548 -12732 19564 -11908
rect 19628 -12732 19644 -11908
rect 20960 -11908 21056 -11892
rect 19967 -11960 20689 -11959
rect 19967 -12680 19968 -11960
rect 20688 -12680 20689 -11960
rect 19967 -12681 20689 -12680
rect 19548 -12748 19644 -12732
rect 20960 -12732 20976 -11908
rect 21040 -12732 21056 -11908
rect 22372 -11908 22468 -11892
rect 21379 -11960 22101 -11959
rect 21379 -12680 21380 -11960
rect 22100 -12680 22101 -11960
rect 21379 -12681 22101 -12680
rect 20960 -12748 21056 -12732
rect 22372 -12732 22388 -11908
rect 22452 -12732 22468 -11908
rect 23784 -11908 23880 -11892
rect 22791 -11960 23513 -11959
rect 22791 -12680 22792 -11960
rect 23512 -12680 23513 -11960
rect 22791 -12681 23513 -12680
rect 22372 -12748 22468 -12732
rect 23784 -12732 23800 -11908
rect 23864 -12732 23880 -11908
rect 23784 -12748 23880 -12732
rect -22812 -13028 -22716 -13012
rect -23805 -13080 -23083 -13079
rect -23805 -13800 -23804 -13080
rect -23084 -13800 -23083 -13080
rect -23805 -13801 -23083 -13800
rect -22812 -13852 -22796 -13028
rect -22732 -13852 -22716 -13028
rect -21400 -13028 -21304 -13012
rect -22393 -13080 -21671 -13079
rect -22393 -13800 -22392 -13080
rect -21672 -13800 -21671 -13080
rect -22393 -13801 -21671 -13800
rect -22812 -13868 -22716 -13852
rect -21400 -13852 -21384 -13028
rect -21320 -13852 -21304 -13028
rect -19988 -13028 -19892 -13012
rect -20981 -13080 -20259 -13079
rect -20981 -13800 -20980 -13080
rect -20260 -13800 -20259 -13080
rect -20981 -13801 -20259 -13800
rect -21400 -13868 -21304 -13852
rect -19988 -13852 -19972 -13028
rect -19908 -13852 -19892 -13028
rect -18576 -13028 -18480 -13012
rect -19569 -13080 -18847 -13079
rect -19569 -13800 -19568 -13080
rect -18848 -13800 -18847 -13080
rect -19569 -13801 -18847 -13800
rect -19988 -13868 -19892 -13852
rect -18576 -13852 -18560 -13028
rect -18496 -13852 -18480 -13028
rect -17164 -13028 -17068 -13012
rect -18157 -13080 -17435 -13079
rect -18157 -13800 -18156 -13080
rect -17436 -13800 -17435 -13080
rect -18157 -13801 -17435 -13800
rect -18576 -13868 -18480 -13852
rect -17164 -13852 -17148 -13028
rect -17084 -13852 -17068 -13028
rect -15752 -13028 -15656 -13012
rect -16745 -13080 -16023 -13079
rect -16745 -13800 -16744 -13080
rect -16024 -13800 -16023 -13080
rect -16745 -13801 -16023 -13800
rect -17164 -13868 -17068 -13852
rect -15752 -13852 -15736 -13028
rect -15672 -13852 -15656 -13028
rect -14340 -13028 -14244 -13012
rect -15333 -13080 -14611 -13079
rect -15333 -13800 -15332 -13080
rect -14612 -13800 -14611 -13080
rect -15333 -13801 -14611 -13800
rect -15752 -13868 -15656 -13852
rect -14340 -13852 -14324 -13028
rect -14260 -13852 -14244 -13028
rect -12928 -13028 -12832 -13012
rect -13921 -13080 -13199 -13079
rect -13921 -13800 -13920 -13080
rect -13200 -13800 -13199 -13080
rect -13921 -13801 -13199 -13800
rect -14340 -13868 -14244 -13852
rect -12928 -13852 -12912 -13028
rect -12848 -13852 -12832 -13028
rect -11516 -13028 -11420 -13012
rect -12509 -13080 -11787 -13079
rect -12509 -13800 -12508 -13080
rect -11788 -13800 -11787 -13080
rect -12509 -13801 -11787 -13800
rect -12928 -13868 -12832 -13852
rect -11516 -13852 -11500 -13028
rect -11436 -13852 -11420 -13028
rect -10104 -13028 -10008 -13012
rect -11097 -13080 -10375 -13079
rect -11097 -13800 -11096 -13080
rect -10376 -13800 -10375 -13080
rect -11097 -13801 -10375 -13800
rect -11516 -13868 -11420 -13852
rect -10104 -13852 -10088 -13028
rect -10024 -13852 -10008 -13028
rect -8692 -13028 -8596 -13012
rect -9685 -13080 -8963 -13079
rect -9685 -13800 -9684 -13080
rect -8964 -13800 -8963 -13080
rect -9685 -13801 -8963 -13800
rect -10104 -13868 -10008 -13852
rect -8692 -13852 -8676 -13028
rect -8612 -13852 -8596 -13028
rect -7280 -13028 -7184 -13012
rect -8273 -13080 -7551 -13079
rect -8273 -13800 -8272 -13080
rect -7552 -13800 -7551 -13080
rect -8273 -13801 -7551 -13800
rect -8692 -13868 -8596 -13852
rect -7280 -13852 -7264 -13028
rect -7200 -13852 -7184 -13028
rect -5868 -13028 -5772 -13012
rect -6861 -13080 -6139 -13079
rect -6861 -13800 -6860 -13080
rect -6140 -13800 -6139 -13080
rect -6861 -13801 -6139 -13800
rect -7280 -13868 -7184 -13852
rect -5868 -13852 -5852 -13028
rect -5788 -13852 -5772 -13028
rect -4456 -13028 -4360 -13012
rect -5449 -13080 -4727 -13079
rect -5449 -13800 -5448 -13080
rect -4728 -13800 -4727 -13080
rect -5449 -13801 -4727 -13800
rect -5868 -13868 -5772 -13852
rect -4456 -13852 -4440 -13028
rect -4376 -13852 -4360 -13028
rect -3044 -13028 -2948 -13012
rect -4037 -13080 -3315 -13079
rect -4037 -13800 -4036 -13080
rect -3316 -13800 -3315 -13080
rect -4037 -13801 -3315 -13800
rect -4456 -13868 -4360 -13852
rect -3044 -13852 -3028 -13028
rect -2964 -13852 -2948 -13028
rect -1632 -13028 -1536 -13012
rect -2625 -13080 -1903 -13079
rect -2625 -13800 -2624 -13080
rect -1904 -13800 -1903 -13080
rect -2625 -13801 -1903 -13800
rect -3044 -13868 -2948 -13852
rect -1632 -13852 -1616 -13028
rect -1552 -13852 -1536 -13028
rect -220 -13028 -124 -13012
rect -1213 -13080 -491 -13079
rect -1213 -13800 -1212 -13080
rect -492 -13800 -491 -13080
rect -1213 -13801 -491 -13800
rect -1632 -13868 -1536 -13852
rect -220 -13852 -204 -13028
rect -140 -13852 -124 -13028
rect 1192 -13028 1288 -13012
rect 199 -13080 921 -13079
rect 199 -13800 200 -13080
rect 920 -13800 921 -13080
rect 199 -13801 921 -13800
rect -220 -13868 -124 -13852
rect 1192 -13852 1208 -13028
rect 1272 -13852 1288 -13028
rect 2604 -13028 2700 -13012
rect 1611 -13080 2333 -13079
rect 1611 -13800 1612 -13080
rect 2332 -13800 2333 -13080
rect 1611 -13801 2333 -13800
rect 1192 -13868 1288 -13852
rect 2604 -13852 2620 -13028
rect 2684 -13852 2700 -13028
rect 4016 -13028 4112 -13012
rect 3023 -13080 3745 -13079
rect 3023 -13800 3024 -13080
rect 3744 -13800 3745 -13080
rect 3023 -13801 3745 -13800
rect 2604 -13868 2700 -13852
rect 4016 -13852 4032 -13028
rect 4096 -13852 4112 -13028
rect 5428 -13028 5524 -13012
rect 4435 -13080 5157 -13079
rect 4435 -13800 4436 -13080
rect 5156 -13800 5157 -13080
rect 4435 -13801 5157 -13800
rect 4016 -13868 4112 -13852
rect 5428 -13852 5444 -13028
rect 5508 -13852 5524 -13028
rect 6840 -13028 6936 -13012
rect 5847 -13080 6569 -13079
rect 5847 -13800 5848 -13080
rect 6568 -13800 6569 -13080
rect 5847 -13801 6569 -13800
rect 5428 -13868 5524 -13852
rect 6840 -13852 6856 -13028
rect 6920 -13852 6936 -13028
rect 8252 -13028 8348 -13012
rect 7259 -13080 7981 -13079
rect 7259 -13800 7260 -13080
rect 7980 -13800 7981 -13080
rect 7259 -13801 7981 -13800
rect 6840 -13868 6936 -13852
rect 8252 -13852 8268 -13028
rect 8332 -13852 8348 -13028
rect 9664 -13028 9760 -13012
rect 8671 -13080 9393 -13079
rect 8671 -13800 8672 -13080
rect 9392 -13800 9393 -13080
rect 8671 -13801 9393 -13800
rect 8252 -13868 8348 -13852
rect 9664 -13852 9680 -13028
rect 9744 -13852 9760 -13028
rect 11076 -13028 11172 -13012
rect 10083 -13080 10805 -13079
rect 10083 -13800 10084 -13080
rect 10804 -13800 10805 -13080
rect 10083 -13801 10805 -13800
rect 9664 -13868 9760 -13852
rect 11076 -13852 11092 -13028
rect 11156 -13852 11172 -13028
rect 12488 -13028 12584 -13012
rect 11495 -13080 12217 -13079
rect 11495 -13800 11496 -13080
rect 12216 -13800 12217 -13080
rect 11495 -13801 12217 -13800
rect 11076 -13868 11172 -13852
rect 12488 -13852 12504 -13028
rect 12568 -13852 12584 -13028
rect 13900 -13028 13996 -13012
rect 12907 -13080 13629 -13079
rect 12907 -13800 12908 -13080
rect 13628 -13800 13629 -13080
rect 12907 -13801 13629 -13800
rect 12488 -13868 12584 -13852
rect 13900 -13852 13916 -13028
rect 13980 -13852 13996 -13028
rect 15312 -13028 15408 -13012
rect 14319 -13080 15041 -13079
rect 14319 -13800 14320 -13080
rect 15040 -13800 15041 -13080
rect 14319 -13801 15041 -13800
rect 13900 -13868 13996 -13852
rect 15312 -13852 15328 -13028
rect 15392 -13852 15408 -13028
rect 16724 -13028 16820 -13012
rect 15731 -13080 16453 -13079
rect 15731 -13800 15732 -13080
rect 16452 -13800 16453 -13080
rect 15731 -13801 16453 -13800
rect 15312 -13868 15408 -13852
rect 16724 -13852 16740 -13028
rect 16804 -13852 16820 -13028
rect 18136 -13028 18232 -13012
rect 17143 -13080 17865 -13079
rect 17143 -13800 17144 -13080
rect 17864 -13800 17865 -13080
rect 17143 -13801 17865 -13800
rect 16724 -13868 16820 -13852
rect 18136 -13852 18152 -13028
rect 18216 -13852 18232 -13028
rect 19548 -13028 19644 -13012
rect 18555 -13080 19277 -13079
rect 18555 -13800 18556 -13080
rect 19276 -13800 19277 -13080
rect 18555 -13801 19277 -13800
rect 18136 -13868 18232 -13852
rect 19548 -13852 19564 -13028
rect 19628 -13852 19644 -13028
rect 20960 -13028 21056 -13012
rect 19967 -13080 20689 -13079
rect 19967 -13800 19968 -13080
rect 20688 -13800 20689 -13080
rect 19967 -13801 20689 -13800
rect 19548 -13868 19644 -13852
rect 20960 -13852 20976 -13028
rect 21040 -13852 21056 -13028
rect 22372 -13028 22468 -13012
rect 21379 -13080 22101 -13079
rect 21379 -13800 21380 -13080
rect 22100 -13800 22101 -13080
rect 21379 -13801 22101 -13800
rect 20960 -13868 21056 -13852
rect 22372 -13852 22388 -13028
rect 22452 -13852 22468 -13028
rect 23784 -13028 23880 -13012
rect 22791 -13080 23513 -13079
rect 22791 -13800 22792 -13080
rect 23512 -13800 23513 -13080
rect 22791 -13801 23513 -13800
rect 22372 -13868 22468 -13852
rect 23784 -13852 23800 -13028
rect 23864 -13852 23880 -13028
rect 23784 -13868 23880 -13852
rect -22812 -14148 -22716 -14132
rect -23805 -14200 -23083 -14199
rect -23805 -14920 -23804 -14200
rect -23084 -14920 -23083 -14200
rect -23805 -14921 -23083 -14920
rect -22812 -14972 -22796 -14148
rect -22732 -14972 -22716 -14148
rect -21400 -14148 -21304 -14132
rect -22393 -14200 -21671 -14199
rect -22393 -14920 -22392 -14200
rect -21672 -14920 -21671 -14200
rect -22393 -14921 -21671 -14920
rect -22812 -14988 -22716 -14972
rect -21400 -14972 -21384 -14148
rect -21320 -14972 -21304 -14148
rect -19988 -14148 -19892 -14132
rect -20981 -14200 -20259 -14199
rect -20981 -14920 -20980 -14200
rect -20260 -14920 -20259 -14200
rect -20981 -14921 -20259 -14920
rect -21400 -14988 -21304 -14972
rect -19988 -14972 -19972 -14148
rect -19908 -14972 -19892 -14148
rect -18576 -14148 -18480 -14132
rect -19569 -14200 -18847 -14199
rect -19569 -14920 -19568 -14200
rect -18848 -14920 -18847 -14200
rect -19569 -14921 -18847 -14920
rect -19988 -14988 -19892 -14972
rect -18576 -14972 -18560 -14148
rect -18496 -14972 -18480 -14148
rect -17164 -14148 -17068 -14132
rect -18157 -14200 -17435 -14199
rect -18157 -14920 -18156 -14200
rect -17436 -14920 -17435 -14200
rect -18157 -14921 -17435 -14920
rect -18576 -14988 -18480 -14972
rect -17164 -14972 -17148 -14148
rect -17084 -14972 -17068 -14148
rect -15752 -14148 -15656 -14132
rect -16745 -14200 -16023 -14199
rect -16745 -14920 -16744 -14200
rect -16024 -14920 -16023 -14200
rect -16745 -14921 -16023 -14920
rect -17164 -14988 -17068 -14972
rect -15752 -14972 -15736 -14148
rect -15672 -14972 -15656 -14148
rect -14340 -14148 -14244 -14132
rect -15333 -14200 -14611 -14199
rect -15333 -14920 -15332 -14200
rect -14612 -14920 -14611 -14200
rect -15333 -14921 -14611 -14920
rect -15752 -14988 -15656 -14972
rect -14340 -14972 -14324 -14148
rect -14260 -14972 -14244 -14148
rect -12928 -14148 -12832 -14132
rect -13921 -14200 -13199 -14199
rect -13921 -14920 -13920 -14200
rect -13200 -14920 -13199 -14200
rect -13921 -14921 -13199 -14920
rect -14340 -14988 -14244 -14972
rect -12928 -14972 -12912 -14148
rect -12848 -14972 -12832 -14148
rect -11516 -14148 -11420 -14132
rect -12509 -14200 -11787 -14199
rect -12509 -14920 -12508 -14200
rect -11788 -14920 -11787 -14200
rect -12509 -14921 -11787 -14920
rect -12928 -14988 -12832 -14972
rect -11516 -14972 -11500 -14148
rect -11436 -14972 -11420 -14148
rect -10104 -14148 -10008 -14132
rect -11097 -14200 -10375 -14199
rect -11097 -14920 -11096 -14200
rect -10376 -14920 -10375 -14200
rect -11097 -14921 -10375 -14920
rect -11516 -14988 -11420 -14972
rect -10104 -14972 -10088 -14148
rect -10024 -14972 -10008 -14148
rect -8692 -14148 -8596 -14132
rect -9685 -14200 -8963 -14199
rect -9685 -14920 -9684 -14200
rect -8964 -14920 -8963 -14200
rect -9685 -14921 -8963 -14920
rect -10104 -14988 -10008 -14972
rect -8692 -14972 -8676 -14148
rect -8612 -14972 -8596 -14148
rect -7280 -14148 -7184 -14132
rect -8273 -14200 -7551 -14199
rect -8273 -14920 -8272 -14200
rect -7552 -14920 -7551 -14200
rect -8273 -14921 -7551 -14920
rect -8692 -14988 -8596 -14972
rect -7280 -14972 -7264 -14148
rect -7200 -14972 -7184 -14148
rect -5868 -14148 -5772 -14132
rect -6861 -14200 -6139 -14199
rect -6861 -14920 -6860 -14200
rect -6140 -14920 -6139 -14200
rect -6861 -14921 -6139 -14920
rect -7280 -14988 -7184 -14972
rect -5868 -14972 -5852 -14148
rect -5788 -14972 -5772 -14148
rect -4456 -14148 -4360 -14132
rect -5449 -14200 -4727 -14199
rect -5449 -14920 -5448 -14200
rect -4728 -14920 -4727 -14200
rect -5449 -14921 -4727 -14920
rect -5868 -14988 -5772 -14972
rect -4456 -14972 -4440 -14148
rect -4376 -14972 -4360 -14148
rect -3044 -14148 -2948 -14132
rect -4037 -14200 -3315 -14199
rect -4037 -14920 -4036 -14200
rect -3316 -14920 -3315 -14200
rect -4037 -14921 -3315 -14920
rect -4456 -14988 -4360 -14972
rect -3044 -14972 -3028 -14148
rect -2964 -14972 -2948 -14148
rect -1632 -14148 -1536 -14132
rect -2625 -14200 -1903 -14199
rect -2625 -14920 -2624 -14200
rect -1904 -14920 -1903 -14200
rect -2625 -14921 -1903 -14920
rect -3044 -14988 -2948 -14972
rect -1632 -14972 -1616 -14148
rect -1552 -14972 -1536 -14148
rect -220 -14148 -124 -14132
rect -1213 -14200 -491 -14199
rect -1213 -14920 -1212 -14200
rect -492 -14920 -491 -14200
rect -1213 -14921 -491 -14920
rect -1632 -14988 -1536 -14972
rect -220 -14972 -204 -14148
rect -140 -14972 -124 -14148
rect 1192 -14148 1288 -14132
rect 199 -14200 921 -14199
rect 199 -14920 200 -14200
rect 920 -14920 921 -14200
rect 199 -14921 921 -14920
rect -220 -14988 -124 -14972
rect 1192 -14972 1208 -14148
rect 1272 -14972 1288 -14148
rect 2604 -14148 2700 -14132
rect 1611 -14200 2333 -14199
rect 1611 -14920 1612 -14200
rect 2332 -14920 2333 -14200
rect 1611 -14921 2333 -14920
rect 1192 -14988 1288 -14972
rect 2604 -14972 2620 -14148
rect 2684 -14972 2700 -14148
rect 4016 -14148 4112 -14132
rect 3023 -14200 3745 -14199
rect 3023 -14920 3024 -14200
rect 3744 -14920 3745 -14200
rect 3023 -14921 3745 -14920
rect 2604 -14988 2700 -14972
rect 4016 -14972 4032 -14148
rect 4096 -14972 4112 -14148
rect 5428 -14148 5524 -14132
rect 4435 -14200 5157 -14199
rect 4435 -14920 4436 -14200
rect 5156 -14920 5157 -14200
rect 4435 -14921 5157 -14920
rect 4016 -14988 4112 -14972
rect 5428 -14972 5444 -14148
rect 5508 -14972 5524 -14148
rect 6840 -14148 6936 -14132
rect 5847 -14200 6569 -14199
rect 5847 -14920 5848 -14200
rect 6568 -14920 6569 -14200
rect 5847 -14921 6569 -14920
rect 5428 -14988 5524 -14972
rect 6840 -14972 6856 -14148
rect 6920 -14972 6936 -14148
rect 8252 -14148 8348 -14132
rect 7259 -14200 7981 -14199
rect 7259 -14920 7260 -14200
rect 7980 -14920 7981 -14200
rect 7259 -14921 7981 -14920
rect 6840 -14988 6936 -14972
rect 8252 -14972 8268 -14148
rect 8332 -14972 8348 -14148
rect 9664 -14148 9760 -14132
rect 8671 -14200 9393 -14199
rect 8671 -14920 8672 -14200
rect 9392 -14920 9393 -14200
rect 8671 -14921 9393 -14920
rect 8252 -14988 8348 -14972
rect 9664 -14972 9680 -14148
rect 9744 -14972 9760 -14148
rect 11076 -14148 11172 -14132
rect 10083 -14200 10805 -14199
rect 10083 -14920 10084 -14200
rect 10804 -14920 10805 -14200
rect 10083 -14921 10805 -14920
rect 9664 -14988 9760 -14972
rect 11076 -14972 11092 -14148
rect 11156 -14972 11172 -14148
rect 12488 -14148 12584 -14132
rect 11495 -14200 12217 -14199
rect 11495 -14920 11496 -14200
rect 12216 -14920 12217 -14200
rect 11495 -14921 12217 -14920
rect 11076 -14988 11172 -14972
rect 12488 -14972 12504 -14148
rect 12568 -14972 12584 -14148
rect 13900 -14148 13996 -14132
rect 12907 -14200 13629 -14199
rect 12907 -14920 12908 -14200
rect 13628 -14920 13629 -14200
rect 12907 -14921 13629 -14920
rect 12488 -14988 12584 -14972
rect 13900 -14972 13916 -14148
rect 13980 -14972 13996 -14148
rect 15312 -14148 15408 -14132
rect 14319 -14200 15041 -14199
rect 14319 -14920 14320 -14200
rect 15040 -14920 15041 -14200
rect 14319 -14921 15041 -14920
rect 13900 -14988 13996 -14972
rect 15312 -14972 15328 -14148
rect 15392 -14972 15408 -14148
rect 16724 -14148 16820 -14132
rect 15731 -14200 16453 -14199
rect 15731 -14920 15732 -14200
rect 16452 -14920 16453 -14200
rect 15731 -14921 16453 -14920
rect 15312 -14988 15408 -14972
rect 16724 -14972 16740 -14148
rect 16804 -14972 16820 -14148
rect 18136 -14148 18232 -14132
rect 17143 -14200 17865 -14199
rect 17143 -14920 17144 -14200
rect 17864 -14920 17865 -14200
rect 17143 -14921 17865 -14920
rect 16724 -14988 16820 -14972
rect 18136 -14972 18152 -14148
rect 18216 -14972 18232 -14148
rect 19548 -14148 19644 -14132
rect 18555 -14200 19277 -14199
rect 18555 -14920 18556 -14200
rect 19276 -14920 19277 -14200
rect 18555 -14921 19277 -14920
rect 18136 -14988 18232 -14972
rect 19548 -14972 19564 -14148
rect 19628 -14972 19644 -14148
rect 20960 -14148 21056 -14132
rect 19967 -14200 20689 -14199
rect 19967 -14920 19968 -14200
rect 20688 -14920 20689 -14200
rect 19967 -14921 20689 -14920
rect 19548 -14988 19644 -14972
rect 20960 -14972 20976 -14148
rect 21040 -14972 21056 -14148
rect 22372 -14148 22468 -14132
rect 21379 -14200 22101 -14199
rect 21379 -14920 21380 -14200
rect 22100 -14920 22101 -14200
rect 21379 -14921 22101 -14920
rect 20960 -14988 21056 -14972
rect 22372 -14972 22388 -14148
rect 22452 -14972 22468 -14148
rect 23784 -14148 23880 -14132
rect 22791 -14200 23513 -14199
rect 22791 -14920 22792 -14200
rect 23512 -14920 23513 -14200
rect 22791 -14921 23513 -14920
rect 22372 -14988 22468 -14972
rect 23784 -14972 23800 -14148
rect 23864 -14972 23880 -14148
rect 23784 -14988 23880 -14972
rect -22812 -15268 -22716 -15252
rect -23805 -15320 -23083 -15319
rect -23805 -16040 -23804 -15320
rect -23084 -16040 -23083 -15320
rect -23805 -16041 -23083 -16040
rect -22812 -16092 -22796 -15268
rect -22732 -16092 -22716 -15268
rect -21400 -15268 -21304 -15252
rect -22393 -15320 -21671 -15319
rect -22393 -16040 -22392 -15320
rect -21672 -16040 -21671 -15320
rect -22393 -16041 -21671 -16040
rect -22812 -16108 -22716 -16092
rect -21400 -16092 -21384 -15268
rect -21320 -16092 -21304 -15268
rect -19988 -15268 -19892 -15252
rect -20981 -15320 -20259 -15319
rect -20981 -16040 -20980 -15320
rect -20260 -16040 -20259 -15320
rect -20981 -16041 -20259 -16040
rect -21400 -16108 -21304 -16092
rect -19988 -16092 -19972 -15268
rect -19908 -16092 -19892 -15268
rect -18576 -15268 -18480 -15252
rect -19569 -15320 -18847 -15319
rect -19569 -16040 -19568 -15320
rect -18848 -16040 -18847 -15320
rect -19569 -16041 -18847 -16040
rect -19988 -16108 -19892 -16092
rect -18576 -16092 -18560 -15268
rect -18496 -16092 -18480 -15268
rect -17164 -15268 -17068 -15252
rect -18157 -15320 -17435 -15319
rect -18157 -16040 -18156 -15320
rect -17436 -16040 -17435 -15320
rect -18157 -16041 -17435 -16040
rect -18576 -16108 -18480 -16092
rect -17164 -16092 -17148 -15268
rect -17084 -16092 -17068 -15268
rect -15752 -15268 -15656 -15252
rect -16745 -15320 -16023 -15319
rect -16745 -16040 -16744 -15320
rect -16024 -16040 -16023 -15320
rect -16745 -16041 -16023 -16040
rect -17164 -16108 -17068 -16092
rect -15752 -16092 -15736 -15268
rect -15672 -16092 -15656 -15268
rect -14340 -15268 -14244 -15252
rect -15333 -15320 -14611 -15319
rect -15333 -16040 -15332 -15320
rect -14612 -16040 -14611 -15320
rect -15333 -16041 -14611 -16040
rect -15752 -16108 -15656 -16092
rect -14340 -16092 -14324 -15268
rect -14260 -16092 -14244 -15268
rect -12928 -15268 -12832 -15252
rect -13921 -15320 -13199 -15319
rect -13921 -16040 -13920 -15320
rect -13200 -16040 -13199 -15320
rect -13921 -16041 -13199 -16040
rect -14340 -16108 -14244 -16092
rect -12928 -16092 -12912 -15268
rect -12848 -16092 -12832 -15268
rect -11516 -15268 -11420 -15252
rect -12509 -15320 -11787 -15319
rect -12509 -16040 -12508 -15320
rect -11788 -16040 -11787 -15320
rect -12509 -16041 -11787 -16040
rect -12928 -16108 -12832 -16092
rect -11516 -16092 -11500 -15268
rect -11436 -16092 -11420 -15268
rect -10104 -15268 -10008 -15252
rect -11097 -15320 -10375 -15319
rect -11097 -16040 -11096 -15320
rect -10376 -16040 -10375 -15320
rect -11097 -16041 -10375 -16040
rect -11516 -16108 -11420 -16092
rect -10104 -16092 -10088 -15268
rect -10024 -16092 -10008 -15268
rect -8692 -15268 -8596 -15252
rect -9685 -15320 -8963 -15319
rect -9685 -16040 -9684 -15320
rect -8964 -16040 -8963 -15320
rect -9685 -16041 -8963 -16040
rect -10104 -16108 -10008 -16092
rect -8692 -16092 -8676 -15268
rect -8612 -16092 -8596 -15268
rect -7280 -15268 -7184 -15252
rect -8273 -15320 -7551 -15319
rect -8273 -16040 -8272 -15320
rect -7552 -16040 -7551 -15320
rect -8273 -16041 -7551 -16040
rect -8692 -16108 -8596 -16092
rect -7280 -16092 -7264 -15268
rect -7200 -16092 -7184 -15268
rect -5868 -15268 -5772 -15252
rect -6861 -15320 -6139 -15319
rect -6861 -16040 -6860 -15320
rect -6140 -16040 -6139 -15320
rect -6861 -16041 -6139 -16040
rect -7280 -16108 -7184 -16092
rect -5868 -16092 -5852 -15268
rect -5788 -16092 -5772 -15268
rect -4456 -15268 -4360 -15252
rect -5449 -15320 -4727 -15319
rect -5449 -16040 -5448 -15320
rect -4728 -16040 -4727 -15320
rect -5449 -16041 -4727 -16040
rect -5868 -16108 -5772 -16092
rect -4456 -16092 -4440 -15268
rect -4376 -16092 -4360 -15268
rect -3044 -15268 -2948 -15252
rect -4037 -15320 -3315 -15319
rect -4037 -16040 -4036 -15320
rect -3316 -16040 -3315 -15320
rect -4037 -16041 -3315 -16040
rect -4456 -16108 -4360 -16092
rect -3044 -16092 -3028 -15268
rect -2964 -16092 -2948 -15268
rect -1632 -15268 -1536 -15252
rect -2625 -15320 -1903 -15319
rect -2625 -16040 -2624 -15320
rect -1904 -16040 -1903 -15320
rect -2625 -16041 -1903 -16040
rect -3044 -16108 -2948 -16092
rect -1632 -16092 -1616 -15268
rect -1552 -16092 -1536 -15268
rect -220 -15268 -124 -15252
rect -1213 -15320 -491 -15319
rect -1213 -16040 -1212 -15320
rect -492 -16040 -491 -15320
rect -1213 -16041 -491 -16040
rect -1632 -16108 -1536 -16092
rect -220 -16092 -204 -15268
rect -140 -16092 -124 -15268
rect 1192 -15268 1288 -15252
rect 199 -15320 921 -15319
rect 199 -16040 200 -15320
rect 920 -16040 921 -15320
rect 199 -16041 921 -16040
rect -220 -16108 -124 -16092
rect 1192 -16092 1208 -15268
rect 1272 -16092 1288 -15268
rect 2604 -15268 2700 -15252
rect 1611 -15320 2333 -15319
rect 1611 -16040 1612 -15320
rect 2332 -16040 2333 -15320
rect 1611 -16041 2333 -16040
rect 1192 -16108 1288 -16092
rect 2604 -16092 2620 -15268
rect 2684 -16092 2700 -15268
rect 4016 -15268 4112 -15252
rect 3023 -15320 3745 -15319
rect 3023 -16040 3024 -15320
rect 3744 -16040 3745 -15320
rect 3023 -16041 3745 -16040
rect 2604 -16108 2700 -16092
rect 4016 -16092 4032 -15268
rect 4096 -16092 4112 -15268
rect 5428 -15268 5524 -15252
rect 4435 -15320 5157 -15319
rect 4435 -16040 4436 -15320
rect 5156 -16040 5157 -15320
rect 4435 -16041 5157 -16040
rect 4016 -16108 4112 -16092
rect 5428 -16092 5444 -15268
rect 5508 -16092 5524 -15268
rect 6840 -15268 6936 -15252
rect 5847 -15320 6569 -15319
rect 5847 -16040 5848 -15320
rect 6568 -16040 6569 -15320
rect 5847 -16041 6569 -16040
rect 5428 -16108 5524 -16092
rect 6840 -16092 6856 -15268
rect 6920 -16092 6936 -15268
rect 8252 -15268 8348 -15252
rect 7259 -15320 7981 -15319
rect 7259 -16040 7260 -15320
rect 7980 -16040 7981 -15320
rect 7259 -16041 7981 -16040
rect 6840 -16108 6936 -16092
rect 8252 -16092 8268 -15268
rect 8332 -16092 8348 -15268
rect 9664 -15268 9760 -15252
rect 8671 -15320 9393 -15319
rect 8671 -16040 8672 -15320
rect 9392 -16040 9393 -15320
rect 8671 -16041 9393 -16040
rect 8252 -16108 8348 -16092
rect 9664 -16092 9680 -15268
rect 9744 -16092 9760 -15268
rect 11076 -15268 11172 -15252
rect 10083 -15320 10805 -15319
rect 10083 -16040 10084 -15320
rect 10804 -16040 10805 -15320
rect 10083 -16041 10805 -16040
rect 9664 -16108 9760 -16092
rect 11076 -16092 11092 -15268
rect 11156 -16092 11172 -15268
rect 12488 -15268 12584 -15252
rect 11495 -15320 12217 -15319
rect 11495 -16040 11496 -15320
rect 12216 -16040 12217 -15320
rect 11495 -16041 12217 -16040
rect 11076 -16108 11172 -16092
rect 12488 -16092 12504 -15268
rect 12568 -16092 12584 -15268
rect 13900 -15268 13996 -15252
rect 12907 -15320 13629 -15319
rect 12907 -16040 12908 -15320
rect 13628 -16040 13629 -15320
rect 12907 -16041 13629 -16040
rect 12488 -16108 12584 -16092
rect 13900 -16092 13916 -15268
rect 13980 -16092 13996 -15268
rect 15312 -15268 15408 -15252
rect 14319 -15320 15041 -15319
rect 14319 -16040 14320 -15320
rect 15040 -16040 15041 -15320
rect 14319 -16041 15041 -16040
rect 13900 -16108 13996 -16092
rect 15312 -16092 15328 -15268
rect 15392 -16092 15408 -15268
rect 16724 -15268 16820 -15252
rect 15731 -15320 16453 -15319
rect 15731 -16040 15732 -15320
rect 16452 -16040 16453 -15320
rect 15731 -16041 16453 -16040
rect 15312 -16108 15408 -16092
rect 16724 -16092 16740 -15268
rect 16804 -16092 16820 -15268
rect 18136 -15268 18232 -15252
rect 17143 -15320 17865 -15319
rect 17143 -16040 17144 -15320
rect 17864 -16040 17865 -15320
rect 17143 -16041 17865 -16040
rect 16724 -16108 16820 -16092
rect 18136 -16092 18152 -15268
rect 18216 -16092 18232 -15268
rect 19548 -15268 19644 -15252
rect 18555 -15320 19277 -15319
rect 18555 -16040 18556 -15320
rect 19276 -16040 19277 -15320
rect 18555 -16041 19277 -16040
rect 18136 -16108 18232 -16092
rect 19548 -16092 19564 -15268
rect 19628 -16092 19644 -15268
rect 20960 -15268 21056 -15252
rect 19967 -15320 20689 -15319
rect 19967 -16040 19968 -15320
rect 20688 -16040 20689 -15320
rect 19967 -16041 20689 -16040
rect 19548 -16108 19644 -16092
rect 20960 -16092 20976 -15268
rect 21040 -16092 21056 -15268
rect 22372 -15268 22468 -15252
rect 21379 -15320 22101 -15319
rect 21379 -16040 21380 -15320
rect 22100 -16040 22101 -15320
rect 21379 -16041 22101 -16040
rect 20960 -16108 21056 -16092
rect 22372 -16092 22388 -15268
rect 22452 -16092 22468 -15268
rect 23784 -15268 23880 -15252
rect 22791 -15320 23513 -15319
rect 22791 -16040 22792 -15320
rect 23512 -16040 23513 -15320
rect 22791 -16041 23513 -16040
rect 22372 -16108 22468 -16092
rect 23784 -16092 23800 -15268
rect 23864 -16092 23880 -15268
rect 23784 -16108 23880 -16092
rect -22812 -16388 -22716 -16372
rect -23805 -16440 -23083 -16439
rect -23805 -17160 -23804 -16440
rect -23084 -17160 -23083 -16440
rect -23805 -17161 -23083 -17160
rect -22812 -17212 -22796 -16388
rect -22732 -17212 -22716 -16388
rect -21400 -16388 -21304 -16372
rect -22393 -16440 -21671 -16439
rect -22393 -17160 -22392 -16440
rect -21672 -17160 -21671 -16440
rect -22393 -17161 -21671 -17160
rect -22812 -17228 -22716 -17212
rect -21400 -17212 -21384 -16388
rect -21320 -17212 -21304 -16388
rect -19988 -16388 -19892 -16372
rect -20981 -16440 -20259 -16439
rect -20981 -17160 -20980 -16440
rect -20260 -17160 -20259 -16440
rect -20981 -17161 -20259 -17160
rect -21400 -17228 -21304 -17212
rect -19988 -17212 -19972 -16388
rect -19908 -17212 -19892 -16388
rect -18576 -16388 -18480 -16372
rect -19569 -16440 -18847 -16439
rect -19569 -17160 -19568 -16440
rect -18848 -17160 -18847 -16440
rect -19569 -17161 -18847 -17160
rect -19988 -17228 -19892 -17212
rect -18576 -17212 -18560 -16388
rect -18496 -17212 -18480 -16388
rect -17164 -16388 -17068 -16372
rect -18157 -16440 -17435 -16439
rect -18157 -17160 -18156 -16440
rect -17436 -17160 -17435 -16440
rect -18157 -17161 -17435 -17160
rect -18576 -17228 -18480 -17212
rect -17164 -17212 -17148 -16388
rect -17084 -17212 -17068 -16388
rect -15752 -16388 -15656 -16372
rect -16745 -16440 -16023 -16439
rect -16745 -17160 -16744 -16440
rect -16024 -17160 -16023 -16440
rect -16745 -17161 -16023 -17160
rect -17164 -17228 -17068 -17212
rect -15752 -17212 -15736 -16388
rect -15672 -17212 -15656 -16388
rect -14340 -16388 -14244 -16372
rect -15333 -16440 -14611 -16439
rect -15333 -17160 -15332 -16440
rect -14612 -17160 -14611 -16440
rect -15333 -17161 -14611 -17160
rect -15752 -17228 -15656 -17212
rect -14340 -17212 -14324 -16388
rect -14260 -17212 -14244 -16388
rect -12928 -16388 -12832 -16372
rect -13921 -16440 -13199 -16439
rect -13921 -17160 -13920 -16440
rect -13200 -17160 -13199 -16440
rect -13921 -17161 -13199 -17160
rect -14340 -17228 -14244 -17212
rect -12928 -17212 -12912 -16388
rect -12848 -17212 -12832 -16388
rect -11516 -16388 -11420 -16372
rect -12509 -16440 -11787 -16439
rect -12509 -17160 -12508 -16440
rect -11788 -17160 -11787 -16440
rect -12509 -17161 -11787 -17160
rect -12928 -17228 -12832 -17212
rect -11516 -17212 -11500 -16388
rect -11436 -17212 -11420 -16388
rect -10104 -16388 -10008 -16372
rect -11097 -16440 -10375 -16439
rect -11097 -17160 -11096 -16440
rect -10376 -17160 -10375 -16440
rect -11097 -17161 -10375 -17160
rect -11516 -17228 -11420 -17212
rect -10104 -17212 -10088 -16388
rect -10024 -17212 -10008 -16388
rect -8692 -16388 -8596 -16372
rect -9685 -16440 -8963 -16439
rect -9685 -17160 -9684 -16440
rect -8964 -17160 -8963 -16440
rect -9685 -17161 -8963 -17160
rect -10104 -17228 -10008 -17212
rect -8692 -17212 -8676 -16388
rect -8612 -17212 -8596 -16388
rect -7280 -16388 -7184 -16372
rect -8273 -16440 -7551 -16439
rect -8273 -17160 -8272 -16440
rect -7552 -17160 -7551 -16440
rect -8273 -17161 -7551 -17160
rect -8692 -17228 -8596 -17212
rect -7280 -17212 -7264 -16388
rect -7200 -17212 -7184 -16388
rect -5868 -16388 -5772 -16372
rect -6861 -16440 -6139 -16439
rect -6861 -17160 -6860 -16440
rect -6140 -17160 -6139 -16440
rect -6861 -17161 -6139 -17160
rect -7280 -17228 -7184 -17212
rect -5868 -17212 -5852 -16388
rect -5788 -17212 -5772 -16388
rect -4456 -16388 -4360 -16372
rect -5449 -16440 -4727 -16439
rect -5449 -17160 -5448 -16440
rect -4728 -17160 -4727 -16440
rect -5449 -17161 -4727 -17160
rect -5868 -17228 -5772 -17212
rect -4456 -17212 -4440 -16388
rect -4376 -17212 -4360 -16388
rect -3044 -16388 -2948 -16372
rect -4037 -16440 -3315 -16439
rect -4037 -17160 -4036 -16440
rect -3316 -17160 -3315 -16440
rect -4037 -17161 -3315 -17160
rect -4456 -17228 -4360 -17212
rect -3044 -17212 -3028 -16388
rect -2964 -17212 -2948 -16388
rect -1632 -16388 -1536 -16372
rect -2625 -16440 -1903 -16439
rect -2625 -17160 -2624 -16440
rect -1904 -17160 -1903 -16440
rect -2625 -17161 -1903 -17160
rect -3044 -17228 -2948 -17212
rect -1632 -17212 -1616 -16388
rect -1552 -17212 -1536 -16388
rect -220 -16388 -124 -16372
rect -1213 -16440 -491 -16439
rect -1213 -17160 -1212 -16440
rect -492 -17160 -491 -16440
rect -1213 -17161 -491 -17160
rect -1632 -17228 -1536 -17212
rect -220 -17212 -204 -16388
rect -140 -17212 -124 -16388
rect 1192 -16388 1288 -16372
rect 199 -16440 921 -16439
rect 199 -17160 200 -16440
rect 920 -17160 921 -16440
rect 199 -17161 921 -17160
rect -220 -17228 -124 -17212
rect 1192 -17212 1208 -16388
rect 1272 -17212 1288 -16388
rect 2604 -16388 2700 -16372
rect 1611 -16440 2333 -16439
rect 1611 -17160 1612 -16440
rect 2332 -17160 2333 -16440
rect 1611 -17161 2333 -17160
rect 1192 -17228 1288 -17212
rect 2604 -17212 2620 -16388
rect 2684 -17212 2700 -16388
rect 4016 -16388 4112 -16372
rect 3023 -16440 3745 -16439
rect 3023 -17160 3024 -16440
rect 3744 -17160 3745 -16440
rect 3023 -17161 3745 -17160
rect 2604 -17228 2700 -17212
rect 4016 -17212 4032 -16388
rect 4096 -17212 4112 -16388
rect 5428 -16388 5524 -16372
rect 4435 -16440 5157 -16439
rect 4435 -17160 4436 -16440
rect 5156 -17160 5157 -16440
rect 4435 -17161 5157 -17160
rect 4016 -17228 4112 -17212
rect 5428 -17212 5444 -16388
rect 5508 -17212 5524 -16388
rect 6840 -16388 6936 -16372
rect 5847 -16440 6569 -16439
rect 5847 -17160 5848 -16440
rect 6568 -17160 6569 -16440
rect 5847 -17161 6569 -17160
rect 5428 -17228 5524 -17212
rect 6840 -17212 6856 -16388
rect 6920 -17212 6936 -16388
rect 8252 -16388 8348 -16372
rect 7259 -16440 7981 -16439
rect 7259 -17160 7260 -16440
rect 7980 -17160 7981 -16440
rect 7259 -17161 7981 -17160
rect 6840 -17228 6936 -17212
rect 8252 -17212 8268 -16388
rect 8332 -17212 8348 -16388
rect 9664 -16388 9760 -16372
rect 8671 -16440 9393 -16439
rect 8671 -17160 8672 -16440
rect 9392 -17160 9393 -16440
rect 8671 -17161 9393 -17160
rect 8252 -17228 8348 -17212
rect 9664 -17212 9680 -16388
rect 9744 -17212 9760 -16388
rect 11076 -16388 11172 -16372
rect 10083 -16440 10805 -16439
rect 10083 -17160 10084 -16440
rect 10804 -17160 10805 -16440
rect 10083 -17161 10805 -17160
rect 9664 -17228 9760 -17212
rect 11076 -17212 11092 -16388
rect 11156 -17212 11172 -16388
rect 12488 -16388 12584 -16372
rect 11495 -16440 12217 -16439
rect 11495 -17160 11496 -16440
rect 12216 -17160 12217 -16440
rect 11495 -17161 12217 -17160
rect 11076 -17228 11172 -17212
rect 12488 -17212 12504 -16388
rect 12568 -17212 12584 -16388
rect 13900 -16388 13996 -16372
rect 12907 -16440 13629 -16439
rect 12907 -17160 12908 -16440
rect 13628 -17160 13629 -16440
rect 12907 -17161 13629 -17160
rect 12488 -17228 12584 -17212
rect 13900 -17212 13916 -16388
rect 13980 -17212 13996 -16388
rect 15312 -16388 15408 -16372
rect 14319 -16440 15041 -16439
rect 14319 -17160 14320 -16440
rect 15040 -17160 15041 -16440
rect 14319 -17161 15041 -17160
rect 13900 -17228 13996 -17212
rect 15312 -17212 15328 -16388
rect 15392 -17212 15408 -16388
rect 16724 -16388 16820 -16372
rect 15731 -16440 16453 -16439
rect 15731 -17160 15732 -16440
rect 16452 -17160 16453 -16440
rect 15731 -17161 16453 -17160
rect 15312 -17228 15408 -17212
rect 16724 -17212 16740 -16388
rect 16804 -17212 16820 -16388
rect 18136 -16388 18232 -16372
rect 17143 -16440 17865 -16439
rect 17143 -17160 17144 -16440
rect 17864 -17160 17865 -16440
rect 17143 -17161 17865 -17160
rect 16724 -17228 16820 -17212
rect 18136 -17212 18152 -16388
rect 18216 -17212 18232 -16388
rect 19548 -16388 19644 -16372
rect 18555 -16440 19277 -16439
rect 18555 -17160 18556 -16440
rect 19276 -17160 19277 -16440
rect 18555 -17161 19277 -17160
rect 18136 -17228 18232 -17212
rect 19548 -17212 19564 -16388
rect 19628 -17212 19644 -16388
rect 20960 -16388 21056 -16372
rect 19967 -16440 20689 -16439
rect 19967 -17160 19968 -16440
rect 20688 -17160 20689 -16440
rect 19967 -17161 20689 -17160
rect 19548 -17228 19644 -17212
rect 20960 -17212 20976 -16388
rect 21040 -17212 21056 -16388
rect 22372 -16388 22468 -16372
rect 21379 -16440 22101 -16439
rect 21379 -17160 21380 -16440
rect 22100 -17160 22101 -16440
rect 21379 -17161 22101 -17160
rect 20960 -17228 21056 -17212
rect 22372 -17212 22388 -16388
rect 22452 -17212 22468 -16388
rect 23784 -16388 23880 -16372
rect 22791 -16440 23513 -16439
rect 22791 -17160 22792 -16440
rect 23512 -17160 23513 -16440
rect 22791 -17161 23513 -17160
rect 22372 -17228 22468 -17212
rect 23784 -17212 23800 -16388
rect 23864 -17212 23880 -16388
rect 23784 -17228 23880 -17212
rect -22812 -17508 -22716 -17492
rect -23805 -17560 -23083 -17559
rect -23805 -18280 -23804 -17560
rect -23084 -18280 -23083 -17560
rect -23805 -18281 -23083 -18280
rect -22812 -18332 -22796 -17508
rect -22732 -18332 -22716 -17508
rect -21400 -17508 -21304 -17492
rect -22393 -17560 -21671 -17559
rect -22393 -18280 -22392 -17560
rect -21672 -18280 -21671 -17560
rect -22393 -18281 -21671 -18280
rect -22812 -18348 -22716 -18332
rect -21400 -18332 -21384 -17508
rect -21320 -18332 -21304 -17508
rect -19988 -17508 -19892 -17492
rect -20981 -17560 -20259 -17559
rect -20981 -18280 -20980 -17560
rect -20260 -18280 -20259 -17560
rect -20981 -18281 -20259 -18280
rect -21400 -18348 -21304 -18332
rect -19988 -18332 -19972 -17508
rect -19908 -18332 -19892 -17508
rect -18576 -17508 -18480 -17492
rect -19569 -17560 -18847 -17559
rect -19569 -18280 -19568 -17560
rect -18848 -18280 -18847 -17560
rect -19569 -18281 -18847 -18280
rect -19988 -18348 -19892 -18332
rect -18576 -18332 -18560 -17508
rect -18496 -18332 -18480 -17508
rect -17164 -17508 -17068 -17492
rect -18157 -17560 -17435 -17559
rect -18157 -18280 -18156 -17560
rect -17436 -18280 -17435 -17560
rect -18157 -18281 -17435 -18280
rect -18576 -18348 -18480 -18332
rect -17164 -18332 -17148 -17508
rect -17084 -18332 -17068 -17508
rect -15752 -17508 -15656 -17492
rect -16745 -17560 -16023 -17559
rect -16745 -18280 -16744 -17560
rect -16024 -18280 -16023 -17560
rect -16745 -18281 -16023 -18280
rect -17164 -18348 -17068 -18332
rect -15752 -18332 -15736 -17508
rect -15672 -18332 -15656 -17508
rect -14340 -17508 -14244 -17492
rect -15333 -17560 -14611 -17559
rect -15333 -18280 -15332 -17560
rect -14612 -18280 -14611 -17560
rect -15333 -18281 -14611 -18280
rect -15752 -18348 -15656 -18332
rect -14340 -18332 -14324 -17508
rect -14260 -18332 -14244 -17508
rect -12928 -17508 -12832 -17492
rect -13921 -17560 -13199 -17559
rect -13921 -18280 -13920 -17560
rect -13200 -18280 -13199 -17560
rect -13921 -18281 -13199 -18280
rect -14340 -18348 -14244 -18332
rect -12928 -18332 -12912 -17508
rect -12848 -18332 -12832 -17508
rect -11516 -17508 -11420 -17492
rect -12509 -17560 -11787 -17559
rect -12509 -18280 -12508 -17560
rect -11788 -18280 -11787 -17560
rect -12509 -18281 -11787 -18280
rect -12928 -18348 -12832 -18332
rect -11516 -18332 -11500 -17508
rect -11436 -18332 -11420 -17508
rect -10104 -17508 -10008 -17492
rect -11097 -17560 -10375 -17559
rect -11097 -18280 -11096 -17560
rect -10376 -18280 -10375 -17560
rect -11097 -18281 -10375 -18280
rect -11516 -18348 -11420 -18332
rect -10104 -18332 -10088 -17508
rect -10024 -18332 -10008 -17508
rect -8692 -17508 -8596 -17492
rect -9685 -17560 -8963 -17559
rect -9685 -18280 -9684 -17560
rect -8964 -18280 -8963 -17560
rect -9685 -18281 -8963 -18280
rect -10104 -18348 -10008 -18332
rect -8692 -18332 -8676 -17508
rect -8612 -18332 -8596 -17508
rect -7280 -17508 -7184 -17492
rect -8273 -17560 -7551 -17559
rect -8273 -18280 -8272 -17560
rect -7552 -18280 -7551 -17560
rect -8273 -18281 -7551 -18280
rect -8692 -18348 -8596 -18332
rect -7280 -18332 -7264 -17508
rect -7200 -18332 -7184 -17508
rect -5868 -17508 -5772 -17492
rect -6861 -17560 -6139 -17559
rect -6861 -18280 -6860 -17560
rect -6140 -18280 -6139 -17560
rect -6861 -18281 -6139 -18280
rect -7280 -18348 -7184 -18332
rect -5868 -18332 -5852 -17508
rect -5788 -18332 -5772 -17508
rect -4456 -17508 -4360 -17492
rect -5449 -17560 -4727 -17559
rect -5449 -18280 -5448 -17560
rect -4728 -18280 -4727 -17560
rect -5449 -18281 -4727 -18280
rect -5868 -18348 -5772 -18332
rect -4456 -18332 -4440 -17508
rect -4376 -18332 -4360 -17508
rect -3044 -17508 -2948 -17492
rect -4037 -17560 -3315 -17559
rect -4037 -18280 -4036 -17560
rect -3316 -18280 -3315 -17560
rect -4037 -18281 -3315 -18280
rect -4456 -18348 -4360 -18332
rect -3044 -18332 -3028 -17508
rect -2964 -18332 -2948 -17508
rect -1632 -17508 -1536 -17492
rect -2625 -17560 -1903 -17559
rect -2625 -18280 -2624 -17560
rect -1904 -18280 -1903 -17560
rect -2625 -18281 -1903 -18280
rect -3044 -18348 -2948 -18332
rect -1632 -18332 -1616 -17508
rect -1552 -18332 -1536 -17508
rect -220 -17508 -124 -17492
rect -1213 -17560 -491 -17559
rect -1213 -18280 -1212 -17560
rect -492 -18280 -491 -17560
rect -1213 -18281 -491 -18280
rect -1632 -18348 -1536 -18332
rect -220 -18332 -204 -17508
rect -140 -18332 -124 -17508
rect 1192 -17508 1288 -17492
rect 199 -17560 921 -17559
rect 199 -18280 200 -17560
rect 920 -18280 921 -17560
rect 199 -18281 921 -18280
rect -220 -18348 -124 -18332
rect 1192 -18332 1208 -17508
rect 1272 -18332 1288 -17508
rect 2604 -17508 2700 -17492
rect 1611 -17560 2333 -17559
rect 1611 -18280 1612 -17560
rect 2332 -18280 2333 -17560
rect 1611 -18281 2333 -18280
rect 1192 -18348 1288 -18332
rect 2604 -18332 2620 -17508
rect 2684 -18332 2700 -17508
rect 4016 -17508 4112 -17492
rect 3023 -17560 3745 -17559
rect 3023 -18280 3024 -17560
rect 3744 -18280 3745 -17560
rect 3023 -18281 3745 -18280
rect 2604 -18348 2700 -18332
rect 4016 -18332 4032 -17508
rect 4096 -18332 4112 -17508
rect 5428 -17508 5524 -17492
rect 4435 -17560 5157 -17559
rect 4435 -18280 4436 -17560
rect 5156 -18280 5157 -17560
rect 4435 -18281 5157 -18280
rect 4016 -18348 4112 -18332
rect 5428 -18332 5444 -17508
rect 5508 -18332 5524 -17508
rect 6840 -17508 6936 -17492
rect 5847 -17560 6569 -17559
rect 5847 -18280 5848 -17560
rect 6568 -18280 6569 -17560
rect 5847 -18281 6569 -18280
rect 5428 -18348 5524 -18332
rect 6840 -18332 6856 -17508
rect 6920 -18332 6936 -17508
rect 8252 -17508 8348 -17492
rect 7259 -17560 7981 -17559
rect 7259 -18280 7260 -17560
rect 7980 -18280 7981 -17560
rect 7259 -18281 7981 -18280
rect 6840 -18348 6936 -18332
rect 8252 -18332 8268 -17508
rect 8332 -18332 8348 -17508
rect 9664 -17508 9760 -17492
rect 8671 -17560 9393 -17559
rect 8671 -18280 8672 -17560
rect 9392 -18280 9393 -17560
rect 8671 -18281 9393 -18280
rect 8252 -18348 8348 -18332
rect 9664 -18332 9680 -17508
rect 9744 -18332 9760 -17508
rect 11076 -17508 11172 -17492
rect 10083 -17560 10805 -17559
rect 10083 -18280 10084 -17560
rect 10804 -18280 10805 -17560
rect 10083 -18281 10805 -18280
rect 9664 -18348 9760 -18332
rect 11076 -18332 11092 -17508
rect 11156 -18332 11172 -17508
rect 12488 -17508 12584 -17492
rect 11495 -17560 12217 -17559
rect 11495 -18280 11496 -17560
rect 12216 -18280 12217 -17560
rect 11495 -18281 12217 -18280
rect 11076 -18348 11172 -18332
rect 12488 -18332 12504 -17508
rect 12568 -18332 12584 -17508
rect 13900 -17508 13996 -17492
rect 12907 -17560 13629 -17559
rect 12907 -18280 12908 -17560
rect 13628 -18280 13629 -17560
rect 12907 -18281 13629 -18280
rect 12488 -18348 12584 -18332
rect 13900 -18332 13916 -17508
rect 13980 -18332 13996 -17508
rect 15312 -17508 15408 -17492
rect 14319 -17560 15041 -17559
rect 14319 -18280 14320 -17560
rect 15040 -18280 15041 -17560
rect 14319 -18281 15041 -18280
rect 13900 -18348 13996 -18332
rect 15312 -18332 15328 -17508
rect 15392 -18332 15408 -17508
rect 16724 -17508 16820 -17492
rect 15731 -17560 16453 -17559
rect 15731 -18280 15732 -17560
rect 16452 -18280 16453 -17560
rect 15731 -18281 16453 -18280
rect 15312 -18348 15408 -18332
rect 16724 -18332 16740 -17508
rect 16804 -18332 16820 -17508
rect 18136 -17508 18232 -17492
rect 17143 -17560 17865 -17559
rect 17143 -18280 17144 -17560
rect 17864 -18280 17865 -17560
rect 17143 -18281 17865 -18280
rect 16724 -18348 16820 -18332
rect 18136 -18332 18152 -17508
rect 18216 -18332 18232 -17508
rect 19548 -17508 19644 -17492
rect 18555 -17560 19277 -17559
rect 18555 -18280 18556 -17560
rect 19276 -18280 19277 -17560
rect 18555 -18281 19277 -18280
rect 18136 -18348 18232 -18332
rect 19548 -18332 19564 -17508
rect 19628 -18332 19644 -17508
rect 20960 -17508 21056 -17492
rect 19967 -17560 20689 -17559
rect 19967 -18280 19968 -17560
rect 20688 -18280 20689 -17560
rect 19967 -18281 20689 -18280
rect 19548 -18348 19644 -18332
rect 20960 -18332 20976 -17508
rect 21040 -18332 21056 -17508
rect 22372 -17508 22468 -17492
rect 21379 -17560 22101 -17559
rect 21379 -18280 21380 -17560
rect 22100 -18280 22101 -17560
rect 21379 -18281 22101 -18280
rect 20960 -18348 21056 -18332
rect 22372 -18332 22388 -17508
rect 22452 -18332 22468 -17508
rect 23784 -17508 23880 -17492
rect 22791 -17560 23513 -17559
rect 22791 -18280 22792 -17560
rect 23512 -18280 23513 -17560
rect 22791 -18281 23513 -18280
rect 22372 -18348 22468 -18332
rect 23784 -18332 23800 -17508
rect 23864 -18332 23880 -17508
rect 23784 -18348 23880 -18332
<< properties >>
string FIXED_BBOX 22712 17480 23592 18360
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 4 l 4 val 35.04 carea 2.00 cperi 0.19 nx 34 ny 33 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
<< end >>
