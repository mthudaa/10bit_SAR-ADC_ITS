magic
tech sky130A
magscale 1 2
timestamp 1749656160
<< nwell >>
rect 2369 -56 3107 1053
rect 2369 -115 3033 -56
<< pwell >>
rect -53 -149 1001 -115
rect 225 -201 1001 -149
rect -53 -3725 1001 -201
<< locali >>
rect -9799 1913 -9768 1947
rect -9734 1913 -9672 1947
rect -9638 1913 -9576 1947
rect -9542 1913 -9480 1947
rect -9446 1913 -9384 1947
rect -9350 1913 -9288 1947
rect -9254 1913 -9192 1947
rect -9158 1913 -9096 1947
rect -9062 1913 -9000 1947
rect -8966 1913 -8904 1947
rect -8870 1913 -8808 1947
rect -8774 1913 -8712 1947
rect -8678 1913 -8616 1947
rect -8582 1913 -8520 1947
rect -8486 1913 -8424 1947
rect -8390 1913 -8328 1947
rect -8294 1913 -8232 1947
rect -8198 1913 -8136 1947
rect -8102 1913 -8040 1947
rect -8006 1913 -7944 1947
rect -7910 1913 -7848 1947
rect -7814 1913 -7752 1947
rect -7718 1913 -7656 1947
rect -7622 1913 -7560 1947
rect -7526 1913 -7464 1947
rect -7430 1913 -7368 1947
rect -7334 1913 -7272 1947
rect -7238 1913 -7176 1947
rect -7142 1913 -7080 1947
rect -7046 1913 -6984 1947
rect -6950 1913 -6888 1947
rect -6854 1913 -6792 1947
rect -6758 1913 -6696 1947
rect -6662 1913 -6600 1947
rect -6566 1913 -6504 1947
rect -6470 1913 -6408 1947
rect -6374 1913 -6312 1947
rect -6278 1913 -6216 1947
rect -6182 1913 -6120 1947
rect -6086 1913 -6024 1947
rect -5990 1913 -5928 1947
rect -5894 1913 -5832 1947
rect -5798 1913 -5736 1947
rect -5702 1913 -5640 1947
rect -5606 1913 -5544 1947
rect -5510 1913 -5448 1947
rect -5414 1913 -5352 1947
rect -5318 1913 -5256 1947
rect -5222 1913 -5160 1947
rect -5126 1913 -5064 1947
rect -5030 1913 -4968 1947
rect -4934 1913 -4872 1947
rect -4838 1913 -4776 1947
rect -4742 1913 -4680 1947
rect -4646 1913 -4584 1947
rect -4550 1913 -4488 1947
rect -4454 1913 -4392 1947
rect -4358 1913 -4296 1947
rect -4262 1913 -4200 1947
rect -4166 1913 -4104 1947
rect -4070 1913 -4008 1947
rect -3974 1913 -3912 1947
rect -3878 1913 -3816 1947
rect -3782 1913 -3720 1947
rect -3686 1913 -3624 1947
rect -3590 1913 -3528 1947
rect -3494 1913 -3432 1947
rect -3398 1913 -3336 1947
rect -3302 1913 -3240 1947
rect -3206 1913 -3144 1947
rect -3110 1913 -3048 1947
rect -3014 1913 -2952 1947
rect -2918 1913 -2856 1947
rect -2822 1913 -2760 1947
rect -2726 1913 -2664 1947
rect -2630 1913 -2568 1947
rect -2534 1913 -2472 1947
rect -2438 1913 -2376 1947
rect -2342 1913 -2280 1947
rect -2246 1913 -2184 1947
rect -2150 1913 -2088 1947
rect -2054 1913 -1992 1947
rect -1958 1913 -1896 1947
rect -1862 1913 -1800 1947
rect -1766 1913 -1704 1947
rect -1670 1913 -1608 1947
rect -1574 1913 -1512 1947
rect -1478 1913 -1416 1947
rect -1382 1913 -1320 1947
rect -1286 1913 -1224 1947
rect -1190 1913 -1128 1947
rect -1094 1913 -1032 1947
rect -998 1913 -936 1947
rect -902 1913 -840 1947
rect -806 1913 -744 1947
rect -710 1913 -648 1947
rect -614 1913 -552 1947
rect -518 1913 -456 1947
rect -422 1913 -360 1947
rect -326 1913 -264 1947
rect -230 1913 -168 1947
rect -134 1913 -72 1947
rect -38 1913 24 1947
rect 58 1913 120 1947
rect 154 1913 216 1947
rect 250 1913 312 1947
rect 346 1913 408 1947
rect 442 1913 504 1947
rect 538 1913 600 1947
rect 634 1913 696 1947
rect 730 1913 792 1947
rect 826 1913 888 1947
rect 922 1913 984 1947
rect 1018 1913 1080 1947
rect 1114 1913 1176 1947
rect 1210 1913 1272 1947
rect 1306 1913 1368 1947
rect 1402 1913 1464 1947
rect 1498 1913 1529 1947
rect 79 367 237 1913
rect -9799 -4101 -9768 -4067
rect -9734 -4101 -9672 -4067
rect -9638 -4101 -9576 -4067
rect -9542 -4101 -9480 -4067
rect -9446 -4101 -9384 -4067
rect -9350 -4101 -9288 -4067
rect -9254 -4101 -9192 -4067
rect -9158 -4101 -9096 -4067
rect -9062 -4101 -9000 -4067
rect -8966 -4101 -8904 -4067
rect -8870 -4101 -8808 -4067
rect -8774 -4101 -8712 -4067
rect -8678 -4101 -8616 -4067
rect -8582 -4101 -8520 -4067
rect -8486 -4101 -8424 -4067
rect -8390 -4101 -8328 -4067
rect -8294 -4101 -8232 -4067
rect -8198 -4101 -8136 -4067
rect -8102 -4101 -8040 -4067
rect -8006 -4101 -7944 -4067
rect -7910 -4101 -7848 -4067
rect -7814 -4101 -7752 -4067
rect -7718 -4101 -7656 -4067
rect -7622 -4101 -7560 -4067
rect -7526 -4101 -7464 -4067
rect -7430 -4101 -7368 -4067
rect -7334 -4101 -7272 -4067
rect -7238 -4101 -7176 -4067
rect -7142 -4101 -7080 -4067
rect -7046 -4101 -6984 -4067
rect -6950 -4101 -6888 -4067
rect -6854 -4101 -6792 -4067
rect -6758 -4101 -6696 -4067
rect -6662 -4101 -6600 -4067
rect -6566 -4101 -6504 -4067
rect -6470 -4101 -6408 -4067
rect -6374 -4101 -6312 -4067
rect -6278 -4101 -6216 -4067
rect -6182 -4101 -6120 -4067
rect -6086 -4101 -6024 -4067
rect -5990 -4101 -5928 -4067
rect -5894 -4101 -5832 -4067
rect -5798 -4101 -5736 -4067
rect -5702 -4101 -5640 -4067
rect -5606 -4101 -5544 -4067
rect -5510 -4101 -5448 -4067
rect -5414 -4101 -5352 -4067
rect -5318 -4101 -5256 -4067
rect -5222 -4101 -5160 -4067
rect -5126 -4101 -5064 -4067
rect -5030 -4101 -4968 -4067
rect -4934 -4101 -4872 -4067
rect -4838 -4101 -4776 -4067
rect -4742 -4101 -4680 -4067
rect -4646 -4101 -4584 -4067
rect -4550 -4101 -4488 -4067
rect -4454 -4101 -4392 -4067
rect -4358 -4101 -4296 -4067
rect -4262 -4101 -4200 -4067
rect -4166 -4101 -4104 -4067
rect -4070 -4101 -4008 -4067
rect -3974 -4101 -3912 -4067
rect -3878 -4101 -3816 -4067
rect -3782 -4101 -3720 -4067
rect -3686 -4101 -3624 -4067
rect -3590 -4101 -3528 -4067
rect -3494 -4101 -3432 -4067
rect -3398 -4101 -3336 -4067
rect -3302 -4101 -3240 -4067
rect -3206 -4101 -3144 -4067
rect -3110 -4101 -3048 -4067
rect -3014 -4101 -2952 -4067
rect -2918 -4101 -2856 -4067
rect -2822 -4101 -2760 -4067
rect -2726 -4101 -2664 -4067
rect -2630 -4101 -2568 -4067
rect -2534 -4101 -2472 -4067
rect -2438 -4101 -2376 -4067
rect -2342 -4101 -2280 -4067
rect -2246 -4101 -2184 -4067
rect -2150 -4101 -2088 -4067
rect -2054 -4101 -1992 -4067
rect -1958 -4101 -1896 -4067
rect -1862 -4101 -1800 -4067
rect -1766 -4101 -1704 -4067
rect -1670 -4101 -1608 -4067
rect -1574 -4101 -1512 -4067
rect -1478 -4101 -1416 -4067
rect -1382 -4101 -1320 -4067
rect -1286 -4101 -1224 -4067
rect -1190 -4101 -1128 -4067
rect -1094 -4101 -1032 -4067
rect -998 -4101 -936 -4067
rect -902 -4101 -840 -4067
rect -806 -4101 -744 -4067
rect -710 -4101 -648 -4067
rect -614 -4101 -552 -4067
rect -518 -4101 -456 -4067
rect -422 -4101 -360 -4067
rect -326 -4101 -264 -4067
rect -230 -4101 -168 -4067
rect -134 -4101 -72 -4067
rect -38 -4101 24 -4067
rect 58 -4101 120 -4067
rect 154 -4101 216 -4067
rect 250 -4101 312 -4067
rect 346 -4101 408 -4067
rect 442 -4101 504 -4067
rect 538 -4101 600 -4067
rect 634 -4101 696 -4067
rect 730 -4101 792 -4067
rect 826 -4101 888 -4067
rect 922 -4101 984 -4067
rect 1018 -4101 1080 -4067
rect 1114 -4101 1176 -4067
rect 1210 -4101 1272 -4067
rect 1306 -4101 1368 -4067
rect 1402 -4101 1464 -4067
rect 1498 -4101 1529 -4067
<< viali >>
rect -9768 1913 -9734 1947
rect -9672 1913 -9638 1947
rect -9576 1913 -9542 1947
rect -9480 1913 -9446 1947
rect -9384 1913 -9350 1947
rect -9288 1913 -9254 1947
rect -9192 1913 -9158 1947
rect -9096 1913 -9062 1947
rect -9000 1913 -8966 1947
rect -8904 1913 -8870 1947
rect -8808 1913 -8774 1947
rect -8712 1913 -8678 1947
rect -8616 1913 -8582 1947
rect -8520 1913 -8486 1947
rect -8424 1913 -8390 1947
rect -8328 1913 -8294 1947
rect -8232 1913 -8198 1947
rect -8136 1913 -8102 1947
rect -8040 1913 -8006 1947
rect -7944 1913 -7910 1947
rect -7848 1913 -7814 1947
rect -7752 1913 -7718 1947
rect -7656 1913 -7622 1947
rect -7560 1913 -7526 1947
rect -7464 1913 -7430 1947
rect -7368 1913 -7334 1947
rect -7272 1913 -7238 1947
rect -7176 1913 -7142 1947
rect -7080 1913 -7046 1947
rect -6984 1913 -6950 1947
rect -6888 1913 -6854 1947
rect -6792 1913 -6758 1947
rect -6696 1913 -6662 1947
rect -6600 1913 -6566 1947
rect -6504 1913 -6470 1947
rect -6408 1913 -6374 1947
rect -6312 1913 -6278 1947
rect -6216 1913 -6182 1947
rect -6120 1913 -6086 1947
rect -6024 1913 -5990 1947
rect -5928 1913 -5894 1947
rect -5832 1913 -5798 1947
rect -5736 1913 -5702 1947
rect -5640 1913 -5606 1947
rect -5544 1913 -5510 1947
rect -5448 1913 -5414 1947
rect -5352 1913 -5318 1947
rect -5256 1913 -5222 1947
rect -5160 1913 -5126 1947
rect -5064 1913 -5030 1947
rect -4968 1913 -4934 1947
rect -4872 1913 -4838 1947
rect -4776 1913 -4742 1947
rect -4680 1913 -4646 1947
rect -4584 1913 -4550 1947
rect -4488 1913 -4454 1947
rect -4392 1913 -4358 1947
rect -4296 1913 -4262 1947
rect -4200 1913 -4166 1947
rect -4104 1913 -4070 1947
rect -4008 1913 -3974 1947
rect -3912 1913 -3878 1947
rect -3816 1913 -3782 1947
rect -3720 1913 -3686 1947
rect -3624 1913 -3590 1947
rect -3528 1913 -3494 1947
rect -3432 1913 -3398 1947
rect -3336 1913 -3302 1947
rect -3240 1913 -3206 1947
rect -3144 1913 -3110 1947
rect -3048 1913 -3014 1947
rect -2952 1913 -2918 1947
rect -2856 1913 -2822 1947
rect -2760 1913 -2726 1947
rect -2664 1913 -2630 1947
rect -2568 1913 -2534 1947
rect -2472 1913 -2438 1947
rect -2376 1913 -2342 1947
rect -2280 1913 -2246 1947
rect -2184 1913 -2150 1947
rect -2088 1913 -2054 1947
rect -1992 1913 -1958 1947
rect -1896 1913 -1862 1947
rect -1800 1913 -1766 1947
rect -1704 1913 -1670 1947
rect -1608 1913 -1574 1947
rect -1512 1913 -1478 1947
rect -1416 1913 -1382 1947
rect -1320 1913 -1286 1947
rect -1224 1913 -1190 1947
rect -1128 1913 -1094 1947
rect -1032 1913 -998 1947
rect -936 1913 -902 1947
rect -840 1913 -806 1947
rect -744 1913 -710 1947
rect -648 1913 -614 1947
rect -552 1913 -518 1947
rect -456 1913 -422 1947
rect -360 1913 -326 1947
rect -264 1913 -230 1947
rect -168 1913 -134 1947
rect -72 1913 -38 1947
rect 24 1913 58 1947
rect 120 1913 154 1947
rect 216 1913 250 1947
rect 312 1913 346 1947
rect 408 1913 442 1947
rect 504 1913 538 1947
rect 600 1913 634 1947
rect 696 1913 730 1947
rect 792 1913 826 1947
rect 888 1913 922 1947
rect 984 1913 1018 1947
rect 1080 1913 1114 1947
rect 1176 1913 1210 1947
rect 1272 1913 1306 1947
rect 1368 1913 1402 1947
rect 1464 1913 1498 1947
rect 79 333 237 367
rect 2721 139 2755 471
rect 237 -3689 395 -3655
rect -9768 -4101 -9734 -4067
rect -9672 -4101 -9638 -4067
rect -9576 -4101 -9542 -4067
rect -9480 -4101 -9446 -4067
rect -9384 -4101 -9350 -4067
rect -9288 -4101 -9254 -4067
rect -9192 -4101 -9158 -4067
rect -9096 -4101 -9062 -4067
rect -9000 -4101 -8966 -4067
rect -8904 -4101 -8870 -4067
rect -8808 -4101 -8774 -4067
rect -8712 -4101 -8678 -4067
rect -8616 -4101 -8582 -4067
rect -8520 -4101 -8486 -4067
rect -8424 -4101 -8390 -4067
rect -8328 -4101 -8294 -4067
rect -8232 -4101 -8198 -4067
rect -8136 -4101 -8102 -4067
rect -8040 -4101 -8006 -4067
rect -7944 -4101 -7910 -4067
rect -7848 -4101 -7814 -4067
rect -7752 -4101 -7718 -4067
rect -7656 -4101 -7622 -4067
rect -7560 -4101 -7526 -4067
rect -7464 -4101 -7430 -4067
rect -7368 -4101 -7334 -4067
rect -7272 -4101 -7238 -4067
rect -7176 -4101 -7142 -4067
rect -7080 -4101 -7046 -4067
rect -6984 -4101 -6950 -4067
rect -6888 -4101 -6854 -4067
rect -6792 -4101 -6758 -4067
rect -6696 -4101 -6662 -4067
rect -6600 -4101 -6566 -4067
rect -6504 -4101 -6470 -4067
rect -6408 -4101 -6374 -4067
rect -6312 -4101 -6278 -4067
rect -6216 -4101 -6182 -4067
rect -6120 -4101 -6086 -4067
rect -6024 -4101 -5990 -4067
rect -5928 -4101 -5894 -4067
rect -5832 -4101 -5798 -4067
rect -5736 -4101 -5702 -4067
rect -5640 -4101 -5606 -4067
rect -5544 -4101 -5510 -4067
rect -5448 -4101 -5414 -4067
rect -5352 -4101 -5318 -4067
rect -5256 -4101 -5222 -4067
rect -5160 -4101 -5126 -4067
rect -5064 -4101 -5030 -4067
rect -4968 -4101 -4934 -4067
rect -4872 -4101 -4838 -4067
rect -4776 -4101 -4742 -4067
rect -4680 -4101 -4646 -4067
rect -4584 -4101 -4550 -4067
rect -4488 -4101 -4454 -4067
rect -4392 -4101 -4358 -4067
rect -4296 -4101 -4262 -4067
rect -4200 -4101 -4166 -4067
rect -4104 -4101 -4070 -4067
rect -4008 -4101 -3974 -4067
rect -3912 -4101 -3878 -4067
rect -3816 -4101 -3782 -4067
rect -3720 -4101 -3686 -4067
rect -3624 -4101 -3590 -4067
rect -3528 -4101 -3494 -4067
rect -3432 -4101 -3398 -4067
rect -3336 -4101 -3302 -4067
rect -3240 -4101 -3206 -4067
rect -3144 -4101 -3110 -4067
rect -3048 -4101 -3014 -4067
rect -2952 -4101 -2918 -4067
rect -2856 -4101 -2822 -4067
rect -2760 -4101 -2726 -4067
rect -2664 -4101 -2630 -4067
rect -2568 -4101 -2534 -4067
rect -2472 -4101 -2438 -4067
rect -2376 -4101 -2342 -4067
rect -2280 -4101 -2246 -4067
rect -2184 -4101 -2150 -4067
rect -2088 -4101 -2054 -4067
rect -1992 -4101 -1958 -4067
rect -1896 -4101 -1862 -4067
rect -1800 -4101 -1766 -4067
rect -1704 -4101 -1670 -4067
rect -1608 -4101 -1574 -4067
rect -1512 -4101 -1478 -4067
rect -1416 -4101 -1382 -4067
rect -1320 -4101 -1286 -4067
rect -1224 -4101 -1190 -4067
rect -1128 -4101 -1094 -4067
rect -1032 -4101 -998 -4067
rect -936 -4101 -902 -4067
rect -840 -4101 -806 -4067
rect -744 -4101 -710 -4067
rect -648 -4101 -614 -4067
rect -552 -4101 -518 -4067
rect -456 -4101 -422 -4067
rect -360 -4101 -326 -4067
rect -264 -4101 -230 -4067
rect -168 -4101 -134 -4067
rect -72 -4101 -38 -4067
rect 24 -4101 58 -4067
rect 120 -4101 154 -4067
rect 216 -4101 250 -4067
rect 312 -4101 346 -4067
rect 408 -4101 442 -4067
rect 504 -4101 538 -4067
rect 600 -4101 634 -4067
rect 696 -4101 730 -4067
rect 792 -4101 826 -4067
rect 888 -4101 922 -4067
rect 984 -4101 1018 -4067
rect 1080 -4101 1114 -4067
rect 1176 -4101 1210 -4067
rect 1272 -4101 1306 -4067
rect 1368 -4101 1402 -4067
rect 1464 -4101 1498 -4067
<< metal1 >>
rect -9799 1947 1529 1978
rect -9799 1913 -9768 1947
rect -9734 1913 -9672 1947
rect -9638 1913 -9576 1947
rect -9542 1913 -9480 1947
rect -9446 1913 -9384 1947
rect -9350 1913 -9288 1947
rect -9254 1913 -9192 1947
rect -9158 1913 -9096 1947
rect -9062 1913 -9000 1947
rect -8966 1913 -8904 1947
rect -8870 1913 -8808 1947
rect -8774 1913 -8712 1947
rect -8678 1913 -8616 1947
rect -8582 1913 -8520 1947
rect -8486 1913 -8424 1947
rect -8390 1913 -8328 1947
rect -8294 1913 -8232 1947
rect -8198 1913 -8136 1947
rect -8102 1913 -8040 1947
rect -8006 1913 -7944 1947
rect -7910 1913 -7848 1947
rect -7814 1913 -7752 1947
rect -7718 1913 -7656 1947
rect -7622 1913 -7560 1947
rect -7526 1913 -7464 1947
rect -7430 1913 -7368 1947
rect -7334 1913 -7272 1947
rect -7238 1913 -7176 1947
rect -7142 1913 -7080 1947
rect -7046 1913 -6984 1947
rect -6950 1913 -6888 1947
rect -6854 1913 -6792 1947
rect -6758 1913 -6696 1947
rect -6662 1913 -6600 1947
rect -6566 1913 -6504 1947
rect -6470 1913 -6408 1947
rect -6374 1913 -6312 1947
rect -6278 1913 -6216 1947
rect -6182 1913 -6120 1947
rect -6086 1913 -6024 1947
rect -5990 1913 -5928 1947
rect -5894 1913 -5832 1947
rect -5798 1913 -5736 1947
rect -5702 1913 -5640 1947
rect -5606 1913 -5544 1947
rect -5510 1913 -5448 1947
rect -5414 1913 -5352 1947
rect -5318 1913 -5256 1947
rect -5222 1913 -5160 1947
rect -5126 1913 -5064 1947
rect -5030 1913 -4968 1947
rect -4934 1913 -4872 1947
rect -4838 1913 -4776 1947
rect -4742 1913 -4680 1947
rect -4646 1913 -4584 1947
rect -4550 1913 -4488 1947
rect -4454 1913 -4392 1947
rect -4358 1913 -4296 1947
rect -4262 1913 -4200 1947
rect -4166 1913 -4104 1947
rect -4070 1913 -4008 1947
rect -3974 1913 -3912 1947
rect -3878 1913 -3816 1947
rect -3782 1913 -3720 1947
rect -3686 1913 -3624 1947
rect -3590 1913 -3528 1947
rect -3494 1913 -3432 1947
rect -3398 1913 -3336 1947
rect -3302 1913 -3240 1947
rect -3206 1913 -3144 1947
rect -3110 1913 -3048 1947
rect -3014 1913 -2952 1947
rect -2918 1913 -2856 1947
rect -2822 1913 -2760 1947
rect -2726 1913 -2664 1947
rect -2630 1913 -2568 1947
rect -2534 1913 -2472 1947
rect -2438 1913 -2376 1947
rect -2342 1913 -2280 1947
rect -2246 1913 -2184 1947
rect -2150 1913 -2088 1947
rect -2054 1913 -1992 1947
rect -1958 1913 -1896 1947
rect -1862 1913 -1800 1947
rect -1766 1913 -1704 1947
rect -1670 1913 -1608 1947
rect -1574 1913 -1512 1947
rect -1478 1913 -1416 1947
rect -1382 1913 -1320 1947
rect -1286 1913 -1224 1947
rect -1190 1913 -1128 1947
rect -1094 1913 -1032 1947
rect -998 1913 -936 1947
rect -902 1913 -840 1947
rect -806 1913 -744 1947
rect -710 1913 -648 1947
rect -614 1913 -552 1947
rect -518 1913 -456 1947
rect -422 1913 -360 1947
rect -326 1913 -264 1947
rect -230 1913 -168 1947
rect -134 1913 -72 1947
rect -38 1913 24 1947
rect 58 1913 120 1947
rect 154 1913 216 1947
rect 250 1913 312 1947
rect 346 1913 408 1947
rect 442 1913 504 1947
rect 538 1913 600 1947
rect 634 1913 696 1947
rect 730 1913 792 1947
rect 826 1913 888 1947
rect 922 1913 984 1947
rect 1018 1913 1080 1947
rect 1114 1913 1176 1947
rect 1210 1913 1272 1947
rect 1306 1913 1368 1947
rect 1402 1913 1464 1947
rect 1498 1913 1529 1947
rect -9799 1882 1529 1913
rect 79 1053 237 1882
rect 79 981 2523 1053
rect 79 507 237 981
rect 79 455 448 507
rect 500 455 510 507
rect 79 373 237 455
rect 67 367 249 373
rect 67 333 79 367
rect 237 333 249 367
rect 67 327 249 333
rect 91 220 137 327
rect 215 104 225 254
rect 277 104 287 254
rect -281 -45 -271 59
rect -167 -45 -157 59
rect 122 11 132 63
rect 184 11 194 63
rect 2451 33 2523 981
rect 2551 874 2963 926
rect 3015 874 3025 926
rect 2607 471 2870 505
rect 2607 139 2712 471
rect 2764 139 2870 471
rect 2607 105 2870 139
rect 2953 105 2963 505
rect 3015 105 3025 505
rect 2860 12 2870 64
rect 2922 12 2932 64
rect -281 -97 2712 -45
rect 2764 -97 2774 -45
rect -281 -201 -271 -97
rect -167 -201 -157 -97
rect 215 -201 225 -149
rect 277 -201 857 -149
rect 909 -201 2870 -149
rect 2922 -201 2932 -149
rect 122 -293 132 -241
rect 184 -293 194 -241
rect 438 -293 448 -241
rect 500 -293 510 -241
rect 29 -425 39 -325
rect 91 -425 101 -325
rect 215 -425 225 -325
rect 277 -425 287 -325
rect 345 -1825 355 -325
rect 407 -1825 417 -325
rect 531 -1847 541 -325
rect 593 -377 2963 -325
rect 3015 -377 3025 -325
rect 593 -1795 603 -377
rect 661 -1763 671 -963
rect 723 -1763 733 -963
rect 847 -1763 857 -963
rect 909 -1763 919 -963
rect 593 -1847 764 -1795
rect 816 -1847 1433 -1795
rect 29 -1955 39 -1903
rect 91 -1955 671 -1903
rect 723 -1955 733 -1903
rect 29 -3515 39 -3115
rect 91 -3515 101 -3115
rect 215 -3515 225 -3115
rect 277 -3515 287 -3115
rect 345 -3515 355 -2015
rect 407 -3515 417 -2015
rect 531 -3515 541 -2015
rect 593 -3515 603 -2015
rect 754 -2045 764 -1993
rect 816 -2045 826 -1993
rect 661 -2877 671 -2077
rect 723 -2877 733 -2077
rect 817 -2451 851 -2443
rect 817 -2503 1433 -2451
rect 817 -2511 851 -2503
rect 129 -3587 1433 -3553
rect 215 -3701 225 -3649
rect 277 -3655 541 -3649
rect 395 -3689 541 -3655
rect 277 -3701 541 -3689
rect 593 -3701 603 -3649
rect 237 -4036 395 -3701
rect -9799 -4067 1529 -4036
rect -9799 -4101 -9768 -4067
rect -9734 -4101 -9672 -4067
rect -9638 -4101 -9576 -4067
rect -9542 -4101 -9480 -4067
rect -9446 -4101 -9384 -4067
rect -9350 -4101 -9288 -4067
rect -9254 -4101 -9192 -4067
rect -9158 -4101 -9096 -4067
rect -9062 -4101 -9000 -4067
rect -8966 -4101 -8904 -4067
rect -8870 -4101 -8808 -4067
rect -8774 -4101 -8712 -4067
rect -8678 -4101 -8616 -4067
rect -8582 -4101 -8520 -4067
rect -8486 -4101 -8424 -4067
rect -8390 -4101 -8328 -4067
rect -8294 -4101 -8232 -4067
rect -8198 -4101 -8136 -4067
rect -8102 -4101 -8040 -4067
rect -8006 -4101 -7944 -4067
rect -7910 -4101 -7848 -4067
rect -7814 -4101 -7752 -4067
rect -7718 -4101 -7656 -4067
rect -7622 -4101 -7560 -4067
rect -7526 -4101 -7464 -4067
rect -7430 -4101 -7368 -4067
rect -7334 -4101 -7272 -4067
rect -7238 -4101 -7176 -4067
rect -7142 -4101 -7080 -4067
rect -7046 -4101 -6984 -4067
rect -6950 -4101 -6888 -4067
rect -6854 -4101 -6792 -4067
rect -6758 -4101 -6696 -4067
rect -6662 -4101 -6600 -4067
rect -6566 -4101 -6504 -4067
rect -6470 -4101 -6408 -4067
rect -6374 -4101 -6312 -4067
rect -6278 -4101 -6216 -4067
rect -6182 -4101 -6120 -4067
rect -6086 -4101 -6024 -4067
rect -5990 -4101 -5928 -4067
rect -5894 -4101 -5832 -4067
rect -5798 -4101 -5736 -4067
rect -5702 -4101 -5640 -4067
rect -5606 -4101 -5544 -4067
rect -5510 -4101 -5448 -4067
rect -5414 -4101 -5352 -4067
rect -5318 -4101 -5256 -4067
rect -5222 -4101 -5160 -4067
rect -5126 -4101 -5064 -4067
rect -5030 -4101 -4968 -4067
rect -4934 -4101 -4872 -4067
rect -4838 -4101 -4776 -4067
rect -4742 -4101 -4680 -4067
rect -4646 -4101 -4584 -4067
rect -4550 -4101 -4488 -4067
rect -4454 -4101 -4392 -4067
rect -4358 -4101 -4296 -4067
rect -4262 -4101 -4200 -4067
rect -4166 -4101 -4104 -4067
rect -4070 -4101 -4008 -4067
rect -3974 -4101 -3912 -4067
rect -3878 -4101 -3816 -4067
rect -3782 -4101 -3720 -4067
rect -3686 -4101 -3624 -4067
rect -3590 -4101 -3528 -4067
rect -3494 -4101 -3432 -4067
rect -3398 -4101 -3336 -4067
rect -3302 -4101 -3240 -4067
rect -3206 -4101 -3144 -4067
rect -3110 -4101 -3048 -4067
rect -3014 -4101 -2952 -4067
rect -2918 -4101 -2856 -4067
rect -2822 -4101 -2760 -4067
rect -2726 -4101 -2664 -4067
rect -2630 -4101 -2568 -4067
rect -2534 -4101 -2472 -4067
rect -2438 -4101 -2376 -4067
rect -2342 -4101 -2280 -4067
rect -2246 -4101 -2184 -4067
rect -2150 -4101 -2088 -4067
rect -2054 -4101 -1992 -4067
rect -1958 -4101 -1896 -4067
rect -1862 -4101 -1800 -4067
rect -1766 -4101 -1704 -4067
rect -1670 -4101 -1608 -4067
rect -1574 -4101 -1512 -4067
rect -1478 -4101 -1416 -4067
rect -1382 -4101 -1320 -4067
rect -1286 -4101 -1224 -4067
rect -1190 -4101 -1128 -4067
rect -1094 -4101 -1032 -4067
rect -998 -4101 -936 -4067
rect -902 -4101 -840 -4067
rect -806 -4101 -744 -4067
rect -710 -4101 -648 -4067
rect -614 -4101 -552 -4067
rect -518 -4101 -456 -4067
rect -422 -4101 -360 -4067
rect -326 -4101 -264 -4067
rect -230 -4101 -168 -4067
rect -134 -4101 -72 -4067
rect -38 -4101 24 -4067
rect 58 -4101 120 -4067
rect 154 -4101 216 -4067
rect 250 -4101 312 -4067
rect 346 -4101 408 -4067
rect 442 -4101 504 -4067
rect 538 -4101 600 -4067
rect 634 -4101 696 -4067
rect 730 -4101 792 -4067
rect 826 -4101 888 -4067
rect 922 -4101 984 -4067
rect 1018 -4101 1080 -4067
rect 1114 -4101 1176 -4067
rect 1210 -4101 1272 -4067
rect 1306 -4101 1368 -4067
rect 1402 -4101 1464 -4067
rect 1498 -4101 1529 -4067
rect -9799 -4132 1529 -4101
<< via1 >>
rect 448 455 500 507
rect 225 104 277 254
rect -271 -45 -167 59
rect 132 11 184 63
rect 2963 874 3015 926
rect 2712 139 2721 471
rect 2721 139 2755 471
rect 2755 139 2764 471
rect 2963 105 3015 505
rect 2870 12 2922 64
rect 2712 -97 2764 -45
rect -271 -201 -167 -97
rect 225 -201 277 -149
rect 857 -201 909 -149
rect 2870 -201 2922 -149
rect 132 -293 184 -241
rect 448 -293 500 -241
rect 39 -425 91 -325
rect 225 -425 277 -325
rect 355 -1825 407 -325
rect 541 -1847 593 -325
rect 2963 -377 3015 -325
rect 671 -1763 723 -963
rect 857 -1763 909 -963
rect 764 -1847 816 -1795
rect 39 -1955 91 -1903
rect 671 -1955 723 -1903
rect 39 -3515 91 -3115
rect 225 -3515 277 -3115
rect 355 -3515 407 -2015
rect 541 -3515 593 -2015
rect 764 -2045 816 -1993
rect 671 -2877 723 -2077
rect 225 -3655 277 -3649
rect 225 -3689 237 -3655
rect 237 -3689 277 -3655
rect 225 -3701 277 -3689
rect 541 -3701 593 -3649
<< metal2 >>
rect 2963 926 3015 936
rect 448 507 500 517
rect 2963 505 3015 874
rect 225 254 277 264
rect -271 59 -167 69
rect -271 -55 -167 -45
rect 132 63 184 73
rect 132 -77 184 11
rect 128 -87 184 -77
rect -271 -97 -167 -87
rect 128 -153 184 -143
rect -271 -211 -167 -201
rect 132 -241 184 -153
rect 132 -303 184 -293
rect 225 -149 277 104
rect 39 -325 91 -315
rect 39 -1903 91 -425
rect 225 -325 277 -201
rect 448 -241 500 455
rect 2712 471 2764 481
rect 2712 -45 2764 139
rect 2712 -107 2764 -97
rect 2870 64 2922 74
rect 448 -303 500 -293
rect 857 -149 909 -139
rect 225 -435 277 -425
rect 355 -325 407 -315
rect 39 -2543 91 -1955
rect 35 -2553 91 -2543
rect 35 -2713 91 -2609
rect 35 -2779 91 -2769
rect 39 -3115 91 -2779
rect 355 -2015 407 -1825
rect 541 -325 593 -315
rect 541 -1857 593 -1847
rect 671 -963 723 -953
rect 671 -1903 723 -1763
rect 857 -963 909 -201
rect 2870 -149 2922 12
rect 2870 -211 2922 -201
rect 2963 -325 3015 105
rect 2963 -387 3015 -377
rect 857 -1773 909 -1763
rect 39 -3525 91 -3515
rect 225 -3115 277 -3105
rect 225 -3649 277 -3515
rect 355 -3525 407 -3515
rect 541 -2015 593 -2005
rect 671 -2077 723 -1955
rect 764 -1795 816 -1785
rect 764 -1993 816 -1847
rect 764 -2055 816 -2045
rect 671 -2887 723 -2877
rect 225 -3711 277 -3701
rect 541 -3649 593 -3515
rect 541 -3711 593 -3701
<< via2 >>
rect -271 -45 -167 59
rect -271 -201 -167 -97
rect 128 -143 184 -87
rect 35 -2609 91 -2553
rect 35 -2769 91 -2713
<< metal3 >>
rect -281 59 -157 64
rect -281 -45 -271 59
rect -167 -45 -157 59
rect -281 -97 -157 -45
rect -281 -201 -271 -97
rect -167 -201 -157 -97
rect 118 -87 1433 -82
rect 118 -143 128 -87
rect 184 -143 1433 -87
rect 118 -148 1433 -143
rect -281 -206 -157 -201
rect 25 -2553 101 -2548
rect 25 -2609 35 -2553
rect 91 -2609 101 -2553
rect -505 -2713 -495 -2609
rect -375 -2713 101 -2609
rect 25 -2769 35 -2713
rect 91 -2769 101 -2713
rect 25 -2774 101 -2769
<< via3 >>
rect -271 -45 -167 59
rect -271 -201 -167 -97
rect -495 -2713 -375 -2609
<< metal4 >>
rect -9543 1523 -9335 1627
rect -9543 215 -9439 1523
rect -375 843 -167 947
rect -9543 111 -9229 215
rect -9543 -1197 -9439 111
rect -271 60 -167 843
rect -272 59 -166 60
rect -272 -45 -271 59
rect -167 -45 -166 59
rect -272 -97 -166 -45
rect -272 -201 -271 -97
rect -167 -201 -166 -97
rect -272 -202 -166 -201
rect -271 -465 -167 -202
rect -375 -569 -167 -465
rect -9543 -1301 -9224 -1197
rect -9543 -2609 -9439 -1301
rect -271 -1877 -167 -569
rect -375 -1981 -167 -1877
rect -496 -2609 -374 -2608
rect -9543 -2713 -9231 -2609
rect -496 -2713 -495 -2609
rect -375 -2713 -374 -2609
rect -496 -2714 -374 -2713
rect -271 -3289 -167 -1981
rect -375 -3393 -167 -3289
use sky130_fd_pr__nfet_01v8_J4Y94J  sky130_fd_pr__nfet_01v8_J4Y94J_0
timestamp 1749313676
transform 1 0 790 0 1 -2446
box -211 -579 211 579
use sky130_fd_pr__cap_mim_m3_1_9XU9T9  XC1
timestamp 1749307785
transform 0 1 -4855 1 0 -1077
box -2704 -4480 2704 4480
use sky130_fd_pr__pfet_01v8_27QFPY  XM1
timestamp 1749310734
transform 1 0 158 0 1 144
box -211 -259 211 259
use sky130_fd_pr__pfet_01v8_MGASDN  XM2
timestamp 1749313676
transform 1 0 2580 0 1 469
box -211 -584 211 584
use sky130_fd_pr__pfet_01v8_LGMQDL  XM3
timestamp 1749313676
transform 1 0 2896 0 1 269
box -211 -384 211 384
use sky130_fd_pr__nfet_01v8_CQKS6Z  XM4
timestamp 1749307785
transform 1 0 158 0 1 -344
box -211 -229 211 229
use sky130_fd_pr__nfet_01v8_46WN23  XM5
timestamp 1749310734
transform 1 0 158 0 1 -3346
box -211 -379 211 379
use sky130_fd_pr__nfet_01v8_J47Z3J  XM6
timestamp 1749313676
transform 1 0 790 0 1 -1394
box -211 -579 211 579
use sky130_fd_pr__nfet_01v8_D4Y996  XM8
timestamp 1749307785
transform 1 0 474 0 1 -1044
box -211 -929 211 929
use sky130_fd_pr__nfet_01v8_D47ZC5  XM9
timestamp 1749310734
transform 1 0 474 0 1 -2796
box -211 -929 211 929
<< labels >>
flabel viali 1464 1913 1498 1947 0 FreeSans 400 0 0 0 VDD
port 0 nsew
flabel viali 1464 -4101 1498 -4067 0 FreeSans 400 0 0 0 VSS
port 1 nsew
flabel metal1 1390 -2494 1424 -2460 0 FreeSans 400 0 0 0 IN
port 2 nsew
flabel metal1 1389 -1839 1423 -1805 0 FreeSans 400 0 0 0 VGS
port 3 nsew
flabel metal1 1399 -3587 1433 -3553 0 FreeSans 400 0 0 0 CK
port 5 nsew
flabel metal3 1378 -139 1412 -105 0 FreeSans 400 0 0 0 CKB
port 7 nsew
<< end >>
