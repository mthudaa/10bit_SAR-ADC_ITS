magic
tech sky130A
magscale 1 2
timestamp 1749223325
<< nwell >>
rect -875 248 805 998
rect -875 4 249 248
<< pwell >>
rect 249 4 805 206
rect -875 -417 805 4
rect -875 -482 805 -451
<< psubdiff >>
rect -819 -76 -785 -52
rect -819 -276 -785 -252
rect 159 -76 193 -52
rect 159 -276 193 -252
<< nsubdiff >>
rect -819 692 -785 716
rect -819 92 -785 116
rect 159 692 193 716
rect 159 92 193 116
<< psubdiffcont >>
rect -819 -252 -785 -76
rect 159 -252 193 -76
<< nsubdiffcont >>
rect -819 116 -785 692
rect 159 116 193 692
<< poly >>
rect -671 -62 -471 98
rect -155 -58 45 102
<< locali >>
rect -875 933 -844 967
rect -810 933 -748 967
rect -714 933 -652 967
rect -618 933 -556 967
rect -522 933 -460 967
rect -426 933 -364 967
rect -330 933 -268 967
rect -234 933 -172 967
rect -138 933 -76 967
rect -42 933 20 967
rect 54 933 116 967
rect 150 933 212 967
rect 246 933 308 967
rect 342 933 404 967
rect 438 933 500 967
rect 534 933 596 967
rect 630 933 692 967
rect 726 933 788 967
rect 822 933 853 967
rect -819 692 -785 933
rect -459 704 -425 933
rect 159 692 193 933
rect -819 100 -785 116
rect -717 57 -683 207
rect -717 23 -77 57
rect -819 -76 -785 -60
rect -717 -64 -683 23
rect 57 14 91 172
rect 193 565 482 599
rect 159 100 193 116
rect 57 -20 367 14
rect 57 -68 91 -20
rect 159 -67 193 -60
rect -819 -417 -785 -252
rect 159 -76 386 -67
rect 193 -101 386 -76
rect -201 -417 -167 -266
rect 159 -417 193 -252
rect -875 -451 -844 -417
rect -810 -451 -748 -417
rect -714 -451 -652 -417
rect -618 -451 -556 -417
rect -522 -451 -460 -417
rect -426 -451 -364 -417
rect -330 -451 -268 -417
rect -234 -451 -172 -417
rect -138 -451 -76 -417
rect -42 -451 20 -417
rect 54 -451 116 -417
rect 150 -451 212 -417
rect 246 -451 308 -417
rect 342 -451 404 -417
rect 438 -451 500 -417
rect 534 -451 596 -417
rect 630 -451 692 -417
rect 726 -451 788 -417
rect 822 -451 853 -417
<< viali >>
rect -844 933 -810 967
rect -748 933 -714 967
rect -652 933 -618 967
rect -556 933 -522 967
rect -460 933 -426 967
rect -364 933 -330 967
rect -268 933 -234 967
rect -172 933 -138 967
rect -76 933 -42 967
rect 20 933 54 967
rect 116 933 150 967
rect 212 933 246 967
rect 308 933 342 967
rect 404 933 438 967
rect 500 933 534 967
rect 596 933 630 967
rect 692 933 726 967
rect 788 933 822 967
rect 518 202 552 236
rect 750 210 784 244
rect -844 -451 -810 -417
rect -748 -451 -714 -417
rect -652 -451 -618 -417
rect -556 -451 -522 -417
rect -460 -451 -426 -417
rect -364 -451 -330 -417
rect -268 -451 -234 -417
rect -172 -451 -138 -417
rect -76 -451 -42 -417
rect 20 -451 54 -417
rect 116 -451 150 -417
rect 212 -451 246 -417
rect 308 -451 342 -417
rect 404 -451 438 -417
rect 500 -451 534 -417
rect 596 -451 630 -417
rect 692 -451 726 -417
rect 788 -451 822 -417
<< metal1 >>
rect -875 967 853 998
rect -875 933 -844 967
rect -810 933 -748 967
rect -714 933 -652 967
rect -618 933 -556 967
rect -522 933 -460 967
rect -426 933 -364 967
rect -330 933 -268 967
rect -234 933 -172 967
rect -138 933 -76 967
rect -42 933 20 967
rect 54 933 116 967
rect 150 933 212 967
rect 246 933 308 967
rect 342 933 404 967
rect 438 933 500 967
rect 534 933 596 967
rect 630 933 692 967
rect 726 933 788 967
rect 822 933 853 967
rect -875 902 853 933
rect -875 825 -259 859
rect -635 785 -625 794
rect -875 751 -625 785
rect -635 742 -625 751
rect -517 742 -507 794
rect -367 791 -259 825
rect 736 569 767 902
rect 492 186 502 252
rect 568 186 578 252
rect 738 244 842 253
rect 738 210 750 244
rect 784 210 842 244
rect 738 201 842 210
rect -875 -336 -259 -302
rect 735 -386 767 -101
rect -875 -417 853 -386
rect -875 -451 -844 -417
rect -810 -451 -748 -417
rect -714 -451 -652 -417
rect -618 -451 -556 -417
rect -522 -451 -460 -417
rect -426 -451 -364 -417
rect -330 -451 -268 -417
rect -234 -451 -172 -417
rect -138 -451 -76 -417
rect -42 -451 20 -417
rect 54 -451 116 -417
rect 150 -451 212 -417
rect 246 -451 308 -417
rect 342 -451 404 -417
rect 438 -451 500 -417
rect 534 -451 596 -417
rect 630 -451 692 -417
rect 726 -451 788 -417
rect 822 -451 853 -417
rect -875 -482 853 -451
<< via1 >>
rect -625 742 -517 794
rect 502 236 568 252
rect 502 202 518 236
rect 518 202 552 236
rect 552 202 568 236
rect 502 186 568 202
<< metal2 >>
rect -625 796 -517 806
rect -625 730 -517 740
rect 502 801 568 811
rect 502 252 568 735
rect 502 176 568 186
<< via2 >>
rect -625 794 -517 796
rect -625 742 -517 794
rect -625 740 -517 742
rect 502 735 568 801
<< metal3 >>
rect 492 801 578 806
rect -635 796 502 801
rect -635 740 -625 796
rect -517 740 502 796
rect -635 735 502 740
rect 568 735 578 801
rect 492 730 578 735
use sky130_fd_pr__nfet_01v8_3KLK8B  sky130_fd_pr__nfet_01v8_3KLK8B_0
timestamp 1749060920
transform 1 0 -313 0 1 -195
box -158 -157 158 157
use sky130_fd_pr__nfet_01v8_WVKZ6V  sky130_fd_pr__nfet_01v8_WVKZ6V_0
timestamp 1749054394
transform 1 0 -55 0 1 -164
box -158 -126 158 126
use sky130_fd_pr__pfet_01v8_GLM8QU  sky130_fd_pr__pfet_01v8_GLM8QU_0
timestamp 1749060920
transform 1 0 -55 0 1 368
box -194 -364 194 398
use sky130_fd_pr__pfet_01v8_JKM84M  sky130_fd_pr__pfet_01v8_JKM84M_0
timestamp 1749060920
transform 1 0 -571 0 1 440
box -194 -398 194 364
use sky130_fd_sc_hs__and2_1  sky130_fd_sc_hs__and2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749223325
transform 1 0 287 0 1 -84
box -38 -49 518 715
use sky130_fd_pr__pfet_01v8_JKM84M  XM1
timestamp 1749060920
transform 1 0 -313 0 1 440
box -194 -398 194 364
use sky130_fd_pr__nfet_01v8_WVKZ6V  XM5
timestamp 1749054394
transform 1 0 -571 0 1 -164
box -158 -126 158 126
<< labels >>
flabel nwell -813 930 -783 960 0 FreeSans 400 0 0 0 VDD
port 0 nsew
flabel metal1 -831 -452 -801 -422 0 FreeSans 400 0 0 0 VSS
port 1 nsew
flabel metal1 -875 825 -841 859 0 FreeSans 400 0 0 0 VINP
port 2 nsew
flabel metal1 -875 -336 -841 -302 0 FreeSans 400 0 0 0 VINN
port 3 nsew
flabel metal1 784 201 842 253 0 FreeSans 400 0 0 0 OUT
port 5 nsew
flabel metal1 -875 751 -841 785 0 FreeSans 400 0 0 0 IN
port 7 nsew
<< end >>
