magic
tech sky130A
magscale 1 2
timestamp 1748790007
<< viali >>
rect 142 1527 7228 1561
rect 142 -123 3740 -89
<< metal1 >>
rect 106 1561 7264 1597
rect 106 1527 142 1561
rect 7228 1527 7264 1561
rect 106 1521 7264 1527
rect 325 1447 7045 1521
rect 106 1301 176 1401
rect 228 1301 284 1401
rect 325 1061 7045 1255
rect 106 915 284 1015
rect 106 569 7264 869
rect 106 423 284 523
rect 316 183 3566 377
rect 166 37 176 137
rect 228 37 284 137
rect 316 -83 3566 -9
rect 106 -89 7264 -83
rect 106 -123 142 -89
rect 3740 -123 7264 -89
rect 106 -159 7264 -123
<< via1 >>
rect 176 1301 228 1401
rect 176 37 228 137
<< metal2 >>
rect 176 1401 228 1411
rect 176 137 228 1301
rect 176 27 228 37
use sky130_fd_pr__nfet_01v8_K9ZN2D  sky130_fd_pr__nfet_01v8_K9ZN2D_0
timestamp 1746379951
transform 0 1 1941 -1 0 87
box -246 -1835 246 1835
use sky130_fd_pr__pfet_01v8_D9Q5W2  sky130_fd_pr__pfet_01v8_D9Q5W2_0
timestamp 1746379951
transform 0 1 3685 -1 0 965
box -246 -3579 246 3579
use sky130_fd_pr__pfet_01v8_D9Q5W2  XM1
timestamp 1746379951
transform 0 1 3685 -1 0 1351
box -246 -3579 246 3579
use sky130_fd_pr__nfet_01v8_K9ZN2D  XM3
timestamp 1746379951
transform 0 1 1941 -1 0 473
box -246 -1835 246 1835
<< labels >>
flabel metal1 122 1555 130 1564 0 FreeSans 400 0 0 0 VDD
port 0 nsew
flabel metal1 119 1343 127 1352 0 FreeSans 400 0 0 0 IN
port 1 nsew
flabel metal1 122 959 130 968 0 FreeSans 400 0 0 0 CKB
port 2 nsew
flabel metal1 120 466 128 475 0 FreeSans 400 0 0 0 CK
port 3 nsew
flabel metal1 123 -126 131 -117 0 FreeSans 400 0 0 0 VSS
port 4 nsew
flabel metal1 7220 701 7228 710 0 FreeSans 400 0 0 0 OUT
port 6 nsew
<< end >>
