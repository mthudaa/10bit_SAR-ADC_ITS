magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect 142 1527 168 1561
rect 202 1527 240 1561
rect 274 1527 312 1561
rect 346 1527 384 1561
rect 418 1527 456 1561
rect 490 1527 528 1561
rect 562 1527 600 1561
rect 634 1527 672 1561
rect 706 1527 744 1561
rect 778 1527 816 1561
rect 850 1527 888 1561
rect 922 1527 960 1561
rect 994 1527 1032 1561
rect 1066 1527 1104 1561
rect 1138 1527 1176 1561
rect 1210 1527 1248 1561
rect 1282 1527 1320 1561
rect 1354 1527 1392 1561
rect 1426 1527 1464 1561
rect 1498 1527 1536 1561
rect 1570 1527 1608 1561
rect 1642 1527 1680 1561
rect 1714 1527 1752 1561
rect 1786 1527 1824 1561
rect 1858 1527 1896 1561
rect 1930 1527 1968 1561
rect 2002 1527 2040 1561
rect 2074 1527 2112 1561
rect 2146 1527 2184 1561
rect 2218 1527 2256 1561
rect 2290 1527 2328 1561
rect 2362 1527 2400 1561
rect 2434 1527 2472 1561
rect 2506 1527 2544 1561
rect 2578 1527 2616 1561
rect 2650 1527 2688 1561
rect 2722 1527 2760 1561
rect 2794 1527 2832 1561
rect 2866 1527 2904 1561
rect 2938 1527 2976 1561
rect 3010 1527 3048 1561
rect 3082 1527 3120 1561
rect 3154 1527 3192 1561
rect 3226 1527 3264 1561
rect 3298 1527 3336 1561
rect 3370 1527 3408 1561
rect 3442 1527 3480 1561
rect 3514 1527 3552 1561
rect 3586 1527 3624 1561
rect 3658 1527 3696 1561
rect 3730 1527 3768 1561
rect 3802 1527 3840 1561
rect 3874 1527 3912 1561
rect 3946 1527 3984 1561
rect 4018 1527 4056 1561
rect 4090 1527 4128 1561
rect 4162 1527 4200 1561
rect 4234 1527 4272 1561
rect 4306 1527 4344 1561
rect 4378 1527 4416 1561
rect 4450 1527 4488 1561
rect 4522 1527 4560 1561
rect 4594 1527 4632 1561
rect 4666 1527 4704 1561
rect 4738 1527 4776 1561
rect 4810 1527 4848 1561
rect 4882 1527 4920 1561
rect 4954 1527 4992 1561
rect 5026 1527 5064 1561
rect 5098 1527 5136 1561
rect 5170 1527 5208 1561
rect 5242 1527 5280 1561
rect 5314 1527 5352 1561
rect 5386 1527 5424 1561
rect 5458 1527 5496 1561
rect 5530 1527 5568 1561
rect 5602 1527 5640 1561
rect 5674 1527 5712 1561
rect 5746 1527 5784 1561
rect 5818 1527 5856 1561
rect 5890 1527 5928 1561
rect 5962 1527 6000 1561
rect 6034 1527 6072 1561
rect 6106 1527 6144 1561
rect 6178 1527 6216 1561
rect 6250 1527 6288 1561
rect 6322 1527 6360 1561
rect 6394 1527 6432 1561
rect 6466 1527 6504 1561
rect 6538 1527 6576 1561
rect 6610 1527 6648 1561
rect 6682 1527 6720 1561
rect 6754 1527 6792 1561
rect 6826 1527 6864 1561
rect 6898 1527 6936 1561
rect 6970 1527 7008 1561
rect 7042 1527 7080 1561
rect 7114 1527 7152 1561
rect 7186 1527 7224 1561
rect 7258 1527 7296 1561
rect 7330 1527 7368 1561
rect 7402 1527 7440 1561
rect 7474 1527 7512 1561
rect 7546 1527 7584 1561
rect 7618 1527 7656 1561
rect 7690 1527 7728 1561
rect 7762 1527 7800 1561
rect 7834 1527 7872 1561
rect 7906 1527 7944 1561
rect 7978 1527 8016 1561
rect 8050 1527 8088 1561
rect 8122 1527 8160 1561
rect 8194 1527 8232 1561
rect 8266 1527 8304 1561
rect 8338 1527 8376 1561
rect 8410 1527 8448 1561
rect 8482 1527 8520 1561
rect 8554 1527 8592 1561
rect 8626 1527 8664 1561
rect 8698 1527 8736 1561
rect 8770 1527 8808 1561
rect 8842 1527 8880 1561
rect 8914 1527 8940 1561
rect 142 -123 148 -89
rect 182 -123 220 -89
rect 254 -123 292 -89
rect 326 -123 364 -89
rect 398 -123 436 -89
rect 470 -123 508 -89
rect 542 -123 580 -89
rect 614 -123 652 -89
rect 686 -123 724 -89
rect 758 -123 796 -89
rect 830 -123 868 -89
rect 902 -123 940 -89
rect 974 -123 1012 -89
rect 1046 -123 1084 -89
rect 1118 -123 1156 -89
rect 1190 -123 1228 -89
rect 1262 -123 1300 -89
rect 1334 -123 1372 -89
rect 1406 -123 1444 -89
rect 1478 -123 1516 -89
rect 1550 -123 1588 -89
rect 1622 -123 1660 -89
rect 1694 -123 1732 -89
rect 1766 -123 1804 -89
rect 1838 -123 1876 -89
rect 1910 -123 1948 -89
rect 1982 -123 2020 -89
rect 2054 -123 2092 -89
rect 2126 -123 2164 -89
rect 2198 -123 2236 -89
rect 2270 -123 2308 -89
rect 2342 -123 2380 -89
rect 2414 -123 2452 -89
rect 2486 -123 2524 -89
rect 2558 -123 2596 -89
rect 2630 -123 2668 -89
rect 2702 -123 2740 -89
rect 2774 -123 2812 -89
rect 2846 -123 2884 -89
rect 2918 -123 2956 -89
rect 2990 -123 3028 -89
rect 3062 -123 3100 -89
rect 3134 -123 3172 -89
rect 3206 -123 3244 -89
rect 3278 -123 3316 -89
rect 3350 -123 3388 -89
rect 3422 -123 3460 -89
rect 3494 -123 3532 -89
rect 3566 -123 3604 -89
rect 3638 -123 3676 -89
rect 3710 -123 3748 -89
rect 3782 -123 3820 -89
rect 3854 -123 3892 -89
rect 3926 -123 3964 -89
rect 3998 -123 4036 -89
rect 4070 -123 4108 -89
rect 4142 -123 4180 -89
rect 4214 -123 4252 -89
rect 4286 -123 4324 -89
rect 4358 -123 4396 -89
rect 4430 -123 4468 -89
rect 4502 -123 4540 -89
rect 4574 -123 4580 -89
<< viali >>
rect 168 1527 202 1561
rect 240 1527 274 1561
rect 312 1527 346 1561
rect 384 1527 418 1561
rect 456 1527 490 1561
rect 528 1527 562 1561
rect 600 1527 634 1561
rect 672 1527 706 1561
rect 744 1527 778 1561
rect 816 1527 850 1561
rect 888 1527 922 1561
rect 960 1527 994 1561
rect 1032 1527 1066 1561
rect 1104 1527 1138 1561
rect 1176 1527 1210 1561
rect 1248 1527 1282 1561
rect 1320 1527 1354 1561
rect 1392 1527 1426 1561
rect 1464 1527 1498 1561
rect 1536 1527 1570 1561
rect 1608 1527 1642 1561
rect 1680 1527 1714 1561
rect 1752 1527 1786 1561
rect 1824 1527 1858 1561
rect 1896 1527 1930 1561
rect 1968 1527 2002 1561
rect 2040 1527 2074 1561
rect 2112 1527 2146 1561
rect 2184 1527 2218 1561
rect 2256 1527 2290 1561
rect 2328 1527 2362 1561
rect 2400 1527 2434 1561
rect 2472 1527 2506 1561
rect 2544 1527 2578 1561
rect 2616 1527 2650 1561
rect 2688 1527 2722 1561
rect 2760 1527 2794 1561
rect 2832 1527 2866 1561
rect 2904 1527 2938 1561
rect 2976 1527 3010 1561
rect 3048 1527 3082 1561
rect 3120 1527 3154 1561
rect 3192 1527 3226 1561
rect 3264 1527 3298 1561
rect 3336 1527 3370 1561
rect 3408 1527 3442 1561
rect 3480 1527 3514 1561
rect 3552 1527 3586 1561
rect 3624 1527 3658 1561
rect 3696 1527 3730 1561
rect 3768 1527 3802 1561
rect 3840 1527 3874 1561
rect 3912 1527 3946 1561
rect 3984 1527 4018 1561
rect 4056 1527 4090 1561
rect 4128 1527 4162 1561
rect 4200 1527 4234 1561
rect 4272 1527 4306 1561
rect 4344 1527 4378 1561
rect 4416 1527 4450 1561
rect 4488 1527 4522 1561
rect 4560 1527 4594 1561
rect 4632 1527 4666 1561
rect 4704 1527 4738 1561
rect 4776 1527 4810 1561
rect 4848 1527 4882 1561
rect 4920 1527 4954 1561
rect 4992 1527 5026 1561
rect 5064 1527 5098 1561
rect 5136 1527 5170 1561
rect 5208 1527 5242 1561
rect 5280 1527 5314 1561
rect 5352 1527 5386 1561
rect 5424 1527 5458 1561
rect 5496 1527 5530 1561
rect 5568 1527 5602 1561
rect 5640 1527 5674 1561
rect 5712 1527 5746 1561
rect 5784 1527 5818 1561
rect 5856 1527 5890 1561
rect 5928 1527 5962 1561
rect 6000 1527 6034 1561
rect 6072 1527 6106 1561
rect 6144 1527 6178 1561
rect 6216 1527 6250 1561
rect 6288 1527 6322 1561
rect 6360 1527 6394 1561
rect 6432 1527 6466 1561
rect 6504 1527 6538 1561
rect 6576 1527 6610 1561
rect 6648 1527 6682 1561
rect 6720 1527 6754 1561
rect 6792 1527 6826 1561
rect 6864 1527 6898 1561
rect 6936 1527 6970 1561
rect 7008 1527 7042 1561
rect 7080 1527 7114 1561
rect 7152 1527 7186 1561
rect 7224 1527 7258 1561
rect 7296 1527 7330 1561
rect 7368 1527 7402 1561
rect 7440 1527 7474 1561
rect 7512 1527 7546 1561
rect 7584 1527 7618 1561
rect 7656 1527 7690 1561
rect 7728 1527 7762 1561
rect 7800 1527 7834 1561
rect 7872 1527 7906 1561
rect 7944 1527 7978 1561
rect 8016 1527 8050 1561
rect 8088 1527 8122 1561
rect 8160 1527 8194 1561
rect 8232 1527 8266 1561
rect 8304 1527 8338 1561
rect 8376 1527 8410 1561
rect 8448 1527 8482 1561
rect 8520 1527 8554 1561
rect 8592 1527 8626 1561
rect 8664 1527 8698 1561
rect 8736 1527 8770 1561
rect 8808 1527 8842 1561
rect 8880 1527 8914 1561
rect 148 -123 182 -89
rect 220 -123 254 -89
rect 292 -123 326 -89
rect 364 -123 398 -89
rect 436 -123 470 -89
rect 508 -123 542 -89
rect 580 -123 614 -89
rect 652 -123 686 -89
rect 724 -123 758 -89
rect 796 -123 830 -89
rect 868 -123 902 -89
rect 940 -123 974 -89
rect 1012 -123 1046 -89
rect 1084 -123 1118 -89
rect 1156 -123 1190 -89
rect 1228 -123 1262 -89
rect 1300 -123 1334 -89
rect 1372 -123 1406 -89
rect 1444 -123 1478 -89
rect 1516 -123 1550 -89
rect 1588 -123 1622 -89
rect 1660 -123 1694 -89
rect 1732 -123 1766 -89
rect 1804 -123 1838 -89
rect 1876 -123 1910 -89
rect 1948 -123 1982 -89
rect 2020 -123 2054 -89
rect 2092 -123 2126 -89
rect 2164 -123 2198 -89
rect 2236 -123 2270 -89
rect 2308 -123 2342 -89
rect 2380 -123 2414 -89
rect 2452 -123 2486 -89
rect 2524 -123 2558 -89
rect 2596 -123 2630 -89
rect 2668 -123 2702 -89
rect 2740 -123 2774 -89
rect 2812 -123 2846 -89
rect 2884 -123 2918 -89
rect 2956 -123 2990 -89
rect 3028 -123 3062 -89
rect 3100 -123 3134 -89
rect 3172 -123 3206 -89
rect 3244 -123 3278 -89
rect 3316 -123 3350 -89
rect 3388 -123 3422 -89
rect 3460 -123 3494 -89
rect 3532 -123 3566 -89
rect 3604 -123 3638 -89
rect 3676 -123 3710 -89
rect 3748 -123 3782 -89
rect 3820 -123 3854 -89
rect 3892 -123 3926 -89
rect 3964 -123 3998 -89
rect 4036 -123 4070 -89
rect 4108 -123 4142 -89
rect 4180 -123 4214 -89
rect 4252 -123 4286 -89
rect 4324 -123 4358 -89
rect 4396 -123 4430 -89
rect 4468 -123 4502 -89
rect 4540 -123 4574 -89
<< metal1 >>
rect 106 1561 8976 1597
rect 106 1527 168 1561
rect 202 1527 240 1561
rect 274 1527 312 1561
rect 346 1527 384 1561
rect 418 1527 456 1561
rect 490 1527 528 1561
rect 562 1527 600 1561
rect 634 1527 672 1561
rect 706 1527 744 1561
rect 778 1527 816 1561
rect 850 1527 888 1561
rect 922 1527 960 1561
rect 994 1527 1032 1561
rect 1066 1527 1104 1561
rect 1138 1527 1176 1561
rect 1210 1527 1248 1561
rect 1282 1527 1320 1561
rect 1354 1527 1392 1561
rect 1426 1527 1464 1561
rect 1498 1527 1536 1561
rect 1570 1527 1608 1561
rect 1642 1527 1680 1561
rect 1714 1527 1752 1561
rect 1786 1527 1824 1561
rect 1858 1527 1896 1561
rect 1930 1527 1968 1561
rect 2002 1527 2040 1561
rect 2074 1527 2112 1561
rect 2146 1527 2184 1561
rect 2218 1527 2256 1561
rect 2290 1527 2328 1561
rect 2362 1527 2400 1561
rect 2434 1527 2472 1561
rect 2506 1527 2544 1561
rect 2578 1527 2616 1561
rect 2650 1527 2688 1561
rect 2722 1527 2760 1561
rect 2794 1527 2832 1561
rect 2866 1527 2904 1561
rect 2938 1527 2976 1561
rect 3010 1527 3048 1561
rect 3082 1527 3120 1561
rect 3154 1527 3192 1561
rect 3226 1527 3264 1561
rect 3298 1527 3336 1561
rect 3370 1527 3408 1561
rect 3442 1527 3480 1561
rect 3514 1527 3552 1561
rect 3586 1527 3624 1561
rect 3658 1527 3696 1561
rect 3730 1527 3768 1561
rect 3802 1527 3840 1561
rect 3874 1527 3912 1561
rect 3946 1527 3984 1561
rect 4018 1527 4056 1561
rect 4090 1527 4128 1561
rect 4162 1527 4200 1561
rect 4234 1527 4272 1561
rect 4306 1527 4344 1561
rect 4378 1527 4416 1561
rect 4450 1527 4488 1561
rect 4522 1527 4560 1561
rect 4594 1527 4632 1561
rect 4666 1527 4704 1561
rect 4738 1527 4776 1561
rect 4810 1527 4848 1561
rect 4882 1527 4920 1561
rect 4954 1527 4992 1561
rect 5026 1527 5064 1561
rect 5098 1527 5136 1561
rect 5170 1527 5208 1561
rect 5242 1527 5280 1561
rect 5314 1527 5352 1561
rect 5386 1527 5424 1561
rect 5458 1527 5496 1561
rect 5530 1527 5568 1561
rect 5602 1527 5640 1561
rect 5674 1527 5712 1561
rect 5746 1527 5784 1561
rect 5818 1527 5856 1561
rect 5890 1527 5928 1561
rect 5962 1527 6000 1561
rect 6034 1527 6072 1561
rect 6106 1527 6144 1561
rect 6178 1527 6216 1561
rect 6250 1527 6288 1561
rect 6322 1527 6360 1561
rect 6394 1527 6432 1561
rect 6466 1527 6504 1561
rect 6538 1527 6576 1561
rect 6610 1527 6648 1561
rect 6682 1527 6720 1561
rect 6754 1527 6792 1561
rect 6826 1527 6864 1561
rect 6898 1527 6936 1561
rect 6970 1527 7008 1561
rect 7042 1527 7080 1561
rect 7114 1527 7152 1561
rect 7186 1527 7224 1561
rect 7258 1527 7296 1561
rect 7330 1527 7368 1561
rect 7402 1527 7440 1561
rect 7474 1527 7512 1561
rect 7546 1527 7584 1561
rect 7618 1527 7656 1561
rect 7690 1527 7728 1561
rect 7762 1527 7800 1561
rect 7834 1527 7872 1561
rect 7906 1527 7944 1561
rect 7978 1527 8016 1561
rect 8050 1527 8088 1561
rect 8122 1527 8160 1561
rect 8194 1527 8232 1561
rect 8266 1527 8304 1561
rect 8338 1527 8376 1561
rect 8410 1527 8448 1561
rect 8482 1527 8520 1561
rect 8554 1527 8592 1561
rect 8626 1527 8664 1561
rect 8698 1527 8736 1561
rect 8770 1527 8808 1561
rect 8842 1527 8880 1561
rect 8914 1527 8976 1561
rect 106 1521 8976 1527
rect 325 1447 8757 1521
rect 106 1377 284 1401
rect 106 1325 176 1377
rect 228 1325 284 1377
rect 106 1301 284 1325
rect 337 1061 8757 1255
rect 106 915 284 1015
rect 106 569 8976 869
rect 106 423 284 523
rect 316 183 4406 377
rect 166 113 284 137
rect 166 61 176 113
rect 228 61 284 113
rect 166 37 284 61
rect 316 -83 4406 -9
rect 106 -89 8976 -83
rect 106 -123 148 -89
rect 182 -123 220 -89
rect 254 -123 292 -89
rect 326 -123 364 -89
rect 398 -123 436 -89
rect 470 -123 508 -89
rect 542 -123 580 -89
rect 614 -123 652 -89
rect 686 -123 724 -89
rect 758 -123 796 -89
rect 830 -123 868 -89
rect 902 -123 940 -89
rect 974 -123 1012 -89
rect 1046 -123 1084 -89
rect 1118 -123 1156 -89
rect 1190 -123 1228 -89
rect 1262 -123 1300 -89
rect 1334 -123 1372 -89
rect 1406 -123 1444 -89
rect 1478 -123 1516 -89
rect 1550 -123 1588 -89
rect 1622 -123 1660 -89
rect 1694 -123 1732 -89
rect 1766 -123 1804 -89
rect 1838 -123 1876 -89
rect 1910 -123 1948 -89
rect 1982 -123 2020 -89
rect 2054 -123 2092 -89
rect 2126 -123 2164 -89
rect 2198 -123 2236 -89
rect 2270 -123 2308 -89
rect 2342 -123 2380 -89
rect 2414 -123 2452 -89
rect 2486 -123 2524 -89
rect 2558 -123 2596 -89
rect 2630 -123 2668 -89
rect 2702 -123 2740 -89
rect 2774 -123 2812 -89
rect 2846 -123 2884 -89
rect 2918 -123 2956 -89
rect 2990 -123 3028 -89
rect 3062 -123 3100 -89
rect 3134 -123 3172 -89
rect 3206 -123 3244 -89
rect 3278 -123 3316 -89
rect 3350 -123 3388 -89
rect 3422 -123 3460 -89
rect 3494 -123 3532 -89
rect 3566 -123 3604 -89
rect 3638 -123 3676 -89
rect 3710 -123 3748 -89
rect 3782 -123 3820 -89
rect 3854 -123 3892 -89
rect 3926 -123 3964 -89
rect 3998 -123 4036 -89
rect 4070 -123 4108 -89
rect 4142 -123 4180 -89
rect 4214 -123 4252 -89
rect 4286 -123 4324 -89
rect 4358 -123 4396 -89
rect 4430 -123 4468 -89
rect 4502 -123 4540 -89
rect 4574 -123 8976 -89
rect 106 -159 8976 -123
<< via1 >>
rect 176 1325 228 1377
rect 176 61 228 113
<< metal2 >>
rect 176 1377 228 1411
rect 176 113 228 1325
rect 176 27 228 61
use sky130_fd_pr__nfet_01v8_MKNP2D  sky130_fd_pr__nfet_01v8_MKNP2D_0
timestamp 1750100919
transform 0 1 2361 -1 0 87
box -236 -2245 236 2245
use sky130_fd_pr__pfet_01v8_C9QZQZ  sky130_fd_pr__pfet_01v8_C9QZQZ_0
timestamp 1750100919
transform 0 1 4541 -1 0 965
box -246 -4435 246 4435
use sky130_fd_pr__pfet_01v8_C9QZQZ  XM1
timestamp 1750100919
transform 0 1 4541 -1 0 1351
box -246 -4435 246 4435
use sky130_fd_pr__nfet_01v8_MKNP2D  XM3
timestamp 1750100919
transform 0 1 2361 -1 0 473
box -236 -2245 236 2245
<< labels >>
flabel metal1 s 120 1555 128 1563 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 117 1345 122 1350 0 FreeSans 500 0 0 0 IN
port 2 nsew
flabel metal1 s 120 961 125 966 0 FreeSans 500 0 0 0 CKB
port 3 nsew
flabel metal1 s 120 469 125 474 0 FreeSans 500 0 0 0 CK
port 4 nsew
flabel metal1 s 122 -124 127 -119 0 FreeSans 500 0 0 0 VSS
port 5 nsew
flabel metal1 s 8943 715 8948 720 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
