magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< metal1 >>
rect -1094 -22116 -38 -22090
rect -1094 -22168 -1072 -22116
rect -1020 -22168 -1008 -22116
rect -956 -22168 -38 -22116
rect -1094 -22194 -38 -22168
rect 47481 -22116 48486 -22090
rect 47481 -22168 48348 -22116
rect 48400 -22168 48412 -22116
rect 48464 -22168 48486 -22116
rect 47481 -22194 48486 -22168
rect 45426 -22324 45546 -22298
rect 45426 -22376 45460 -22324
rect 45512 -22376 45546 -22324
rect 45426 -22402 45546 -22376
rect 40620 -22532 40740 -22506
rect 40620 -22584 40654 -22532
rect 40706 -22584 40740 -22532
rect 40620 -22610 40740 -22584
rect 35818 -22740 35938 -22714
rect 35818 -22792 35852 -22740
rect 35904 -22792 35938 -22740
rect 35818 -22818 35938 -22792
rect 31016 -22948 31136 -22922
rect 31016 -23000 31050 -22948
rect 31102 -23000 31136 -22948
rect 31016 -23026 31136 -23000
rect 26219 -23156 26339 -23130
rect 26219 -23208 26253 -23156
rect 26305 -23208 26339 -23156
rect 26219 -23234 26339 -23208
rect 21412 -23364 21532 -23338
rect 21412 -23416 21446 -23364
rect 21498 -23416 21532 -23364
rect 21412 -23442 21532 -23416
rect 16612 -23572 16732 -23546
rect 16612 -23624 16646 -23572
rect 16698 -23624 16732 -23572
rect 16612 -23650 16732 -23624
rect 11808 -23780 11928 -23754
rect 11808 -23832 11842 -23780
rect 11894 -23832 11928 -23780
rect 11808 -23858 11928 -23832
rect 7006 -23988 7126 -23962
rect 7006 -24040 7040 -23988
rect 7092 -24040 7126 -23988
rect 7006 -24066 7126 -24040
rect 2204 -24196 2324 -24170
rect 2204 -24248 2238 -24196
rect 2290 -24248 2324 -24196
rect 2204 -24274 2324 -24248
rect 4128 -39935 4228 -39795
rect 4328 -39935 4428 -39595
rect 8930 -39935 9030 -39795
rect 9130 -39935 9230 -39595
rect 13732 -39935 13832 -39799
rect 13932 -39935 14032 -39595
rect 18534 -39935 18634 -39795
rect 18734 -39935 18834 -39595
rect 23336 -39935 23436 -39795
rect 23536 -39935 23636 -39595
rect 28138 -39935 28238 -39795
rect 28338 -39935 28438 -39595
rect 32940 -39935 33040 -39795
rect 33140 -39935 33240 -39595
rect 37742 -39935 37842 -39795
rect 37942 -39935 38042 -39595
rect 42544 -39935 42644 -39795
rect 42744 -39935 42844 -39595
rect 47346 -39935 47446 -39795
rect 47546 -39935 47646 -39595
<< via1 >>
rect -1072 -22168 -1020 -22116
rect -1008 -22168 -956 -22116
rect 48348 -22168 48400 -22116
rect 48412 -22168 48464 -22116
rect 45460 -22376 45512 -22324
rect 40654 -22584 40706 -22532
rect 35852 -22792 35904 -22740
rect 31050 -23000 31102 -22948
rect 26253 -23208 26305 -23156
rect 21446 -23416 21498 -23364
rect 16646 -23624 16698 -23572
rect 11842 -23832 11894 -23780
rect 7040 -24040 7092 -23988
rect 2238 -24248 2290 -24196
<< metal2 >>
rect -1084 -22116 -944 -22080
rect -1084 -22168 -1072 -22116
rect -1020 -22168 -1008 -22116
rect -956 -22168 -944 -22116
rect -1084 -39295 -944 -22168
rect -804 -38295 -664 -22090
rect -524 -38095 -384 -22090
rect 45436 -22324 45536 -22288
rect 45436 -22376 45460 -22324
rect 45512 -22376 45536 -22324
rect 40630 -22532 40730 -22496
rect 40630 -22584 40654 -22532
rect 40706 -22584 40730 -22532
rect 35828 -22740 35928 -22704
rect 35828 -22792 35852 -22740
rect 35904 -22792 35928 -22740
rect 31026 -22948 31126 -22912
rect 31026 -23000 31050 -22948
rect 31102 -23000 31126 -22948
rect 26229 -23156 26329 -23120
rect 26229 -23208 26253 -23156
rect 26305 -23208 26329 -23156
rect 21422 -23364 21522 -23328
rect 21422 -23416 21446 -23364
rect 21498 -23416 21522 -23364
rect 16622 -23572 16722 -23536
rect 16622 -23624 16646 -23572
rect 16698 -23624 16722 -23572
rect 11818 -23780 11918 -23744
rect 11818 -23832 11842 -23780
rect 11894 -23832 11918 -23780
rect 7016 -23988 7116 -23952
rect 7016 -24040 7040 -23988
rect 7092 -24040 7116 -23988
rect 2214 -24196 2314 -24160
rect 2214 -24248 2238 -24196
rect 2290 -24248 2314 -24196
rect 2214 -24514 2314 -24248
rect 7016 -25790 7116 -24040
rect 11818 -27066 11918 -23832
rect 16622 -28342 16722 -23624
rect 21422 -29618 21522 -23416
rect 26229 -30894 26329 -23208
rect 31026 -32170 31126 -23000
rect 35828 -33446 35928 -22792
rect 40630 -34722 40730 -22584
rect 45436 -35998 45536 -22376
rect 47776 -38095 47916 -22090
rect -524 -38195 -46 -38095
rect 47392 -38195 47916 -38095
rect 48056 -38295 48196 -22090
rect -804 -38395 -63 -38295
rect 47337 -38395 48196 -38295
rect 48336 -22116 48476 -22080
rect 48336 -22168 48348 -22116
rect 48400 -22168 48412 -22116
rect 48464 -22168 48476 -22116
rect 48336 -39295 48476 -22168
rect -1084 -39395 -129 -39295
rect 47347 -39395 48476 -39295
<< metal4 >>
rect 1621 14830 45489 14926
use cdac_sw_10b  cdac_sw_10b_0
timestamp 1750100919
transform 0 -1 4488 1 0 -39416
box -519 -43168 15012 4742
use x10b_cap_array  x10b_cap_array_0
timestamp 1750100919
transform 1 0 44991 0 1 13844
box -45174 -38128 2594 1082
<< labels >>
flabel metal2 s -471 -38074 -431 -38034 0 FreeSans 1000 0 0 0 VSS
port 1 nsew
flabel metal2 s -756 -38069 -716 -38029 0 FreeSans 1000 0 0 0 VDD
port 2 nsew
flabel metal2 s -1044 -38074 -1004 -38034 0 FreeSans 1000 0 0 0 VCM
port 3 nsew
flabel metal1 s 4160 -39905 4200 -39865 0 FreeSans 1000 0 0 0 SW_IN[0]
port 4 nsew
flabel metal1 s 8957 -39902 8997 -39862 0 FreeSans 1000 0 0 0 SW_IN[1]
port 5 nsew
flabel metal1 s 13755 -39914 13795 -39874 0 FreeSans 1000 0 0 0 SW_IN[2]
port 6 nsew
flabel metal1 s 18561 -39918 18601 -39878 0 FreeSans 1000 0 0 0 SW_IN[3]
port 7 nsew
flabel metal1 s 23354 -39923 23394 -39883 0 FreeSans 1000 0 0 0 SW_IN[4]
port 8 nsew
flabel metal1 s 28164 -39914 28204 -39874 0 FreeSans 1000 0 0 0 SW_IN[5]
port 9 nsew
flabel metal1 s 32969 -39916 33009 -39876 0 FreeSans 1000 0 0 0 SW_IN[6]
port 10 nsew
flabel metal1 s 37770 -39911 37810 -39871 0 FreeSans 1000 0 0 0 SW_IN[7]
port 11 nsew
flabel metal1 s 42576 -39911 42616 -39871 0 FreeSans 1000 0 0 0 SW_IN[8]
port 12 nsew
flabel metal1 s 47374 -39910 47414 -39870 0 FreeSans 1000 0 0 0 SW_IN[9]
port 13 nsew
flabel metal1 s 4355 -39667 4395 -39627 0 FreeSans 1000 0 0 0 CF[0]
port 14 nsew
flabel metal1 s 9157 -39658 9197 -39618 0 FreeSans 1000 0 0 0 CF[1]
port 15 nsew
flabel metal1 s 13962 -39657 14002 -39617 0 FreeSans 1000 0 0 0 CF[2]
port 16 nsew
flabel metal1 s 18760 -39671 18800 -39631 0 FreeSans 1000 0 0 0 CF[3]
port 17 nsew
flabel metal1 s 23565 -39662 23605 -39622 0 FreeSans 1000 0 0 0 CF[4]
port 18 nsew
flabel metal1 s 28367 -39661 28407 -39621 0 FreeSans 1000 0 0 0 CF[5]
port 19 nsew
flabel metal1 s 33165 -39670 33205 -39630 0 FreeSans 1000 0 0 0 CF[6]
port 20 nsew
flabel metal1 s 37970 -39663 38010 -39623 0 FreeSans 1000 0 0 0 CF[7]
port 21 nsew
flabel metal1 s 42769 -39670 42809 -39630 0 FreeSans 1000 0 0 0 CF[8]
port 22 nsew
flabel metal1 s 47575 -39663 47615 -39623 0 FreeSans 1000 0 0 0 CF[9]
port 23 nsew
flabel metal4 s 1621 14830 1717 14926 0 FreeSans 1000 0 0 0 VC
port 24 nsew
<< end >>
