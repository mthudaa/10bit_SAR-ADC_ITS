magic
tech sky130A
magscale 1 2
timestamp 1749307785
<< error_p >>
rect -29 791 29 797
rect -29 757 -17 791
rect -29 751 29 757
<< pwell >>
rect -211 -929 211 929
<< nmos >>
rect -15 -781 15 719
<< ndiff >>
rect -73 707 -15 719
rect -73 -769 -61 707
rect -27 -769 -15 707
rect -73 -781 -15 -769
rect 15 707 73 719
rect 15 -769 27 707
rect 61 -769 73 707
rect 15 -781 73 -769
<< ndiffc >>
rect -61 -769 -27 707
rect 27 -769 61 707
<< psubdiff >>
rect -175 859 -79 893
rect 79 859 175 893
rect -175 797 -141 859
rect 141 797 175 859
rect -175 -859 -141 -797
rect 141 -859 175 -797
rect -175 -893 -79 -859
rect 79 -893 175 -859
<< psubdiffcont >>
rect -79 859 79 893
rect -175 -797 -141 797
rect 141 -797 175 797
rect -79 -893 79 -859
<< poly >>
rect -33 791 33 807
rect -33 757 -17 791
rect 17 757 33 791
rect -33 741 33 757
rect -15 719 15 741
rect -15 -807 15 -781
<< polycont >>
rect -17 757 17 791
<< locali >>
rect -175 859 -79 893
rect 79 859 175 893
rect -175 797 -141 859
rect 141 797 175 859
rect -33 757 -17 791
rect 17 757 33 791
rect -61 707 -27 723
rect -61 -785 -27 -769
rect 27 707 61 723
rect 27 -785 61 -769
rect -175 -859 -141 -797
rect 141 -859 175 -797
rect -175 -893 -79 -859
rect 79 -893 175 -859
<< viali >>
rect -17 757 17 791
rect -61 -769 -27 707
rect 27 -769 61 707
<< metal1 >>
rect -29 791 29 797
rect -29 757 -17 791
rect 17 757 29 791
rect -29 751 29 757
rect -67 707 -21 719
rect -67 -769 -61 707
rect -27 -769 -21 707
rect -67 -781 -21 -769
rect 21 707 67 719
rect 21 -769 27 707
rect 61 -769 67 707
rect 21 -781 67 -769
<< properties >>
string FIXED_BBOX -158 -876 158 876
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 7.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
