magic
tech sky130A
magscale 1 2
timestamp 1748431729
<< error_s >>
rect -1815 -50381 -1687 -50379
rect -1768 -50426 -1752 -50410
rect -1750 -50426 -1734 -50410
rect -1784 -50442 -1718 -50426
rect -1768 -50444 -1734 -50442
rect -1784 -50460 -1718 -50444
rect -1768 -50476 -1752 -50460
rect -1750 -50476 -1734 -50460
<< dnwell >>
rect -803 -51536 -203 -50336
<< pwell >>
rect -2264 -52705 -826 -50313
<< psubdiff >>
rect -2154 -50381 -2130 -50347
rect -960 -50381 -936 -50347
rect -2230 -50447 -2196 -50423
rect -894 -50447 -860 -50423
rect -2230 -52595 -2196 -52571
rect -894 -52595 -860 -52571
rect -2154 -52671 -2130 -52637
rect -960 -52671 -936 -52637
<< psubdiffcont >>
rect -2130 -50381 -960 -50347
rect -2230 -52571 -2196 -50447
rect -894 -52571 -860 -50447
rect -2130 -52671 -960 -52637
<< poly >>
rect -1784 -50426 -1718 -50410
rect -1784 -50446 -1768 -50426
rect -1836 -50460 -1768 -50446
rect -1734 -50460 -1718 -50426
rect -1836 -50476 -1718 -50460
rect -1836 -50509 -1806 -50476
rect -1748 -50506 -1718 -50476
<< polycont >>
rect -1768 -50460 -1734 -50426
<< locali >>
rect -826 -50347 -180 -50313
rect -2230 -50381 -2130 -50347
rect -960 -50381 -860 -50347
rect -2230 -50447 -2196 -50381
rect -894 -50447 -860 -50381
rect -2230 -52637 -2196 -52571
rect -826 -51525 -792 -50347
rect -214 -51525 -180 -50347
rect -826 -51559 -180 -51525
rect -894 -52637 -860 -52571
rect -2230 -52671 -2130 -52637
rect -960 -52671 -860 -52637
<< metal1 >>
rect -324 -50490 -314 -50487
rect -2428 -50572 -2088 -50520
rect -2010 -50620 -2000 -50520
rect -1948 -50620 -1938 -50520
rect -645 -50536 -314 -50490
rect -324 -50539 -314 -50536
rect -262 -50539 -252 -50487
rect -2508 -50701 -1988 -50649
rect -2010 -51402 -2000 -51350
rect -1948 -51353 -1938 -51350
rect -1800 -51353 -1754 -51283
rect -1948 -51399 -1754 -51353
rect -758 -51377 -748 -50577
rect -696 -51377 -633 -50577
rect -591 -51287 -415 -50939
rect -591 -51339 -539 -51287
rect -487 -51339 -415 -51287
rect -373 -51339 -314 -50939
rect -262 -51339 -252 -50939
rect -1948 -51402 -1938 -51399
rect -430 -51432 -420 -51380
rect -368 -51432 -358 -51380
rect -2010 -52162 -2000 -52110
rect -1948 -52162 -1888 -52110
<< via1 >>
rect -2000 -50620 -1948 -50520
rect -314 -50539 -262 -50487
rect -2000 -51402 -1948 -51350
rect -748 -51377 -696 -50577
rect -539 -51339 -487 -51287
rect -314 -51339 -262 -50939
rect -420 -51432 -368 -51380
rect -2000 -52162 -1948 -52110
<< metal2 >>
rect -314 -50487 -262 -50477
rect -2000 -50520 -1948 -50510
rect -2000 -51350 -1948 -50620
rect -748 -50577 -696 -50567
rect -314 -50939 -262 -50539
rect -748 -51387 -696 -51377
rect -539 -51287 -487 -51277
rect -2000 -52110 -1948 -51402
rect -539 -51616 -487 -51339
rect -314 -51349 -262 -51339
rect -420 -51380 -368 -51370
rect -420 -51616 -368 -51432
rect -2000 -52172 -1948 -52162
use sky130_fd_pr__cap_mim_m3_1_9RRBT9  sky130_fd_pr__cap_mim_m3_1_9RRBT9_0
timestamp 1748343649
transform 1 0 -888 0 1 -57170
box -3410 -2680 3410 2680
use sky130_fd_pr__nfet_01v8_5KVWZD  sky130_fd_pr__nfet_01v8_5KVWZD_0
timestamp 1748343649
transform 1 0 -1069 0 1 -51509
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_5QF6Z6  sky130_fd_pr__nfet_01v8_5QF6Z6_0
timestamp 1748343649
transform 1 0 -1445 0 1 -51259
box -73 -776 73 776
use sky130_fd_pr__nfet_01v8_A4C6AH  sky130_fd_pr__nfet_01v8_A4C6AH_0
timestamp 1748431729
transform 1 0 -1821 0 1 -50909
box -73 -426 73 426
use sky130_fd_pr__nfet_01v8_A4C6AH  sky130_fd_pr__nfet_01v8_A4C6AH_1
timestamp 1748431729
transform 1 0 -1733 0 1 -50909
box -73 -426 73 426
use sky130_fd_pr__nfet_01v8_SM2BQK  sky130_fd_pr__nfet_01v8_SM2BQK_0
timestamp 1748361277
transform 1 0 -2021 0 1 -50601
box -73 -107 73 107
use sky130_fd_pr__pfet_01v8_27Q7PL  sky130_fd_pr__pfet_01v8_27Q7PL_0
timestamp 1748361277
transform 1 0 -2475 0 1 -50572
box -211 -259 211 259
use sky130_fd_pr__pfet_01v8_AQMHM9  sky130_fd_pr__pfet_01v8_AQMHM9_0
timestamp 1748351693
transform 1 0 -612 0 1 -50941
box -109 -498 109 464
use sky130_fd_pr__pfet_01v8_B3KWHC  sky130_fd_pr__pfet_01v8_B3KWHC_0
timestamp 1748351693
transform 1 0 -394 0 1 -51175
box -109 -264 109 298
use sky130_fd_pr__nfet_01v8_E5C6AZ  XM5
timestamp 1748347152
transform 1 0 -1821 0 1 -52310
box -73 -226 73 226
use sky130_fd_pr__nfet_01v8_5QF6Z6  XM8
timestamp 1748343649
transform 1 0 -1533 0 1 -51259
box -73 -776 73 776
use sky130_fd_pr__nfet_01v8_5KVWZD  XM10
timestamp 1748343649
transform 1 0 -1245 0 1 -51509
box -73 -1026 73 1026
use sky130_fd_pr__nfet_01v8_5KVWZD  XM11
timestamp 1748343649
transform 1 0 -1157 0 1 -51509
box -73 -1026 73 1026
<< end >>
