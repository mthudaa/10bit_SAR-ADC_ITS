magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect -17 369 -11 403
rect 23 369 61 403
rect 95 369 133 403
rect 167 369 205 403
rect 239 369 277 403
rect 311 369 349 403
rect 383 369 421 403
rect 455 369 493 403
rect 527 369 565 403
rect 599 369 637 403
rect 671 369 709 403
rect 743 369 781 403
rect 815 369 853 403
rect 887 369 925 403
rect 959 369 997 403
rect 1031 369 1069 403
rect 1103 369 1141 403
rect 1175 369 1213 403
rect 1247 369 1285 403
rect 1319 369 1357 403
rect 1391 369 1429 403
rect 1463 369 1501 403
rect 1535 369 1573 403
rect 1607 369 1645 403
rect 1679 369 1717 403
rect 1751 369 1789 403
rect 1823 369 1861 403
rect 1895 369 1933 403
rect 1967 369 2005 403
rect 2039 369 2077 403
rect 2111 369 2149 403
rect 2183 369 2221 403
rect 2255 369 2293 403
rect 2327 369 2365 403
rect 2399 369 2437 403
rect 2471 369 2509 403
rect 2543 369 2581 403
rect 2615 369 2653 403
rect 2687 369 2725 403
rect 2759 369 2797 403
rect 2831 369 2869 403
rect 2903 369 2941 403
rect 2975 369 3013 403
rect 3047 369 3085 403
rect 3119 369 3157 403
rect 3191 369 3229 403
rect 3263 369 3301 403
rect 3335 369 3373 403
rect 3407 369 3445 403
rect 3479 369 3517 403
rect 3551 369 3589 403
rect 3623 369 3661 403
rect 3695 369 3733 403
rect 3767 369 3805 403
rect 3839 369 3877 403
rect 3911 369 3949 403
rect 3983 369 4021 403
rect 4055 369 4093 403
rect 4127 369 4165 403
rect 4199 369 4237 403
rect 4271 369 4309 403
rect 4343 369 4381 403
rect 4415 369 4453 403
rect 4487 369 4525 403
rect 4559 369 4597 403
rect 4631 369 4669 403
rect 4703 369 4741 403
rect 4775 369 4813 403
rect 4847 369 4885 403
rect 4919 369 4957 403
rect 4991 369 5029 403
rect 5063 369 5101 403
rect 5135 369 5173 403
rect 5207 369 5245 403
rect 5279 369 5317 403
rect 5351 369 5357 403
rect 5429 -17 5459 17
rect 5493 -17 5531 17
rect 5565 -17 5603 17
rect 5637 -17 5675 17
rect 5709 -17 5747 17
rect 5781 -17 5819 17
rect 5853 -17 5891 17
rect 5925 -17 5963 17
rect 5997 -17 6035 17
rect 6069 -17 6107 17
rect 6141 -17 6179 17
rect 6213 -17 6251 17
rect 6285 -17 6323 17
rect 6357 -17 6395 17
rect 6429 -17 6467 17
rect 6501 -17 6539 17
rect 6573 -17 6611 17
rect 6645 -17 6683 17
rect 6717 -17 6755 17
rect 6789 -17 6827 17
rect 6861 -17 6899 17
rect 6933 -17 6971 17
rect 7005 -17 7043 17
rect 7077 -17 7115 17
rect 7149 -17 7187 17
rect 7221 -17 7259 17
rect 7293 -17 7331 17
rect 7365 -17 7403 17
rect 7437 -17 7475 17
rect 7509 -17 7547 17
rect 7581 -17 7619 17
rect 7653 -17 7691 17
rect 7725 -17 7763 17
rect 7797 -17 7835 17
rect 7869 -17 7907 17
rect 7941 -17 7979 17
rect 8013 -17 8051 17
rect 8085 -17 8123 17
rect 8157 -17 8187 17
<< viali >>
rect -11 369 23 403
rect 61 369 95 403
rect 133 369 167 403
rect 205 369 239 403
rect 277 369 311 403
rect 349 369 383 403
rect 421 369 455 403
rect 493 369 527 403
rect 565 369 599 403
rect 637 369 671 403
rect 709 369 743 403
rect 781 369 815 403
rect 853 369 887 403
rect 925 369 959 403
rect 997 369 1031 403
rect 1069 369 1103 403
rect 1141 369 1175 403
rect 1213 369 1247 403
rect 1285 369 1319 403
rect 1357 369 1391 403
rect 1429 369 1463 403
rect 1501 369 1535 403
rect 1573 369 1607 403
rect 1645 369 1679 403
rect 1717 369 1751 403
rect 1789 369 1823 403
rect 1861 369 1895 403
rect 1933 369 1967 403
rect 2005 369 2039 403
rect 2077 369 2111 403
rect 2149 369 2183 403
rect 2221 369 2255 403
rect 2293 369 2327 403
rect 2365 369 2399 403
rect 2437 369 2471 403
rect 2509 369 2543 403
rect 2581 369 2615 403
rect 2653 369 2687 403
rect 2725 369 2759 403
rect 2797 369 2831 403
rect 2869 369 2903 403
rect 2941 369 2975 403
rect 3013 369 3047 403
rect 3085 369 3119 403
rect 3157 369 3191 403
rect 3229 369 3263 403
rect 3301 369 3335 403
rect 3373 369 3407 403
rect 3445 369 3479 403
rect 3517 369 3551 403
rect 3589 369 3623 403
rect 3661 369 3695 403
rect 3733 369 3767 403
rect 3805 369 3839 403
rect 3877 369 3911 403
rect 3949 369 3983 403
rect 4021 369 4055 403
rect 4093 369 4127 403
rect 4165 369 4199 403
rect 4237 369 4271 403
rect 4309 369 4343 403
rect 4381 369 4415 403
rect 4453 369 4487 403
rect 4525 369 4559 403
rect 4597 369 4631 403
rect 4669 369 4703 403
rect 4741 369 4775 403
rect 4813 369 4847 403
rect 4885 369 4919 403
rect 4957 369 4991 403
rect 5029 369 5063 403
rect 5101 369 5135 403
rect 5173 369 5207 403
rect 5245 369 5279 403
rect 5317 369 5351 403
rect 5459 -17 5493 17
rect 5531 -17 5565 17
rect 5603 -17 5637 17
rect 5675 -17 5709 17
rect 5747 -17 5781 17
rect 5819 -17 5853 17
rect 5891 -17 5925 17
rect 5963 -17 5997 17
rect 6035 -17 6069 17
rect 6107 -17 6141 17
rect 6179 -17 6213 17
rect 6251 -17 6285 17
rect 6323 -17 6357 17
rect 6395 -17 6429 17
rect 6467 -17 6501 17
rect 6539 -17 6573 17
rect 6611 -17 6645 17
rect 6683 -17 6717 17
rect 6755 -17 6789 17
rect 6827 -17 6861 17
rect 6899 -17 6933 17
rect 6971 -17 7005 17
rect 7043 -17 7077 17
rect 7115 -17 7149 17
rect 7187 -17 7221 17
rect 7259 -17 7293 17
rect 7331 -17 7365 17
rect 7403 -17 7437 17
rect 7475 -17 7509 17
rect 7547 -17 7581 17
rect 7619 -17 7653 17
rect 7691 -17 7725 17
rect 7763 -17 7797 17
rect 7835 -17 7869 17
rect 7907 -17 7941 17
rect 7979 -17 8013 17
rect 8051 -17 8085 17
rect 8123 -17 8157 17
<< metal1 >>
rect -53 403 8223 439
rect -53 369 -11 403
rect 23 369 61 403
rect 95 369 133 403
rect 167 369 205 403
rect 239 369 277 403
rect 311 369 349 403
rect 383 369 421 403
rect 455 369 493 403
rect 527 369 565 403
rect 599 369 637 403
rect 671 369 709 403
rect 743 369 781 403
rect 815 369 853 403
rect 887 369 925 403
rect 959 369 997 403
rect 1031 369 1069 403
rect 1103 369 1141 403
rect 1175 369 1213 403
rect 1247 369 1285 403
rect 1319 369 1357 403
rect 1391 369 1429 403
rect 1463 369 1501 403
rect 1535 369 1573 403
rect 1607 369 1645 403
rect 1679 369 1717 403
rect 1751 369 1789 403
rect 1823 369 1861 403
rect 1895 369 1933 403
rect 1967 369 2005 403
rect 2039 369 2077 403
rect 2111 369 2149 403
rect 2183 369 2221 403
rect 2255 369 2293 403
rect 2327 369 2365 403
rect 2399 369 2437 403
rect 2471 369 2509 403
rect 2543 369 2581 403
rect 2615 369 2653 403
rect 2687 369 2725 403
rect 2759 369 2797 403
rect 2831 369 2869 403
rect 2903 369 2941 403
rect 2975 369 3013 403
rect 3047 369 3085 403
rect 3119 369 3157 403
rect 3191 369 3229 403
rect 3263 369 3301 403
rect 3335 369 3373 403
rect 3407 369 3445 403
rect 3479 369 3517 403
rect 3551 369 3589 403
rect 3623 369 3661 403
rect 3695 369 3733 403
rect 3767 369 3805 403
rect 3839 369 3877 403
rect 3911 369 3949 403
rect 3983 369 4021 403
rect 4055 369 4093 403
rect 4127 369 4165 403
rect 4199 369 4237 403
rect 4271 369 4309 403
rect 4343 369 4381 403
rect 4415 369 4453 403
rect 4487 369 4525 403
rect 4559 369 4597 403
rect 4631 369 4669 403
rect 4703 369 4741 403
rect 4775 369 4813 403
rect 4847 369 4885 403
rect 4919 369 4957 403
rect 4991 369 5029 403
rect 5063 369 5101 403
rect 5135 369 5173 403
rect 5207 369 5245 403
rect 5279 369 5317 403
rect 5351 369 8223 403
rect -53 363 8223 369
rect -53 323 7794 324
rect -53 290 8013 323
rect 166 289 8013 290
rect -53 143 125 243
rect 8045 143 8223 243
rect 166 63 8223 97
rect -53 17 8223 23
rect -53 -17 5459 17
rect 5493 -17 5531 17
rect 5565 -17 5603 17
rect 5637 -17 5675 17
rect 5709 -17 5747 17
rect 5781 -17 5819 17
rect 5853 -17 5891 17
rect 5925 -17 5963 17
rect 5997 -17 6035 17
rect 6069 -17 6107 17
rect 6141 -17 6179 17
rect 6213 -17 6251 17
rect 6285 -17 6323 17
rect 6357 -17 6395 17
rect 6429 -17 6467 17
rect 6501 -17 6539 17
rect 6573 -17 6611 17
rect 6645 -17 6683 17
rect 6717 -17 6755 17
rect 6789 -17 6827 17
rect 6861 -17 6899 17
rect 6933 -17 6971 17
rect 7005 -17 7043 17
rect 7077 -17 7115 17
rect 7149 -17 7187 17
rect 7221 -17 7259 17
rect 7293 -17 7331 17
rect 7365 -17 7403 17
rect 7437 -17 7475 17
rect 7509 -17 7547 17
rect 7581 -17 7619 17
rect 7653 -17 7691 17
rect 7725 -17 7763 17
rect 7797 -17 7835 17
rect 7869 -17 7907 17
rect 7941 -17 7979 17
rect 8013 -17 8051 17
rect 8085 -17 8123 17
rect 8157 -17 8223 17
rect -53 -53 8223 -17
use sky130_fd_pr__pfet_01v8_D9QVK3  XM1
timestamp 1750100919
transform 0 1 2670 -1 0 193
box -246 -2723 246 2723
use sky130_fd_pr__nfet_01v8_PHNS9E  XM2
timestamp 1750100919
transform 0 1 6808 -1 0 193
box -236 -1405 236 1405
<< labels >>
flabel metal1 s -39 391 -26 404 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s -34 -25 -21 -12 0 FreeSans 500 0 0 0 VSS
port 2 nsew
flabel metal1 s -40 303 -27 316 0 FreeSans 500 0 0 0 IN
port 3 nsew
flabel metal1 s -39 185 -26 198 0 FreeSans 500 0 0 0 SWP
port 4 nsew
flabel metal1 s 8196 186 8209 199 0 FreeSans 500 0 0 0 SWN
port 5 nsew
flabel metal1 s 8203 74 8216 87 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
