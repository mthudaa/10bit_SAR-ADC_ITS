magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect -17 369 1 403
rect 35 369 73 403
rect 107 369 145 403
rect 179 369 217 403
rect 251 369 289 403
rect 323 369 361 403
rect 395 369 433 403
rect 467 369 505 403
rect 539 369 577 403
rect 611 369 649 403
rect 683 369 721 403
rect 755 369 793 403
rect 827 369 865 403
rect 899 369 937 403
rect 971 369 1009 403
rect 1043 369 1081 403
rect 1115 369 1153 403
rect 1187 369 1225 403
rect 1259 369 1297 403
rect 1331 369 1369 403
rect 1403 369 1441 403
rect 1475 369 1513 403
rect 1547 369 1585 403
rect 1619 369 1657 403
rect 1691 369 1729 403
rect 1763 369 1801 403
rect 1835 369 1873 403
rect 1907 369 1945 403
rect 1979 369 2017 403
rect 2051 369 2089 403
rect 2123 369 2161 403
rect 2195 369 2233 403
rect 2267 369 2305 403
rect 2339 369 2377 403
rect 2411 369 2449 403
rect 2483 369 2521 403
rect 2555 369 2593 403
rect 2627 369 2665 403
rect 2699 369 2737 403
rect 2771 369 2789 403
rect 2861 -17 2873 17
rect 2907 -17 2945 17
rect 2979 -17 3017 17
rect 3051 -17 3089 17
rect 3123 -17 3161 17
rect 3195 -17 3233 17
rect 3267 -17 3305 17
rect 3339 -17 3377 17
rect 3411 -17 3449 17
rect 3483 -17 3521 17
rect 3555 -17 3593 17
rect 3627 -17 3665 17
rect 3699 -17 3737 17
rect 3771 -17 3809 17
rect 3843 -17 3881 17
rect 3915 -17 3953 17
rect 3987 -17 4025 17
rect 4059 -17 4097 17
rect 4131 -17 4169 17
rect 4203 -17 4241 17
rect 4275 -17 4313 17
rect 4347 -17 4359 17
<< viali >>
rect 1 369 35 403
rect 73 369 107 403
rect 145 369 179 403
rect 217 369 251 403
rect 289 369 323 403
rect 361 369 395 403
rect 433 369 467 403
rect 505 369 539 403
rect 577 369 611 403
rect 649 369 683 403
rect 721 369 755 403
rect 793 369 827 403
rect 865 369 899 403
rect 937 369 971 403
rect 1009 369 1043 403
rect 1081 369 1115 403
rect 1153 369 1187 403
rect 1225 369 1259 403
rect 1297 369 1331 403
rect 1369 369 1403 403
rect 1441 369 1475 403
rect 1513 369 1547 403
rect 1585 369 1619 403
rect 1657 369 1691 403
rect 1729 369 1763 403
rect 1801 369 1835 403
rect 1873 369 1907 403
rect 1945 369 1979 403
rect 2017 369 2051 403
rect 2089 369 2123 403
rect 2161 369 2195 403
rect 2233 369 2267 403
rect 2305 369 2339 403
rect 2377 369 2411 403
rect 2449 369 2483 403
rect 2521 369 2555 403
rect 2593 369 2627 403
rect 2665 369 2699 403
rect 2737 369 2771 403
rect 2873 -17 2907 17
rect 2945 -17 2979 17
rect 3017 -17 3051 17
rect 3089 -17 3123 17
rect 3161 -17 3195 17
rect 3233 -17 3267 17
rect 3305 -17 3339 17
rect 3377 -17 3411 17
rect 3449 -17 3483 17
rect 3521 -17 3555 17
rect 3593 -17 3627 17
rect 3665 -17 3699 17
rect 3737 -17 3771 17
rect 3809 -17 3843 17
rect 3881 -17 3915 17
rect 3953 -17 3987 17
rect 4025 -17 4059 17
rect 4097 -17 4131 17
rect 4169 -17 4203 17
rect 4241 -17 4275 17
rect 4313 -17 4347 17
<< metal1 >>
rect -53 403 4395 439
rect -53 369 1 403
rect 35 369 73 403
rect 107 369 145 403
rect 179 369 217 403
rect 251 369 289 403
rect 323 369 361 403
rect 395 369 433 403
rect 467 369 505 403
rect 539 369 577 403
rect 611 369 649 403
rect 683 369 721 403
rect 755 369 793 403
rect 827 369 865 403
rect 899 369 937 403
rect 971 369 1009 403
rect 1043 369 1081 403
rect 1115 369 1153 403
rect 1187 369 1225 403
rect 1259 369 1297 403
rect 1331 369 1369 403
rect 1403 369 1441 403
rect 1475 369 1513 403
rect 1547 369 1585 403
rect 1619 369 1657 403
rect 1691 369 1729 403
rect 1763 369 1801 403
rect 1835 369 1873 403
rect 1907 369 1945 403
rect 1979 369 2017 403
rect 2051 369 2089 403
rect 2123 369 2161 403
rect 2195 369 2233 403
rect 2267 369 2305 403
rect 2339 369 2377 403
rect 2411 369 2449 403
rect 2483 369 2521 403
rect 2555 369 2593 403
rect 2627 369 2665 403
rect 2699 369 2737 403
rect 2771 369 4395 403
rect -53 363 4395 369
rect -53 289 4185 323
rect -53 143 125 243
rect 4217 143 4395 243
rect 166 63 4395 97
rect -53 17 4395 23
rect -53 -17 2873 17
rect 2907 -17 2945 17
rect 2979 -17 3017 17
rect 3051 -17 3089 17
rect 3123 -17 3161 17
rect 3195 -17 3233 17
rect 3267 -17 3305 17
rect 3339 -17 3377 17
rect 3411 -17 3449 17
rect 3483 -17 3521 17
rect 3555 -17 3593 17
rect 3627 -17 3665 17
rect 3699 -17 3737 17
rect 3771 -17 3809 17
rect 3843 -17 3881 17
rect 3915 -17 3953 17
rect 3987 -17 4025 17
rect 4059 -17 4097 17
rect 4131 -17 4169 17
rect 4203 -17 4241 17
rect 4275 -17 4313 17
rect 4347 -17 4395 17
rect -53 -53 4395 -17
use sky130_fd_pr__pfet_01v8_SEQFW4  XM1
timestamp 1750100919
transform 0 1 1386 -1 0 193
box -246 -1439 246 1439
use sky130_fd_pr__nfet_01v8_A9PWNX  XM2
timestamp 1750100919
transform 0 1 3610 -1 0 193
box -236 -775 236 775
<< labels >>
flabel metal1 s -41 393 -32 401 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s -40 -9 -31 -1 0 FreeSans 500 0 0 0 VSS
port 2 nsew
flabel metal1 s -41 302 -32 310 0 FreeSans 500 0 0 0 IN
port 3 nsew
flabel metal1 s -38 189 -29 197 0 FreeSans 500 0 0 0 SWP
port 4 nsew
flabel metal1 s 4374 196 4383 204 0 FreeSans 500 0 0 0 SWN
port 5 nsew
flabel metal1 s 4371 76 4380 84 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
