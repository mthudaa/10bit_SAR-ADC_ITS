../mag/delay_gate_ori.pex.spice