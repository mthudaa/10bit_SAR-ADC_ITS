magic
tech sky130A
magscale 1 2
timestamp 1749226371
<< metal1 >>
rect -18 1178 2668 1276
rect 966 1061 976 1121
rect 1028 1061 1260 1121
rect 1070 941 1080 1001
rect 1132 941 1264 1001
rect 2623 935 2706 975
rect 1471 723 2706 763
rect 1759 644 2706 684
rect 1218 512 1228 608
rect 1324 512 1334 608
rect -18 8 1228 106
rect 1324 8 1334 106
<< via1 >>
rect 976 1061 1028 1121
rect 1080 941 1132 1001
rect 1228 512 1324 608
rect 1228 8 1324 106
<< metal2 >>
rect -18 356 34 1935
rect 86 505 138 2084
rect 976 1121 1028 1131
rect 976 1051 1028 1061
rect 1080 1001 1132 1011
rect 1080 931 1132 941
rect 1228 608 1324 618
rect 1228 106 1324 512
rect 1228 -2 1324 8
use pd_in  pd_in_0
timestamp 1749046477
transform 1 0 590 0 1 1212
box -618 -1214 552 1244
use pd_out  pd_out_0
timestamp 1749226129
transform 1 0 1190 0 1 610
box 0 -98 1516 666
<< labels >>
flabel metal1 401 1208 431 1238 0 FreeSans 400 0 0 0 VDD
port 0 nsew
flabel metal1 392 43 422 73 0 FreeSans 400 0 0 0 VSS
port 1 nsew
flabel metal2 -5 829 25 859 0 FreeSans 400 0 0 0 INP
port 2 nsew
flabel metal2 100 829 130 859 0 FreeSans 400 0 0 0 INN
port 3 nsew
flabel metal1 2672 941 2702 971 0 FreeSans 400 0 0 0 RDY
port 4 nsew
flabel metal1 2669 730 2699 760 0 FreeSans 400 0 0 0 OUTP
port 5 nsew
flabel metal1 2670 648 2700 678 0 FreeSans 400 0 0 0 OUTN
port 6 nsew
<< end >>
