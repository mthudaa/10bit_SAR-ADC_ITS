* PEX produced on Thu Jun 12 04:56:30 PM WIB 2025 using ./iic-pex.sh with m=2 and s=1
* NGSPICE file created from x10b_adc_pex.ext - technology: sky130A

.subckt x10b_adc_pex VCM EN VDDA VDDR CLK CKO DATA[8] DATA[7] DATA[6] DATA[5] DATA[4]
+ DATA[3] DATA[2] DATA[1] DATA[0] VINP VINN VSSR VSSA VSSD VDDD DATA[9]
X0 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=95.7 ps=1.0428k w=0.5 l=0.5
X5 a_68178_51635# sar10b_0.clk_div_0.COUNT\[0\] VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.168 ps=1.24 w=0.84 l=0.15
X6 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7 c1_25688_97972# m3_25356_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8 VSSA a_55121_59650# tdc_0.RDY VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.2997 pd=2.29 as=0.1554 ps=1.16 w=0.74 l=0.15
X9 a_12472_111642# sar10b_0.CF[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X10 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X11 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X12 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X13 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X14 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X15 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X16 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X17 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X18 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X19 VSSD sar10b_0.cyclic_flag_0.FINAL a_67209_55011# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X20 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=9.28 ps=101.12 w=0.5 l=0.5
X21 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=287.10001 ps=2.3628k w=1.5 l=0.5
X22 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X23 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=121.95275 ps=1.15351k w=0.42 l=1
X24 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X25 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X26 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X27 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[9] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X28 a_65643_71265# sar10b_0.net43 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X29 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X30 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X31 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X32 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X33 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X34 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X35 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X36 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X37 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=34.8 ps=286.39999 w=1.5 l=0.5
X38 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X39 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X40 VSSR sar10b_0.SWN[3] a_29939_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X41 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X42 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X43 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X44 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X45 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X46 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X47 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X48 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X49 sar10b_0.net16 a_66785_50875# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.203 ps=1.505 w=1.12 l=0.15
X50 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X51 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X52 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X53 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X54 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X55 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X56 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X57 VSSD a_65407_63634# sar10b_0.net43 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X58 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X59 a_62281_52347# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X60 a_64949_64916# a_64814_65014# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X61 VDDD a_61929_51311# a_62181_51440# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X62 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X63 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X64 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X65 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X66 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X67 VDDD sar10b_0.cyclic_flag_0.FINAL a_67055_68689# VDDD sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.147 ps=1.19 w=0.84 l=0.15
X68 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=5.8 ps=63.2 w=0.5 l=0.5
X69 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X70 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_108738# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X71 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=10.44 ps=113.76 w=0.5 l=0.5
X72 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X73 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X74 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X75 tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A a_51345_58977# VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X76 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X77 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X78 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X79 VSSD a_60690_49683# sar10b_0.net3 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X80 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X81 c1_45456_80052# m3_45124_80012# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X82 a_40248_111636# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X83 c1_n1140_47378# m3_n1472_47338# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X84 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X85 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X86 VDDD a_67084_53565# sar10b_0._17_ VDDD sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.3304 ps=2.83 w=1.12 l=0.15
X87 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=8.12 ps=88.48 w=0.5 l=0.5
X88 a_64149_60339# a_64085_60119# a_64071_60339# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X89 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X90 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X91 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X92 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X93 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X94 VSSD sar10b_0.net16 a_64620_65967# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X95 a_62899_55988# a_61921_55975# a_62697_56343# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X96 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X97 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X98 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X99 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X100 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X101 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X102 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X103 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X104 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X105 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X106 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=207.74103 ps=1.80017k w=1 l=1
X107 a_62185_64695# a_61395_64612# a_61677_64842# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X108 VSSD a_62181_51440# a_62139_51318# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X109 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X110 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X111 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X112 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X113 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X114 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X115 c1_45456_95732# m3_45124_95692# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X116 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X117 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X118 a_62131_67714# a_61153_67587# a_61929_67295# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X119 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X120 VDDD a_68169_64335# a_68421_64288# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X121 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X122 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X123 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X124 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X125 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X126 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X127 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X128 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X129 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=11.6 ps=126.4 w=0.5 l=0.5
X130 VDDD a_64831_56974# sar10b_0.net31 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X131 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X132 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X133 VSSR sar10b_0.SWN[4] a_25137_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X134 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X135 VSSD a_65733_59432# a_65691_59310# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X136 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X137 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X138 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X139 a_62949_56296# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X140 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X141 VDDD sar10b_0.net16 a_64725_68631# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X142 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X143 a_61589_50795# a_61454_50696# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X144 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X145 a_60747_61567# sar10b_0.net9 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X146 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X147 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y sar10b_0.CF[8] VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X148 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X149 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=4.64 ps=50.56 w=0.5 l=0.5
X150 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X151 VDDD a_65068_49569# sar10b_0._10_ VDDD sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.3304 ps=2.83 w=1.12 l=0.15
X152 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X153 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X154 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X155 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X156 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X157 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X158 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X159 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X160 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X161 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X162 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X163 VDDD sar10b_0.net22 a_68946_56639# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X164 VDDD a_64491_48621# sar10b_0.SWN[4] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X165 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=31.32 ps=257.76001 w=1.5 l=0.5
X166 a_60747_57571# sar10b_0.net6 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X167 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X168 VSSD sar10b_0.clk_div_0.COUNT\[2\] sar10b_0._15_ VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1443 ps=1.13 w=0.74 l=0.15
X169 VDDD a_66633_56639# a_66885_56768# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X170 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X171 VDDD sar10b_0.cyclic_flag_0.FINAL a_67209_68331# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X172 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X173 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X174 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=11.6 ps=126.4 w=0.5 l=0.5
X175 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X176 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X177 a_24259_5788# sar10b_0.SWN[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X178 a_67372_52833# sar10b_0._14_ VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.17738 pd=1.195 as=0.12607 ps=1.1 w=0.55 l=0.15
X179 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X180 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X181 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X182 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X183 a_62995_57320# a_62017_57307# a_62793_57675# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X184 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X185 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=20.88 ps=171.84 w=1.5 l=0.5
X186 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A a_41284_111642# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X187 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X188 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X189 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X190 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X191 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_110450# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X192 c1_4508_97972# m3_4176_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X193 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X194 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X195 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X196 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X197 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X198 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X199 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X200 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X201 a_68767_63980# a_68169_64335# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X202 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=4.64 ps=50.56 w=0.5 l=0.5
X203 VDDD sar10b_0.clknet_1_1__leaf_CLK a_65682_51977# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X204 a_65355_53949# sar10b_0.clknet_0_CLK VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X205 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X206 a_64492_67433# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=0.98 as=0.0735 ps=0.77 w=0.42 l=0.15
X207 c1_15804_97972# m3_15472_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X208 a_10731_113461# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X209 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X210 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X211 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X212 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X213 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X214 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X215 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X216 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X217 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X218 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X219 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X220 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X221 VSSR sar10b_0.SWP[3] a_29939_111781# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X222 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X223 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X224 a_66351_68634# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X225 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X226 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X227 c1_41220_97972# m3_40888_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X228 a_63045_57628# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X229 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X230 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X231 VSSD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X232 tdc_0.OUTP tdc_0.phase_detector_0.pd_out_0.B a_54372_59599# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X233 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X234 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X235 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X236 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X237 a_6634_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X238 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X239 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_109594# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X240 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X241 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X242 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y sar10b_0.CF[6] VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X243 c1_27100_21618# m3_26768_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X244 VDDD sar10b_0.clknet_0_CLK a_65355_53949# VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X245 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X246 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X247 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X248 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X249 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X250 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X251 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X252 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X253 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X254 c1_45456_42898# m3_45124_42858# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X255 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X256 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X257 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X258 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X259 VDDD sar10b_0.net3 a_66933_63063# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X260 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X261 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 a_9853_112162# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X262 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X263 sar10b_0.net29 a_60747_49953# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X264 a_68767_67976# a_68169_68331# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X265 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X266 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X267 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X268 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X269 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X270 a_68421_58960# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X271 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X272 VDDD sar10b_0._09_ a_65021_50292# VDDD sky130_fd_pr__pfet_01v8 ad=0.33483 pd=1.765 as=0.1703 ps=1.355 w=0.84 l=0.15
X273 a_66101_58256# a_65966_58354# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X274 a_61035_71265# sar10b_0.net39 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X275 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X276 VSSD sar10b_0.cyclic_flag_0.FINAL a_67142_68689# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1376 ps=1.14 w=0.64 l=0.15
X277 c1_n1140_87892# m3_n1472_87852# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X278 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X279 a_29061_108738# sar10b_0.SWP[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X280 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X281 VSSD a_65577_51311# sar10b_0.clknet_0_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X282 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X283 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X284 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X285 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X286 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_110450# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X287 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X288 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X289 DATA[3] a_68946_53975# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X290 a_63369_59007# a_62593_58639# a_62933_58787# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X291 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X292 a_54372_59599# tdc_0.OUTN VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X293 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X294 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X295 VSSD sar10b_0.cyclic_flag_0.FINAL a_67209_64335# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X296 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X297 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X298 VSSD sar10b_0.net16 a_66453_69663# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X299 a_63663_67678# a_63457_67583# a_62997_67299# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1218 ps=1.42 w=0.42 l=0.15
X300 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X301 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X302 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X303 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=6.96 ps=75.84 w=0.5 l=0.5
X304 a_62222_57356# a_62017_57307# a_61557_57735# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X305 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X306 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X307 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X308 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X309 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X310 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X311 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X312 c1_45456_65492# m3_45124_65452# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X313 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X314 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X315 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X316 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y sar10b_0.CF[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X317 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X318 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X319 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X320 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X321 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X322 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X323 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X324 a_62185_52707# a_61395_52624# a_61677_52854# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X325 CKO a_68562_71291# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X326 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X327 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X328 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X329 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X330 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X331 a_62038_66346# a_61609_66266# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X332 VDDR sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X333 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X334 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_109594# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X335 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=31.32 ps=257.76001 w=1.5 l=0.5
X336 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X337 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X338 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X339 a_66261_56703# a_66197_56924# a_66183_56703# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X340 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X341 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X342 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X343 c1_35572_21618# m3_35240_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X344 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X345 a_65983_64966# a_65385_64631# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X346 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X347 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X348 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X349 a_62277_53632# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X350 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X351 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X352 a_61557_57735# sar10b_0.net2 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X353 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X354 VSSD sar10b_0.net26 a_68946_65963# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X355 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X356 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X357 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X358 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X359 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X360 a_66453_69663# a_66389_69443# a_66375_69663# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X361 a_61086_60642# a_60945_60609# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X362 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X363 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X364 VDDD a_63621_58960# a_63571_58652# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X365 a_67027_69308# a_66049_69295# a_66825_69663# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X366 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X367 c1_45456_57458# m3_45124_57418# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X368 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X369 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X370 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X371 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X372 a_62593_58639# a_62409_59007# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X373 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X374 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X375 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X376 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X377 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X378 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X379 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X380 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X381 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X382 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X383 VSSD a_66666_49313# a_66865_49412# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X384 a_68479_59984# a_67881_60339# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X385 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X386 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X387 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X388 VDDD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X389 a_63457_56931# a_63273_56639# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X390 sar10b_0.clk_div_0.COUNT\[2\] a_66865_52076# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X391 VSSR sar10b_0.SWP[6] a_15533_113041# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X392 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X393 a_65966_58354# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X394 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X395 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X396 a_66762_50329# a_65778_49979# a_66464_50363# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X397 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X398 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X399 a_66183_56703# a_65857_56931# a_66062_57022# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X400 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X401 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X402 VSSD a_65643_48621# sar10b_0.SWN[5] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X403 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X404 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X405 a_67077_69616# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X406 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X407 c1_n1140_32818# m3_n1472_32778# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X408 VSSD sar10b_0.net16 a_62796_63063# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X409 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X410 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X411 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X412 VDDD a_61419_48621# th_dif_sw_0.CKB VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X413 a_65861_49313# a_65682_49313# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X414 VSSD a_68421_66952# a_68379_67056# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X415 a_62185_64695# a_61400_64952# a_61677_64842# VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X416 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X417 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X418 a_66375_69663# a_66049_69295# a_66254_69344# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X419 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X420 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_51345_60437# a_51861_60437# VDDA sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X421 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X422 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X423 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=10.44 ps=85.92 w=1.5 l=0.5
X424 VSSR sar10b_0.SWP[7] a_10731_113461# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X425 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X426 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X427 a_66386_49720# a_65861_49313# a_66216_49358# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X428 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X429 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X430 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X431 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X432 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X433 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X434 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X435 a_19457_110450# sar10b_0.SWP[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X436 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X437 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X438 a_67020_67059# sar10b_0.net46 a_66933_67059# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X439 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X440 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X441 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X442 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X443 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X444 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X445 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X446 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X447 a_53652_59132# tdc_0.phase_detector_0.INP VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X448 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X449 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X450 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X451 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X452 a_64761_51028# a_64188_51135# a_64428_50947# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.07875 ps=0.865 w=0.42 l=0.15
X453 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X454 a_67598_64016# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X455 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X456 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X457 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X458 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X459 VDDR sar10b_0.CF[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X460 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X461 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X462 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y sar10b_0.CF[7] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X463 a_63759_59064# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X464 VSSR sar10b_0.SWN[4] a_25137_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X465 a_24259_5788# sar10b_0.SWN[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X466 a_62796_63063# sar10b_0.net2 a_62709_63063# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X467 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X468 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X469 a_60747_61567# sar10b_0.net9 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X470 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X471 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X472 VDDD sar10b_0.net16 a_61677_52854# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X473 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X474 a_60789_53739# sar10b_0.net5 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X475 a_68379_67056# a_67209_66999# a_68169_66999# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X476 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X477 a_15533_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X478 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X479 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=13.92 ps=114.56 w=1.5 l=0.5
X480 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X481 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[8] a_7670_8700# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X482 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X483 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X484 a_24259_109594# sar10b_0.SWP[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X485 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X486 a_19457_5788# sar10b_0.SWN[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X487 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X488 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X489 VSSR sar10b_0.CF[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X490 VSSD a_60945_64605# a_60747_64605# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X491 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X492 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=10.44 ps=113.76 w=0.5 l=0.5
X493 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X494 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X495 VDDD a_68671_55988# sar10b_0.net20 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X496 VDDD a_61929_56639# a_62181_56768# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X497 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X498 VSSR sar10b_0.SWP[4] a_25137_112201# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X499 a_25137_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X500 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X501 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X502 a_12472_8700# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X503 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X504 a_61454_53360# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X505 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X506 VSSD sar10b_0.net3 a_66924_56403# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X507 a_40248_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X508 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X509 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X510 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X511 a_65996_50650# sar10b_0._01_ VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.08873 pd=0.895 as=0.2544 ps=2.2 w=0.42 l=0.15
X512 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X513 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X514 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X515 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X516 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X517 VDDD a_66464_50363# a_66419_50408# VDDD sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X518 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X519 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X520 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X521 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X522 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X523 a_19457_110450# sar10b_0.SWP[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X524 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X525 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X526 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X527 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X528 c1_10156_21618# m3_9824_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X529 c1_45456_82292# m3_45124_82252# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X530 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X531 a_55282_59893# tdc_0.phase_detector_0.pd_out_0.B VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.2352 ps=1.54 w=1.12 l=0.15
X532 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X533 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X534 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X535 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X536 a_67400_60020# a_66921_60339# a_67310_60020# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X537 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X538 VDDD a_66885_56768# a_66835_57058# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X539 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X540 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X541 a_10731_113461# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X542 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X543 a_61173_49986# a_60945_49953# a_61086_49986# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X544 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_109594# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X545 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X546 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X547 a_68421_68284# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X548 a_n4470_65264# th_dif_sw_0.CK VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.11655 ps=1.055 w=0.74 l=0.15
X549 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X550 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=27.84 ps=229.12 w=1.5 l=0.5
X551 a_66254_69344# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X552 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X553 VDDD EN a_60690_49683# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X554 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X555 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X556 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X557 a_66924_56403# sar10b_0.net40 a_66837_56403# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X558 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X559 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X560 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X561 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X562 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X563 c1_45456_97972# m3_45124_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X564 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X565 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X566 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_51345_60437# VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X567 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X568 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X569 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X570 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X571 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X572 a_24259_109594# sar10b_0.SWP[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X573 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X574 a_66419_50408# a_65778_49979# a_66312_50368# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X575 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X576 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X577 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=6.96 ps=75.84 w=0.5 l=0.5
X578 a_61358_58354# a_61153_58263# a_60693_57975# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X579 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X580 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X581 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X582 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X583 a_60945_49953# a_61395_49960# a_61347_49986# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X584 a_29061_5788# sar10b_0.SWN[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X585 a_5051_5788# sar10b_0.SWN[8] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X586 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X587 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X588 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=9.28 ps=101.12 w=0.5 l=0.5
X589 sar10b_0._06_ a_67055_68689# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1988 ps=1.505 w=1.12 l=0.15
X590 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X591 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X592 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=34.8 ps=286.39999 w=1.5 l=0.5
X593 a_20335_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X594 a_66464_50363# a_66312_50368# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X595 VSSD sar10b_0.net12 a_64809_65963# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X596 a_66795_71265# sar10b_0.net44 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X597 VSSR sar10b_0.SWN[6] a_15533_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X598 a_63339_48621# sar10b_0.net31 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X599 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X600 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X601 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X602 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X603 a_66666_49313# a_65861_49313# a_66368_49417# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X604 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X605 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X606 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X607 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X608 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X609 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X610 VSSD sar10b_0.net3 a_67797_65667# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X611 a_64814_65014# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X612 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X613 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X614 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=17.4 ps=143.2 w=1.5 l=0.5
X615 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X616 a_66210_50650# a_65586_50645# a_66103_50668# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.08873 ps=0.895 w=0.42 l=0.15
X617 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X618 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X619 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=8.12 ps=88.48 w=0.5 l=0.5
X620 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X621 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X622 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X623 VSSA th_dif_sw_0.th_sw_1.CK a_n8277_54565# VSSA sky130_fd_pr__nfet_01v8 ad=2.175 pd=15.58 as=2.175 ps=15.58 w=7.5 l=0.15
X624 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X625 sar10b_0._00_ a_65021_50292# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.33483 ps=1.765 w=1.12 l=0.15
X626 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X627 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X628 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X629 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X630 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X631 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X632 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X633 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X634 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X635 a_65871_59310# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X636 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X637 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X638 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X639 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=17.4 ps=143.2 w=1.5 l=0.5
X640 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X641 a_60945_52617# a_61400_52964# a_61349_53062# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X642 VSSR sar10b_0.SWP[9] a_1127_114301# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X643 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X644 VSSD a_61395_63280# a_61400_63620# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X645 a_61609_66266# a_61400_66284# a_60945_65937# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X646 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X647 VDDD a_61493_56924# a_61448_57022# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X648 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X649 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X650 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X651 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X652 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X653 VDDD a_66080_53027# a_66035_53072# VDDD sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X654 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X655 VDDD a_67733_64115# a_67688_64016# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X656 a_65333_66248# a_65198_66346# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X657 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X658 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X659 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X660 a_62131_51730# a_61153_51603# a_61929_51311# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X661 VSSD a_65119_59984# sar10b_0.net33 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X662 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X663 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X664 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X665 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X666 a_67797_65667# a_67733_65447# a_67719_65667# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X667 c1_n1140_72212# m3_n1472_72172# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X668 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X669 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X670 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X671 a_29061_5788# sar10b_0.SWN[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X672 VDDD sar10b_0._14_ a_67419_52937# VDDD sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.196 ps=1.47 w=1.12 l=0.15
X673 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X674 a_67310_61352# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X675 VDDD a_61395_61948# a_61400_62288# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X676 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X677 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X678 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X679 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X680 a_19457_5788# sar10b_0.SWN[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X681 VSSD sar10b_0.cyclic_flag_0.FINAL a_66921_60339# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X682 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X683 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X684 a_63950_60020# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X685 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X686 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X687 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X688 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X689 VDDD a_62181_58100# a_62131_58390# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X690 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X691 a_67372_52243# sar10b_0.clk_div_0.COUNT\[1\] VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.09625 pd=0.9 as=0.14887 ps=1.195 w=0.55 l=0.15
X692 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X693 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X694 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X695 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X696 a_63169_62635# a_62985_63003# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X697 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X698 VSSD a_64491_71265# sar10b_0.SWP[4] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X699 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X700 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X701 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X702 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X703 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X704 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X705 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X706 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X707 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X708 a_63804_67580# a_63663_67678# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.18405 pd=1.43 as=0.295 ps=2.59 w=1 l=0.15
X709 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X710 a_25137_112201# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X711 a_67688_64016# a_67209_64335# a_67598_64016# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X712 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X713 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X714 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X715 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[1] a_41284_8700# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X716 VSSA th_dif_sw_0.th_sw_1.CK a_n8277_54249# VSSA sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X717 a_67719_65667# a_67393_65299# a_67598_65348# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X718 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X719 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X720 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X721 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X722 VSSD a_60945_49953# a_60747_49953# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X723 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X724 a_66109_49318# sar10b_0._02_ VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X725 VSSR sar10b_0.CF[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X726 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X727 a_63918_50969# a_64188_51135# a_64146_51029# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.05565 ps=0.685 w=0.42 l=0.15
X728 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X729 a_69003_71265# sar10b_0.net46 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X730 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X731 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X732 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X733 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X734 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X735 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X736 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X737 VSSR sar10b_0.SWP[7] a_10731_113461# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X738 a_61347_64638# a_61086_64638# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X739 a_67445_60119# a_67310_60020# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X740 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X741 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X742 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X743 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X744 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X745 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X746 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X747 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X748 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X749 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X750 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X751 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X752 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X753 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X754 a_29061_108738# sar10b_0.SWP[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X755 a_67598_54692# a_67393_54643# a_66933_55071# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X756 VSSD a_66368_49417# a_66386_49720# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X757 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=20.88 ps=171.84 w=1.5 l=0.5
X758 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X759 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X760 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X761 a_25842_111636# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X762 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X763 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X764 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X765 a_24259_109594# sar10b_0.SWP[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X766 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X767 VSSD a_67077_57628# a_67035_57732# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X768 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X769 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X770 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X771 VSSD sar10b_0.clk_div_0.COUNT\[1\] a_67564_50907# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.33275 pd=2.31 as=0.17738 ps=1.195 w=0.55 l=0.15
X772 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X773 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X774 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X775 a_69003_71265# sar10b_0.net46 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X776 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=24.36 ps=200.48 w=1.5 l=0.5
X777 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X778 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X779 VSSR sar10b_0.SWN[3] a_29939_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X780 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X781 a_61589_53459# a_61454_53360# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X782 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X783 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X784 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X785 VSSD a_68671_55988# sar10b_0.net20 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X786 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X787 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_110450# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X788 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X789 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_108738# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X790 a_14655_5788# sar10b_0.SWN[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X791 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X792 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X793 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X794 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X795 a_62527_67630# a_61929_67295# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X796 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X797 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X798 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X799 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X800 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X801 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X802 a_61803_48621# sar10b_0.net28 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X803 VDDD a_67135_58306# sar10b_0.net36 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X804 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X805 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=5.8 ps=63.2 w=0.5 l=0.5
X806 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X807 VDDD sar10b_0.net16 a_62709_63063# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X808 a_67372_52243# a_67696_52265# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.09212 pd=0.885 as=0.11412 ps=0.965 w=0.55 l=0.15
X809 VSSD a_61677_52854# a_61609_52946# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X810 VSSD a_66378_52993# a_66577_52883# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X811 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X812 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X813 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X814 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X815 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X816 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X817 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X818 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X819 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X820 VDDD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X821 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X822 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X823 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X824 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X825 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X826 a_66389_69443# a_66254_69344# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X827 a_67055_68689# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.252 ps=2.28 w=0.84 l=0.15
X828 a_61644_57735# sar10b_0.net2 a_61557_57735# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X829 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X830 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X831 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X832 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X833 a_61609_62270# a_61395_61948# a_60945_61941# VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X834 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X835 a_61358_67678# a_61153_67587# a_60693_67299# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X836 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X837 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X838 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X839 VSSD a_66021_66092# a_65979_65970# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X840 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X841 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X842 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X843 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X844 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X845 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X846 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X847 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X848 a_62702_61352# a_62497_61303# a_62037_61731# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X849 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X850 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X851 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X852 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X853 a_63169_62635# a_62985_63003# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X854 a_10731_113461# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X855 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X856 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X857 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X858 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X859 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X860 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X861 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X862 a_66312_50368# a_65778_49979# a_66205_50408# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.15563 ps=1.215 w=0.42 l=0.15
X863 VDDA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X864 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X865 a_29061_108738# sar10b_0.SWP[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X866 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X867 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X868 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X869 a_62038_50362# a_61609_50282# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X870 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X871 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X872 a_1127_114301# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X873 VSSR sar10b_0.SWP[3] a_29939_111781# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X874 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X875 VDDD sar10b_0.net26 a_68946_65963# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X876 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X877 c1_29924_21618# m3_29592_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X878 VSSD sar10b_0.net16 a_61173_49986# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X879 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X880 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X881 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X882 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X883 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X884 a_68169_59007# a_67393_58639# a_67733_58787# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X885 a_63273_61671# a_62497_61303# a_62837_61451# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X886 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X887 VSSA th_dif_sw_0.CKB a_n4470_53722# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.11655 pd=1.055 as=0.1295 ps=1.09 w=0.74 l=0.15
X888 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X889 a_60693_57975# sar10b_0.net7 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X890 VDDD a_67445_61451# a_67400_61352# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X891 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X892 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X893 a_61677_64842# a_61400_64952# a_62007_64695# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X894 a_61086_49986# a_60945_49953# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X895 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X896 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X897 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X898 a_67135_58306# a_66537_57971# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X899 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X900 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X901 VDDD sar10b_0._12_ a_67439_50041# VDDD sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.147 ps=1.19 w=0.84 l=0.15
X902 a_61395_52624# sar10b_0.net4 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X903 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X904 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X905 a_62187_71265# sar10b_0.net40 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X906 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X907 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X908 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X909 a_68275_55988# a_67297_55975# a_68073_56343# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X910 a_65407_63634# a_64809_63299# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X911 a_62025_51015# a_61065_51015# a_61589_50795# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X912 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X913 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X914 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X915 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X916 VSSD sar10b_0.net16 a_60876_53739# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X917 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X918 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X919 sar10b_0.clk_div_0.COUNT\[0\] a_66865_49412# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X920 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X921 a_20335_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X922 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X923 VSSD a_62181_58100# a_62139_57978# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X924 VSSA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X925 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X926 VDDD a_63045_57628# a_62995_57320# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X927 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X928 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X929 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X930 VSSD a_67423_69308# sar10b_0.net47 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X931 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X932 a_62185_60699# sar10b_0.net8 a_62706_60639# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X933 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=27.84 ps=229.12 w=1.5 l=0.5
X934 a_60945_61941# a_61400_62288# a_61349_62386# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X935 tdc_0.OUTP tdc_0.OUTN VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X936 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X937 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X938 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X939 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X940 a_66344_57356# a_65865_57675# a_66254_57356# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X941 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X942 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X943 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X944 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X945 a_9853_112162# sar10b_0.SWP[7] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X946 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X947 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X948 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X949 a_65013_64695# a_64949_64916# a_64935_64695# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X950 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X951 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X952 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X953 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X954 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X955 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X956 VDDD sar10b_0.clknet_0_CLK a_66153_48647# VDDD sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X957 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X958 VDDD sar10b_0.net5 a_60969_51311# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X959 VSSA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X960 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X961 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X962 c1_n1140_49618# m3_n1472_49578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X963 a_64335_63060# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X964 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X965 a_60747_68227# sar10b_0.net13 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X966 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X967 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X968 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X969 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X970 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X971 VDDD a_68421_58960# a_68371_58652# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X972 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X973 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X974 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X975 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X976 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X977 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X978 a_62181_51440# a_61929_51311# a_62319_51318# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X979 VDDD sar10b_0.clk_div_0.COUNT\[3\] a_67843_52961# VDDD sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X980 a_67393_58639# a_67209_59007# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X981 a_29061_108738# sar10b_0.SWP[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X982 a_62497_61303# a_62313_61671# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X983 a_60876_53739# sar10b_0.net5 a_60789_53739# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X984 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X985 VDDD a_63369_59007# a_63621_58960# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X986 VDDD CLK a_65577_51311# VDDD sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X987 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X988 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X989 a_61929_57971# a_60969_57971# a_61493_58256# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X990 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X991 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X992 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X993 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X994 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X995 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X996 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X997 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X998 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X999 a_67564_50907# sar10b_0.clk_div_0.COUNT\[0\] VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.17738 pd=1.195 as=0.12607 ps=1.1 w=0.55 l=0.15
X1000 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X1001 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1002 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1003 VDDD sar10b_0.net1 a_62185_50043# VDDD sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X1004 VDDD a_60747_58903# sar10b_0.CF[2] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X1005 a_62706_60639# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1006 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1007 a_65733_59432# a_65481_59303# a_65871_59310# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X1008 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1009 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1010 a_67231_56974# a_66633_56639# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1011 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1012 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1013 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X1014 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1015 c1_45456_27218# m3_45124_27178# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1016 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1017 VDDD a_64492_67433# a_64445_67714# VDDD sky130_fd_pr__pfet_01v8 ad=0.0735 pd=0.77 as=0.0567 ps=0.69 w=0.42 l=0.15
X1018 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1019 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1020 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1021 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X1022 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1023 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1024 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1025 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 a_5051_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1026 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1027 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1028 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1029 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1030 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1031 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1032 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1033 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1034 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1035 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1036 a_67733_66779# a_67598_66680# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X1037 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1038 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1039 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1040 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1041 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1042 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1043 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1044 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1045 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1046 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1047 sar10b_0.net12 a_60747_64605# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X1048 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1049 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1050 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1051 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1052 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1053 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1054 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1055 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1056 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X1057 VDDD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1058 a_n4470_53722# th_dif_sw_0.CKB VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.11655 ps=1.055 w=0.74 l=0.15
X1059 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1060 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1061 a_19457_110450# sar10b_0.SWP[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1062 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1063 VDDR sar10b_0.CF[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1064 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1065 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1066 VDDD sar10b_0.clknet_1_1__leaf_CLK a_65586_50645# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1067 VSSR sar10b_0.SWP[6] a_15533_113041# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1068 a_68463_56400# sar10b_0.net3 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X1069 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1070 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y sar10b_0.CF[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1071 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1072 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1073 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1074 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1075 a_67733_54791# a_67598_54692# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X1076 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1077 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1078 VDDD a_61035_48621# sar10b_0.SWN[1] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X1079 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1080 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1081 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1082 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1083 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1084 VDDD a_66537_57971# a_66789_58100# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1085 c1_n1140_51858# m3_n1472_51818# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1086 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1087 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1088 a_68559_59064# sar10b_0.net3 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X1089 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1090 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1091 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1092 a_68276_50645# sar10b_0.clk_div_0.COUNT\[1\] VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1848 ps=1.45 w=1.12 l=0.15
X1093 a_63967_58652# a_63369_59007# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1094 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1095 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1096 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1097 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1098 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1099 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1100 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1101 VDDD a_63945_63003# a_64197_62956# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1102 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1103 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1104 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1105 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1106 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1107 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1108 VSSR sar10b_0.SWP[7] a_10731_113461# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1109 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1110 VSSA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1111 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1112 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1113 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1114 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1115 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1116 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1117 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1118 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1119 a_62131_57058# a_61153_56931# a_61929_56639# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X1120 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1121 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1122 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1123 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1124 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1125 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1126 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1127 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1128 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1129 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1130 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1131 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1132 a_65761_58263# a_65577_57971# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1133 sar10b_0.clknet_0_CLK a_65577_51311# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1134 VDDD sar10b_0.net10 a_63561_60339# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1135 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1136 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1137 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A a_30644_111636# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1138 c1_39808_97972# m3_39476_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1139 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1140 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1141 VDDD a_66197_56924# a_66152_57022# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X1142 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1143 a_61349_53062# a_61086_52650# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X1144 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=6.96 ps=57.28 w=1.5 l=0.5
X1145 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1146 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1147 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1148 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1149 a_61677_52854# a_61400_52964# a_62007_52707# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X1150 a_52504_60961# tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_52417_60961# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.1824 ps=1.85 w=0.64 l=0.15
X1151 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1152 VDDD sar10b_0.net16 a_64149_64635# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X1153 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1154 VSSR sar10b_0.SWN[4] a_25137_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1155 c1_n1140_74452# m3_n1472_74412# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1156 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1157 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1158 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1159 VSSD a_61677_62178# a_61609_62270# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X1160 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1161 VSSD sar10b_0.net19 a_68946_49747# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X1162 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y sar10b_0.CF[9] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1163 a_62181_67424# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X1164 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1165 VDDD a_64780_52239# sar10b_0._11_ VDDD sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.308 ps=2.79 w=1.12 l=0.15
X1166 a_30644_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1167 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1168 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1169 a_62126_56024# a_61921_55975# a_61461_56403# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X1170 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1171 VSSR sar10b_0.SWP[4] a_25137_112201# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1172 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1173 VSSD a_68133_61624# a_68091_61728# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X1174 a_25137_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1175 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1176 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1177 a_62281_52347# a_61496_52091# a_61773_52237# VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X1178 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1179 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1180 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1181 VSSD sar10b_0.net9 a_62409_59007# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1182 a_n4470_65264# th_dif_sw_0.CK VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1183 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1184 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1185 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1186 VDDD a_68479_59984# sar10b_0.net21 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1187 a_66152_57022# a_65673_56639# a_66062_57022# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X1188 a_66080_53027# a_65928_53032# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X1189 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1190 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1191 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y a_1832_8706# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1192 DATA[6] a_68946_61735# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X1193 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1194 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1195 VSSD sar10b_0.net16 a_63862_67359# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.35328 pd=1.84 as=0.0504 ps=0.66 w=0.42 l=0.15
X1196 a_61544_50696# a_61065_51015# a_61454_50696# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X1197 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1198 a_67215_69720# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X1199 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1200 VSSD a_66885_56768# a_66843_56646# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X1201 VDDD sar10b_0.net16 a_63285_60399# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X1202 VSSD sar10b_0.net16 a_61653_51015# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X1203 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1204 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1205 VSSD a_66559_68962# sar10b_0.net46 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X1206 a_60693_67299# sar10b_0.net13 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X1207 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1208 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1209 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1210 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1211 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X1212 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1213 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1214 VSSD a_60690_70625# sar10b_0.net2 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X1215 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X1216 a_66062_57022# a_65673_56639# a_65397_56643# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X1217 a_68169_63003# a_67393_62635# a_67733_62783# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X1218 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1219 a_61395_61948# sar10b_0.net4 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X1220 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1221 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1222 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1223 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1224 a_66927_57978# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X1225 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1226 c1_45456_67732# m3_45124_67692# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1227 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1228 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1229 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1230 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1231 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1232 a_66254_69344# a_65865_69663# a_65589_69723# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X1233 VDDA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1234 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1235 a_62185_66027# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X1236 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1237 c1_45456_44018# m3_45124_43978# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1238 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1239 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1240 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1241 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1242 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1243 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 a_5051_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1244 sar10b_0.net9 a_60747_60609# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X1245 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1246 VSSD sar10b_0._07_ a_64050_51311# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1247 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X1248 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1249 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1250 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1251 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1252 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1253 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1254 a_62933_58787# a_62798_58688# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X1255 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1256 VSSR sar10b_0.SWN[4] a_25137_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1257 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1258 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1259 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1260 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1261 a_63862_67359# a_63804_67580# a_63784_67359# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1262 c1_n1140_89012# m3_n1472_88972# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1263 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1264 a_68083_59984# a_67105_59971# a_67881_60339# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X1265 a_65236_49657# sar10b_0._07_ VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.15535 ps=1.17 w=0.64 l=0.15
X1266 a_61653_51015# a_61589_50795# a_61575_51015# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1267 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1268 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1269 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1270 a_10731_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1271 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1272 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1273 a_64491_48621# sar10b_0.net32 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X1274 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1275 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1276 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1277 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1278 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1279 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1280 VDDD a_68421_68284# a_68371_67976# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X1281 VSSD a_68767_65312# sar10b_0.net25 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X1282 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1283 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1284 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1285 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1286 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1287 a_67020_68391# sar10b_0.net47 a_66933_68391# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1288 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1289 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1290 a_20335_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1291 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1292 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1293 VDDD sar10b_0.clknet_0_CLK a_66153_48647# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1294 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1295 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1296 VSSR sar10b_0.SWN[6] a_15533_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1297 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1298 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X1299 a_61929_67295# a_60969_67295# a_61493_67580# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X1300 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1301 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1302 a_67393_62635# a_67209_63003# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X1303 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1304 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1305 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1306 VSSD a_66577_52883# a_66535_52693# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05565 ps=0.685 w=0.42 l=0.15
X1307 a_68421_66952# a_68169_66999# a_68559_67056# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X1308 VSSD a_64773_60292# a_64731_60396# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X1309 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1310 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1311 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X1312 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1313 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1314 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1315 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1316 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X1317 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1318 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1319 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1320 sar10b_0.clknet_0_CLK a_65577_51311# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X1321 a_61395_52624# sar10b_0.net4 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1322 VDDD a_60747_62899# sar10b_0.CF[5] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X1323 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1324 a_66823_49697# a_65682_49313# a_66666_49313# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X1325 a_63784_67359# a_63457_67583# a_63663_67678# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X1326 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1327 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1328 a_68169_63003# a_67209_63003# a_67733_62783# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X1329 a_68371_66644# a_67393_66631# a_68169_66999# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X1330 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1331 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1332 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1333 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1334 a_67744_51002# sar10b_0.clk_div_0.COUNT\[0\] sar10b_0._12_ VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1554 ps=1.16 w=0.74 l=0.15
X1335 a_61575_51015# a_61249_50647# a_61454_50696# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X1336 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1337 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1338 sar10b_0.net1 a_60690_54641# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1339 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1340 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1341 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1342 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1343 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1344 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X1345 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1346 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1347 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1348 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_108738# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1349 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1350 a_62281_52347# a_61491_52222# a_61773_52237# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X1351 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1352 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1353 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1354 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1355 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1356 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1357 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1358 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1359 a_62793_57675# a_62017_57307# a_62357_57455# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X1360 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1361 VDDD a_61929_57971# a_62181_58100# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1362 VSSR sar10b_0.SWP[9] a_1127_114301# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1363 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1364 VDDD sar10b_0.clk_div_0.COUNT\[2\] a_68178_51635# VDDD sky130_fd_pr__pfet_01v8 ad=0.36323 pd=1.84 as=0.126 ps=1.14 w=0.84 l=0.15
X1365 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1366 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1367 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1368 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1369 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1370 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1371 VSSD sar10b_0.clknet_0_CLK a_65355_53949# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.063 pd=0.72 as=0.0588 ps=0.7 w=0.42 l=0.15
X1372 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X1373 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1374 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1375 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1376 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1377 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1378 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1379 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1380 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1381 c1_n1140_91252# m3_n1472_91212# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1382 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1383 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1384 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1385 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1386 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1387 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1388 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1389 a_67733_64115# a_67598_64016# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X1390 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1391 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1392 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1393 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1394 a_68559_68388# sar10b_0.net3 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X1395 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1396 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1397 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1398 a_41284_111642# sar10b_0.CF[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1399 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1400 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1401 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1402 a_68559_63060# sar10b_0.net3 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X1403 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1404 sar10b_0.net3 a_60690_49683# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.435 as=0.1876 ps=1.455 w=1.12 l=0.15
X1405 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1406 a_n4470_65264# th_dif_sw_0.CK VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1407 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1408 VDDD a_66785_50875# sar10b_0.net16 VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1409 a_62527_56974# a_61929_56639# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X1410 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1411 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1412 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[3] a_31680_8700# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1413 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1414 c1_n1140_36178# m3_n1472_36138# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1415 VSSD sar10b_0._06_ a_67890_69727# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X1416 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1417 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1418 VSSA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1419 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1420 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1421 VSSR sar10b_0.CF[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1422 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1423 a_25137_112201# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1424 VDDA th_dif_sw_0.CK a_n4470_65264# VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1425 VDDD sar10b_0.net6 a_62281_52347# VDDD sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X1426 VDDD sar10b_0._08_ a_68943_51605# VDDD sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.1512 ps=1.39 w=1.12 l=0.15
X1427 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1428 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1429 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1430 VDDD a_60690_49683# sar10b_0.net3 VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1764 ps=1.435 w=1.12 l=0.15
X1431 a_62017_57307# a_61833_57675# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X1432 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1433 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1434 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1435 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1436 a_61677_52854# a_61395_52624# a_62038_53026# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X1437 a_n4470_65264# th_dif_sw_0.CK VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1438 a_68325_56296# a_68073_56343# a_68463_56400# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X1439 a_61349_62386# a_61086_61974# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X1440 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1441 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1442 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1443 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1444 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1445 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1446 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1447 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1448 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1449 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1450 c1_45456_84532# m3_45124_84492# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1451 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1452 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1453 VSSR sar10b_0.SWP[7] a_10731_113461# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1454 a_61358_51694# a_61153_51603# a_60693_51315# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X1455 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1456 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1457 a_24259_5788# sar10b_0.SWN[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1458 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1459 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1460 a_26878_8700# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X1461 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1462 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_108738# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1463 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1464 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1465 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1466 a_62025_53679# a_61249_53311# a_61589_53459# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X1467 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1468 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1469 a_65996_50650# sar10b_0._01_ VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.35502 ps=2.6 w=0.42 l=0.15
X1470 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1471 a_60747_58903# sar10b_0.net7 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X1472 VDDD a_65637_64760# a_65587_65050# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X1473 a_61269_52404# a_61041_52340# a_61182_52404# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X1474 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1475 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1476 VSSD a_62277_50968# a_62235_51072# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X1477 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1478 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1479 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1480 c1_45456_29458# m3_45124_29418# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1481 VSSD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X1482 VDDD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1483 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1484 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1485 c1_272_21618# m3_n60_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1486 VSSD sar10b_0.net16 a_61557_58035# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X1487 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1488 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1489 sar10b_0.SWP[9] a_68946_71059# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X1490 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1491 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1492 VDDD a_62697_56343# a_62949_56296# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1493 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1494 VSSR sar10b_0.SWN[3] a_29939_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1495 a_66255_50749# a_66103_50668# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2226 pd=1.37 as=0.23985 ps=1.735 w=0.84 l=0.15
X1496 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1497 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1498 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1499 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1500 VSSD sar10b_0.net16 a_64437_63363# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X1501 VDDD a_64491_71265# sar10b_0.SWP[4] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X1502 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1503 VDDD a_60945_63273# a_60747_63273# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X1504 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1505 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1506 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1507 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1508 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1509 a_67419_52937# a_67372_52833# sar10b_0._16_ VDDD sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3864 ps=2.93 w=1.12 l=0.15
X1510 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1511 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1512 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1513 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1514 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y a_21040_8706# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X1515 a_67035_69720# a_65865_69663# a_66825_69663# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X1516 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1517 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1518 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1519 VDDR sar10b_0.CF[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1520 DATA[0] a_68562_48647# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X1521 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1522 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1523 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1524 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1525 sar10b_0._14_ a_68178_51635# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.36323 ps=1.84 w=1.12 l=0.15
X1526 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1527 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1528 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1529 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1530 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1531 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1532 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1533 a_67393_67963# a_67209_68331# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X1534 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X1535 a_66747_57978# a_65577_57971# a_66537_57971# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X1536 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1537 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1538 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1539 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1540 VSSD sar10b_0.net12 a_65865_57675# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1541 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1542 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1543 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1544 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1545 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1546 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X1547 VDDD sar10b_0.net6 a_61737_56343# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1548 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1549 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1550 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1551 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1552 a_61557_58035# a_61493_58256# a_61479_58035# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1553 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1554 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1555 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1556 VDDD a_61395_63280# a_61400_63620# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1557 VSSD sar10b_0.cyclic_flag_0.FINAL a_66921_61671# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1558 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_108738# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1559 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1560 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X1561 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1562 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1563 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1564 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1565 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1566 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1567 a_67077_69616# a_66825_69663# a_67215_69720# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X1568 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1569 a_67598_65348# a_67209_65667# a_66933_65727# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X1570 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X1571 VSSD a_64888_67630# sar10b_0.cyclic_flag_0.FINAL VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2072 pd=2.04 as=0.1036 ps=1.02 w=0.74 l=0.15
X1572 a_63273_61671# a_62313_61671# a_62837_61451# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X1573 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1574 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1575 VDDD a_61677_63510# a_61609_63602# VDDD sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X1576 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1577 a_65861_51977# a_65682_51977# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1578 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1579 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1580 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1581 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1582 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1583 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1584 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1585 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1586 a_65577_51311# CLK VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X1587 a_66789_58100# a_66537_57971# a_66927_57978# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X1588 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1589 VDDD a_66079_59638# sar10b_0.net34 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1590 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1591 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X1592 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X1593 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1594 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1595 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1596 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1597 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1598 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1599 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1600 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1601 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1602 a_1127_114301# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1603 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1604 c1_45456_31698# m3_45124_31658# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1605 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1606 VDDD a_62793_57675# a_63045_57628# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1607 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1608 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1609 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1610 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1611 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X1612 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1613 VDDD sar10b_0.cyclic_flag_0.FINAL a_67113_56343# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1614 a_61929_56639# a_61153_56931# a_61493_56924# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X1615 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1616 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1617 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1618 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1619 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1620 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1621 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1622 a_61479_58035# a_61153_58263# a_61358_58354# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X1623 a_61929_51311# a_61153_51603# a_61493_51596# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X1624 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1625 a_66389_57455# a_66254_57356# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X1626 VDDD a_62357_57455# a_62312_57356# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X1627 c1_n1140_76692# m3_n1472_76652# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1628 a_10731_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1629 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1630 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1631 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1632 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1633 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1634 VSSD sar10b_0.net3 a_67020_67059# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X1635 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1636 a_64543_62648# a_63945_63003# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1637 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1638 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1639 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1640 a_61347_65970# a_61086_65970# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X1641 a_67445_61451# a_67310_61352# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X1642 VDDD sar10b_0.net16 a_61677_63510# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X1643 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X1644 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1645 VDDD a_68169_59007# a_68421_58960# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1646 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1647 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1648 a_20335_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1649 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1650 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1651 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1652 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1653 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1654 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1655 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1656 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1657 a_64339_51661# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2562 pd=2.29 as=0.2814 ps=2.35 w=0.84 l=0.15
X1658 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1659 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1660 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1661 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1662 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1663 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1664 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1665 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1666 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1667 a_66205_50408# sar10b_0._03_ VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
X1668 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1669 VDDA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1670 a_66645_60399# sar10b_0.net41 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X1671 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 a_9853_112162# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1672 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1673 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1674 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1675 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1676 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1677 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1678 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1679 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1680 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1681 a_64583_51628# a_64339_51661# a_64454_51311# VDDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X1682 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1683 a_63753_67678# a_63273_67295# a_63663_67678# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X1684 sar10b_0.clknet_0_CLK a_65577_51311# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X1685 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1686 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1687 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1688 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1689 a_62312_57356# a_61833_57675# a_62222_57356# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X1690 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1691 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1692 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1693 a_61358_58354# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X1694 a_64521_60339# a_63745_59971# a_64085_60119# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X1695 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1696 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1697 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1698 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1699 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1700 a_n9133_57045# th_dif_sw_0.th_sw_1.CKB VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.15
X1701 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1702 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1703 a_10731_113461# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1704 VDDD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X1705 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1706 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1707 c1_45456_69972# m3_45124_69932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1708 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1709 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1710 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1711 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1712 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1713 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1714 c1_45456_46258# m3_45124_46218# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1715 c1_27100_97972# m3_26768_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1716 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1717 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1718 VSSD sar10b_0.net9 a_62985_63003# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1719 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1720 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1721 VSSD a_65637_64760# a_65595_64638# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X1722 a_66739_58390# a_65761_58263# a_66537_57971# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X1723 a_66825_57675# a_65865_57675# a_66389_57455# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X1724 a_68271_61728# sar10b_0.net3 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X1725 a_66933_67059# sar10b_0.net46 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X1726 VDDD a_62025_53679# a_62277_53632# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1727 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1728 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1729 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1730 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1731 VDDD sar10b_0.net16 a_61557_57735# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X1732 a_65021_50292# sar10b_0._09_ a_64818_49979# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.0896 ps=0.92 w=0.64 l=0.15
X1733 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1734 a_64454_51311# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.08663 pd=0.865 as=0.1155 ps=0.97 w=0.55 l=0.15
X1735 VDDA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1736 a_68767_58652# a_68169_59007# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1737 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1738 VDDD sar10b_0._00_ a_64761_51028# VDDD sky130_fd_pr__pfet_01v8 ad=0.2972 pd=2.41 as=0.09835 ps=1.005 w=0.42 l=0.15
X1739 VDDD sar10b_0.net16 a_61086_60642# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X1740 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1741 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1742 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X1743 a_62181_51440# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X1744 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X1745 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_109594# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1746 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1747 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1748 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1749 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1750 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1751 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1752 c1_n1140_21618# m3_n1472_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1753 a_67439_50041# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.252 ps=2.28 w=0.84 l=0.15
X1754 VSSD a_61395_52624# a_61400_52964# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X1755 a_66837_56403# sar10b_0.net40 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X1756 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1757 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1758 a_61548_56403# sar10b_0.net2 a_61461_56403# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1759 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1760 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1761 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 a_9853_112162# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1762 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1763 VDDD a_61131_70891# sar10b_0.SWP[0] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X1764 VDDA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1765 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1766 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1767 VSSD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X1768 VSSD a_65577_51311# sar10b_0.clknet_0_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1769 VDDD a_61419_71265# th_dif_sw_0.CK VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X1770 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1771 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1772 VSSR sar10b_0.SWP[6] a_15533_113041# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1773 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1774 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1775 a_60747_68227# sar10b_0.net13 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X1776 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1777 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1778 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1779 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1780 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1781 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1782 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1783 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1784 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1785 a_65595_64638# a_64425_64631# a_65385_64631# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X1786 VDDD a_66825_69663# a_67077_69616# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1787 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1788 a_66021_66092# a_65769_65963# a_66159_65970# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X1789 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1790 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1791 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1792 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=13.92 ps=114.56 w=1.5 l=0.5
X1793 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1794 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1795 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1796 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1797 c1_32748_21618# m3_32416_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1798 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1799 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1800 VDDD sar10b_0.net19 a_68946_49747# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X1801 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1802 a_60693_51315# sar10b_0.net1 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X1803 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1804 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1805 VSSD sar10b_0.net16 a_61557_67359# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X1806 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1807 VSSD a_68421_65620# a_68379_65724# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X1808 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1809 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1810 a_62187_48621# sar10b_0.net30 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X1811 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1812 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1813 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1814 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1815 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1816 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1817 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1818 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1819 VSSD a_60945_63273# a_60747_63273# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X1820 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1821 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1822 VDDD a_66865_49412# a_66773_49313# VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.09975 ps=0.895 w=0.42 l=0.15
X1823 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1824 VDDD sar10b_0.net11 a_64425_64631# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X1825 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1826 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1827 c1_35572_97972# m3_35240_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1828 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1829 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1830 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1831 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1832 a_67020_65727# sar10b_0.net45 a_66933_65727# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1833 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1834 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1835 a_66835_57058# a_65857_56931# a_66633_56639# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X1836 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1837 a_62185_62031# sar10b_0.net9 a_62706_61971# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X1838 VSSD sar10b_0.cyclic_flag_0.FINAL a_67209_59007# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1839 VSSD sar10b_0.net8 a_62313_61671# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X1840 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1841 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1842 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1843 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1844 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X1845 a_63945_63003# a_63169_62635# a_63509_62783# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X1846 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1847 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X1848 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X1849 c1_n1140_93492# m3_n1472_93452# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1850 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1851 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_109594# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1852 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1853 a_9853_5788# sar10b_0.SWN[7] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1854 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1855 VDDD a_66368_49417# a_66323_49318# VDDD sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X1856 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1857 VSSD sar10b_0.net3 a_67509_60339# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X1858 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1859 VDDR sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X1860 VDDD sar10b_0.net16 a_60789_53739# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X1861 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1862 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1863 a_62181_58100# a_61929_57971# a_62319_57978# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X1864 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X1865 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X1866 VSSD a_66785_50875# sar10b_0.net16 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1867 a_61557_67359# a_61493_67580# a_61479_67359# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1868 a_64911_60396# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X1869 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1870 a_68379_65724# a_67209_65667# a_68169_65667# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X1871 VSSD a_60690_53975# sar10b_0.net4 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X1872 a_66885_56768# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X1873 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1874 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1875 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1876 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1877 VDDD a_67423_69308# sar10b_0.net47 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X1878 VSSR sar10b_0.SWP[4] a_25137_112201# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1879 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1880 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y sar10b_0.CF[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1881 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X1882 a_25137_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1883 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1884 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1885 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1886 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1887 VSSD a_62623_50660# sar10b_0.net30 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X1888 a_67598_54692# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X1889 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1890 c1_45456_71092# m3_45124_71052# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1891 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1892 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X1893 a_67372_52243# a_67798_52206# a_67747_51991# VDDD sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X1894 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X1895 a_67231_56974# a_66633_56639# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X1896 a_62706_61971# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X1897 a_29061_5788# sar10b_0.SWN[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1898 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1899 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1900 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1901 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1902 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1903 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X1904 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X1905 DATA[8] a_68946_65963# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X1906 a_n8277_66083# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS VINP VSSA sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X1907 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1908 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1909 a_62837_61451# a_62702_61352# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X1910 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X1911 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1912 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1913 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1914 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1915 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1916 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1917 a_66323_49318# a_65682_49313# a_66216_49358# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X1918 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1919 a_67509_60339# a_67445_60119# a_67431_60339# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X1920 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1921 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1922 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1923 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1924 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1925 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1926 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1927 a_61479_67359# a_61153_67587# a_61358_67678# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X1928 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1929 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X1930 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1931 c1_45456_86772# m3_45124_86732# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1932 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1933 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1934 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1935 a_64809_63299# a_63849_63299# a_64373_63584# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X1936 VDDD a_64373_63584# a_64328_63682# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X1937 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1938 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1939 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1940 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1941 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1942 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1943 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1944 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X1945 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1946 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1947 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1948 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1949 VDDD a_68169_68331# a_68421_68284# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X1950 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X1951 a_60690_49683# EN VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1952 a_63945_63003# a_62985_63003# a_63509_62783# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X1953 a_62185_63363# a_61395_63280# a_61677_63510# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X1954 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1955 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1956 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1957 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X1958 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1959 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1960 VDDD a_66577_52883# a_66485_53077# VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.09975 ps=0.895 w=0.42 l=0.15
X1961 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X1962 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1963 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X1964 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1965 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X1966 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X1967 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1968 a_65587_65050# a_64609_64923# a_65385_64631# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X1969 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X1970 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X1971 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1972 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1973 VDDD sar10b_0.clknet_1_0__leaf_CLK a_65778_49979# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X1974 a_61448_58354# a_60969_57971# a_61358_58354# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X1975 a_65979_65970# a_64809_65963# a_65769_65963# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X1976 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1977 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X1978 a_10731_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1979 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1980 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1981 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1982 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1983 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1984 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1985 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X1986 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X1987 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X1988 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1989 a_61358_67678# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X1990 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1991 a_62798_58688# a_62593_58639# a_62133_59067# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X1992 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1993 a_29061_5788# sar10b_0.SWN[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1994 a_64328_63682# a_63849_63299# a_64238_63682# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X1995 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X1996 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X1997 a_66537_57971# a_65761_58263# a_66101_58256# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X1998 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X1999 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2000 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2001 a_62131_58390# a_61153_58263# a_61929_57971# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X2002 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2003 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2004 VSSD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2005 a_24259_109594# sar10b_0.SWP[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2006 a_19457_5788# sar10b_0.SWN[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2007 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2008 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2009 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2010 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2011 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2012 VSSD a_67084_53565# sar10b_0._17_ VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.2109 ps=2.05 w=0.74 l=0.15
X2013 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2014 a_65481_59303# a_64521_59303# a_65045_59588# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X2015 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2016 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2017 VDDD sar10b_0.net18 a_68562_48647# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X2018 a_66368_49417# a_66216_49358# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X2019 a_68325_56296# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X2020 a_60747_56239# sar10b_0.net5 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X2021 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2022 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2023 VDDD sar10b_0.cyclic_flag_0.FINAL a_67209_66999# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2024 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2025 c1_10156_97972# m3_9824_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2026 VSSD a_66666_51977# a_66865_52076# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X2027 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2028 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2029 a_62007_64695# a_61609_64934# a_61929_64695# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2030 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2031 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2032 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2033 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2034 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X2035 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2036 VDDR sar10b_0.CF[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2037 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2038 a_n8277_66083# th_dif_sw_0.th_sw_1.CK VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X2039 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2040 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2041 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2042 sar10b_0.net3 a_60690_49683# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2043 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2044 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2045 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2046 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X2047 a_68767_67976# a_68169_68331# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2048 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2049 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2050 a_68479_59984# a_67881_60339# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X2051 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2052 a_68767_62648# a_68169_63003# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2053 a_63391_57320# a_62793_57675# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2054 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2055 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2056 a_66386_52384# a_65861_51977# a_66216_52022# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X2057 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2058 VSSR sar10b_0.SWP[3] a_29939_111781# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2059 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2060 VSSD a_61395_61948# a_61400_62288# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X2061 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2062 a_62798_58688# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X2063 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2064 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2065 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2066 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2067 a_9853_5788# sar10b_0.SWN[7] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2068 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2069 a_65761_58263# a_65577_57971# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X2070 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X2071 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2072 a_61929_64695# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2073 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2074 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2075 a_66633_56639# a_65673_56639# a_66197_56924# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X2076 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2077 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2078 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2079 a_61395_61948# sar10b_0.net4 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2080 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2081 VDDD sar10b_0.net3 a_66933_67059# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X2082 a_55121_59650# tdc_0.phase_detector_0.pd_out_0.A VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.17738 pd=1.195 as=0.33275 ps=2.31 w=0.55 l=0.15
X2083 VDDD a_60945_52617# a_60747_52617# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X2084 a_66633_56639# a_65857_56931# a_66197_56924# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X2085 VDDD a_61395_60616# a_61400_60956# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2086 a_68133_61624# a_67881_61671# a_68271_61728# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X2087 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2088 a_24259_109594# sar10b_0.SWP[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2089 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2090 a_19457_5788# sar10b_0.SWN[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2091 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2092 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2093 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2094 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2095 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2096 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2097 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2098 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2099 a_65188_51977# a_64924_52385# a_64780_52239# VDDD sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.3 as=0.275 ps=2.55 w=1 l=0.15
X2100 a_68767_66644# a_68169_66999# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X2101 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X2102 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2103 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2104 VDDD a_67423_57320# sar10b_0.net35 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X2105 VDDD a_61677_60846# a_61609_60938# VDDD sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X2106 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2107 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2108 VDDD a_67733_54791# a_67688_54692# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X2109 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2110 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2111 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2112 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2113 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2114 a_64050_51311# sar10b_0.net3 sar10b_0._08_ VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2115 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2116 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2117 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2118 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2119 VSSR sar10b_0.SWP[6] a_15533_113041# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2120 a_25137_112201# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2121 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2122 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2123 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2124 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2125 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2126 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2127 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2128 VSSD sar10b_0.cyclic_flag_0.FINAL a_67209_63003# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2129 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2130 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2131 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2132 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2133 c1_8744_21618# m3_8412_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2134 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2135 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2136 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2137 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2138 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2139 VSSD a_65577_51311# sar10b_0.clknet_0_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X2140 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2141 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2142 a_63663_67678# a_63273_67295# a_62997_67299# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X2143 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2144 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2145 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[7] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X2146 a_61454_50696# a_61065_51015# a_60789_51075# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X2147 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2148 a_67688_54692# a_67209_55011# a_67598_54692# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X2149 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2150 a_62623_53324# a_62025_53679# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2151 a_65857_56931# a_65673_56639# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X2152 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2153 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2154 VSSD sar10b_0.net3 a_67797_55011# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2155 a_62038_65014# a_61609_64934# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X2156 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2157 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2158 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2159 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2160 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2161 a_61773_52237# a_61496_52091# a_62103_52347# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2162 a_64731_60396# a_63561_60339# a_64521_60339# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2163 VDDD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X2164 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2165 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2166 c1_45456_48498# m3_45124_48458# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2167 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2168 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=24.36 ps=200.48 w=1.5 l=0.5
X2169 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2170 VSSR sar10b_0.SWN[8] a_5929_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2171 sar10b_0.net4 a_60690_53975# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2172 a_62181_56768# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X2173 a_68169_64335# a_67209_64335# a_67733_64115# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X2174 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2175 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2176 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2177 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2178 VDDD a_68767_65312# sar10b_0.net25 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X2179 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2180 w_n9655_63119# a_n9133_63315# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS w_n9655_63119# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X2181 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2182 a_68235_48621# sar10b_0.net35 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X2183 VDDD a_62837_61451# a_62792_61352# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X2184 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2185 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2186 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2187 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2188 a_64773_60292# a_64521_60339# a_64911_60396# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X2189 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2190 a_65385_64631# a_64609_64923# a_64949_64916# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X2191 c1_n1140_23858# m3_n1472_23818# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2192 VSSD a_62181_67424# a_62139_67302# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X2193 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2194 a_67797_55011# a_67733_54791# a_67719_55011# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2195 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2196 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2197 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2198 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2199 a_62697_56343# a_61921_55975# a_62261_56123# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X2200 a_62103_52347# a_61705_51992# a_62025_52347# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2201 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2202 a_62007_52707# a_61609_52946# a_61929_52707# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2203 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2204 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2205 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2206 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2207 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2208 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2209 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2210 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_110450# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2211 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X2212 VSSD EN a_60690_49683# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.2109 ps=2.05 w=0.74 l=0.15
X2213 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2214 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2215 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2216 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2217 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2218 VSSR sar10b_0.SWP[7] a_10731_113461# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2219 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2220 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2221 a_5929_113881# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2222 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2223 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2224 VSSD sar10b_0.net7 a_61833_57675# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2225 a_61448_67678# a_60969_67295# a_61358_67678# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X2226 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2227 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2228 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2229 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2230 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X2231 VSSD a_61419_48621# th_dif_sw_0.CKB VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X2232 a_62792_61352# a_62313_61671# a_62702_61352# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X2233 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2234 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2235 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2236 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2237 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2238 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X2239 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2240 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2241 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2242 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2243 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2244 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2245 a_67843_52961# sar10b_0._14_ a_67372_52833# VDDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X2246 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2247 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2248 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2249 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=1.16 ps=12.64 w=0.5 l=0.5
X2250 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2251 a_67719_55011# a_67393_54643# a_67598_54692# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2252 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2253 VSSD EN a_60690_49683# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2254 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2255 VDDD sar10b_0.net4 a_60969_57971# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2256 a_61929_52707# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X2257 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2258 VSSR sar10b_0.SWN[4] a_25137_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2259 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2260 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2261 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2262 VDDD sar10b_0.net16 a_60693_57975# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X2263 a_64609_64923# a_64425_64631# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X2264 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2265 VDDD sar10b_0.net16 a_61086_49986# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X2266 a_64445_67714# a_63457_67583# a_64238_67295# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.22695 ps=1.83 w=0.42 l=0.15
X2267 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2268 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2269 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2270 a_60747_60235# sar10b_0.net8 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X2271 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2272 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2273 a_10731_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2274 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2275 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2276 a_61921_55975# a_61737_56343# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X2277 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2278 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2279 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2280 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2281 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2282 VSSD a_65061_63428# a_65019_63306# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X2283 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2284 a_62997_67299# sar10b_0.net14 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X2285 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2286 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2287 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2288 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2289 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2290 VSSD a_63339_71265# sar10b_0.SWP[3] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X2291 a_20335_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2292 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2293 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2294 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2295 c1_n1140_38418# m3_n1472_38378# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2296 VDDD a_62623_50660# sar10b_0.net30 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X2297 a_62697_56343# a_61737_56343# a_62261_56123# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X2298 a_65397_56643# sar10b_0.net1 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X2299 a_68133_60292# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X2300 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2301 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2302 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_110450# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2303 VSSD sar10b_0.net16 a_62997_59007# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2304 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2305 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2306 VDDA tdc_0.phase_detector_0.pd_out_0.B tdc_0.OUTP VDDA sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2307 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2308 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2309 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2310 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2311 a_30644_111636# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2312 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2313 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2314 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2315 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2316 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2317 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2318 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2319 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2320 a_67747_51991# a_67696_52265# a_67651_51991# VDDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X2321 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2322 VSSD sar10b_0.net16 a_65388_57975# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2323 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2324 c1_20040_21618# m3_19708_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2325 a_61153_51603# a_60969_51311# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2326 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2327 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2328 VSSD sar10b_0.net16 a_61557_51375# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2329 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2330 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2331 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2332 VDDA CLK a_52417_59293# VDDA sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.147 ps=1.19 w=0.84 l=0.15
X2333 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2334 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2335 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2336 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2337 a_66378_52993# a_65394_52643# a_66080_53027# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X2338 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2339 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2340 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2341 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2342 c1_29924_97972# m3_29592_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2343 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2344 a_61443_52404# a_61182_52404# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X2345 a_9853_112162# sar10b_0.SWP[7] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2346 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2347 sar10b_0._06_ a_67055_68689# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X2348 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2349 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2350 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2351 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X2352 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_109594# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2353 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2354 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2355 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2356 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2357 a_61929_56639# a_60969_56639# a_61493_56924# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X2358 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2359 a_68421_66952# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X2360 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2361 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2362 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2363 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2364 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2365 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2366 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2367 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2368 VSSD a_66368_52081# a_66386_52384# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X2369 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2370 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2371 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2372 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2373 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2374 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2375 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2376 a_65388_57975# sar10b_0.net1 a_65301_57975# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X2377 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2378 VSSD a_66367_66298# sar10b_0.net45 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2379 a_61358_57022# a_61153_56931# a_60693_56643# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X2380 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2381 a_61557_51375# a_61493_51596# a_61479_51375# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2382 VDDD a_69003_48621# sar10b_0.SWN[8] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X2383 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X2384 sar10b_0._04_ sar10b_0._14_ VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2385 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2386 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2387 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2388 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2389 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2390 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X2391 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2392 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2393 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2394 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2395 c1_n1140_40658# m3_n1472_40618# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2396 a_20335_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2397 a_61358_58354# a_60969_57971# a_60693_57975# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X2398 VDDD a_61035_71265# sar10b_0.SWP[1] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X2399 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X2400 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2401 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2402 a_64888_67630# a_64238_67295# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2072 ps=2.04 w=0.74 l=0.15
X2403 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2404 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2405 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2406 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2407 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2408 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2409 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2410 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2411 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2412 a_65765_50645# a_65586_50645# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2413 VSSR sar10b_0.SWP[6] a_15533_113041# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2414 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2415 a_63339_48621# sar10b_0.net31 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2416 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2417 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2418 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2419 VDDR sar10b_0.CF[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2420 VSSD sar10b_0.net3 a_67797_64335# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2421 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A a_31680_111642# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2422 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2423 VSSD a_63525_61624# a_63483_61728# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X2424 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2425 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2426 a_66773_49313# a_65861_49313# a_66666_49313# VDDD sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X2427 a_61929_57971# a_61153_58263# a_61493_58256# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X2428 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2429 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2430 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2431 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2432 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2433 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2434 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2435 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2436 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2437 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2438 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2439 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2440 a_46086_8700# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X2441 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2442 sar10b_0._15_ sar10b_0.clk_div_0.COUNT\[2\] a_68276_50645# VDDD sky130_fd_pr__pfet_01v8 ad=0.308 pd=2.79 as=0.168 ps=1.42 w=1.12 l=0.15
X2443 a_9853_112162# sar10b_0.SWP[7] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2444 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2445 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[9] a_2868_8700# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2446 a_19457_110450# sar10b_0.SWP[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2447 VSSD sar10b_0.net3 a_67020_68391# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2448 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2449 a_61479_51375# a_61153_51603# a_61358_51694# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2450 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2451 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2452 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2453 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y a_35446_8706# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2454 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2455 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2456 VDDD a_62261_56123# a_62216_56024# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X2457 a_64910_59686# a_64705_59595# a_64245_59307# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X2458 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2459 VSSD CLK a_65577_51311# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X2460 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2461 VSSR sar10b_0.SWP[5] a_20335_112621# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2462 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2463 c1_n1140_63252# m3_n1472_63212# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2464 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2465 a_63374_62684# a_63169_62635# a_62709_63063# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X2466 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2467 a_61609_64934# a_61400_64952# a_60945_64605# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X2468 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2469 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X2470 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2471 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y sar10b_0.CF[8] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X2472 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2473 VDDD a_65577_51311# sar10b_0.clknet_0_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2474 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2475 a_63745_59971# a_63561_60339# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2476 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2477 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2478 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2479 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2480 c1_45456_33938# m3_45124_33898# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2481 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2482 a_66737_51029# a_65586_50645# a_66593_50645# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.06615 pd=0.735 as=0.1076 ps=0.985 w=0.42 l=0.15
X2483 VDDR sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2484 tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.pd_out_0.A a_53652_61050# VSSA sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X2485 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2486 a_67797_64335# a_67733_64115# a_67719_64335# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2487 VSSR sar10b_0.SWN[8] a_5929_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2488 a_63483_61728# a_62313_61671# a_63273_61671# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2489 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2490 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2491 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2492 a_67310_60020# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X2493 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2494 c1_n1140_78932# m3_n1472_78892# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2495 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2496 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2497 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2498 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2499 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 a_5051_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2500 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2501 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X2502 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2503 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2504 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2505 a_67084_53565# sar10b_0._10_ a_67252_53653# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1376 ps=1.14 w=0.64 l=0.15
X2506 VSSD a_66785_50875# a_66737_51029# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.06615 ps=0.735 w=0.42 l=0.15
X2507 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2508 a_61358_51694# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X2509 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2510 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2511 a_68083_61316# a_67105_61303# a_67881_61671# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X2512 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2513 c1_n1140_55218# m3_n1472_55178# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2514 VSSD sar10b_0.net16 a_66261_56703# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2515 a_29061_5788# sar10b_0.SWN[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2516 a_62216_56024# a_61737_56343# a_62126_56024# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X2517 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2518 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2519 VSSR sar10b_0.SWP[4] a_25137_112201# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2520 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2521 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2522 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2523 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2524 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A a_6634_111636# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2525 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2526 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2527 VSSD a_64780_52239# sar10b_0._11_ VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.11312 pd=1.065 as=0.1961 ps=2.01 w=0.74 l=0.15
X2528 a_61182_52404# a_61041_52340# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X2529 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2530 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2531 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2532 sar10b_0.net3 a_60690_49683# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2533 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2534 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2535 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2536 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2537 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2538 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2539 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2540 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2541 VDDD a_64188_51135# a_64199_50761# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2542 a_19457_110450# sar10b_0.SWP[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2543 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2544 a_67719_64335# a_67393_63967# a_67598_64016# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2545 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X2546 a_66933_68391# sar10b_0.net47 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X2547 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2548 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2549 tdc_0.phase_detector_0.INP a_52417_60961# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X2550 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2551 VDDD sar10b_0.net4 a_60969_67295# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2552 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2553 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2554 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2555 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2556 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2557 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2558 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2559 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X2560 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2561 VDDD sar10b_0.net16 a_60693_67299# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X2562 VSSD sar10b_0.net16 a_64236_64635# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2563 a_61677_63510# a_61395_63280# a_62038_63682# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X2564 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2565 a_5929_113881# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2566 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2567 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2568 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2569 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2570 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2571 VDDD sar10b_0.net16 a_61677_60846# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X2572 a_61347_63306# a_61086_63306# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X2573 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2574 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2575 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2576 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2577 a_67598_58688# a_67393_58639# a_66933_59067# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X2578 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2579 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2580 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2581 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2582 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_111306# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2583 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2584 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2585 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2586 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2587 VDDD sar10b_0.net12 a_62185_66027# VDDD sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X2588 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X2589 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2590 VDDD a_60747_69559# sar10b_0.CF[9] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X2591 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2592 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2593 a_24259_109594# sar10b_0.SWP[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2594 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X2595 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2596 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2597 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2598 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2599 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2600 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X2601 a_67142_68689# sar10b_0.net16 a_67055_68689# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.1824 ps=1.85 w=0.64 l=0.15
X2602 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2603 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2604 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2605 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X2606 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2607 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2608 sar10b_0.net7 a_60843_52216# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2609 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2610 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2611 a_29061_5788# sar10b_0.SWN[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2612 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2613 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2614 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2615 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2616 VSSD a_60747_65563# sar10b_0.CF[7] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X2617 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2618 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X2619 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2620 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2621 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2622 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2623 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A a_16238_111636# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2624 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2625 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2626 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2627 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2628 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2629 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2630 a_66153_48647# sar10b_0.clknet_0_CLK VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2631 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2632 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2633 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2634 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2635 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2636 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2637 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2638 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2639 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2640 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2641 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2642 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2643 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2644 a_61173_52650# a_60945_52617# a_61086_52650# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X2645 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2646 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2647 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2648 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X2649 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2650 a_68421_65620# a_68169_65667# a_68559_65724# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X2651 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2652 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2653 VSSD sar10b_0.net16 a_66453_57675# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2654 a_68943_51605# sar10b_0._14_ a_68841_51605# VDDD sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.2016 ps=1.48 w=1.12 l=0.15
X2655 DATA[1] a_68946_49747# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X2656 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2657 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2658 a_61609_66266# a_61395_65944# a_60945_65937# VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X2659 c1_24276_21618# m3_23944_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2660 VSSD sar10b_0.net3 a_67509_61671# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2661 VDDD sar10b_0.clk_div_0.COUNT\[0\] a_67611_50645# VDDD sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.196 ps=1.47 w=1.12 l=0.15
X2662 VDDD a_60690_54641# sar10b_0.net1 VDDD sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2663 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2664 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2665 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2666 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2667 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2668 a_66593_50645# a_65586_50645# a_66255_50749# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2226 ps=1.37 w=0.84 l=0.15
X2669 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2670 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2671 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2672 c1_n1140_80052# m3_n1472_80012# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2673 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2674 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2675 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2676 sar10b_0.net15 a_67890_69727# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X2677 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2678 VDDD a_68325_56296# a_68275_55988# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X2679 c1_45456_50738# m3_45124_50698# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2680 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2681 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2682 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2683 sar10b_0.SWN[9] a_68562_49747# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2684 a_60945_52617# a_61395_52624# a_61347_52650# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X2685 a_61358_67678# a_60969_67295# a_60693_67299# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X2686 VSSR sar10b_0.SWP[3] a_29939_111781# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2687 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X2688 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2689 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2690 a_20335_112621# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2691 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2692 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2693 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2694 sar10b_0.clk_div_0.COUNT\[3\] a_66577_52883# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X2695 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X2696 VSSD sar10b_0.net21 a_68946_53975# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X2697 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2698 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2699 c1_n1140_95732# m3_n1472_95692# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2700 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2701 a_66453_57675# a_66389_57455# a_66375_57675# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2702 VDDD a_67445_60119# a_67400_60020# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X2703 VSSD sar10b_0.clknet_1_0__leaf_CLK a_65778_49979# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X2704 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2705 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2706 a_61677_63510# a_61400_63620# a_62007_63363# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X2707 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2708 a_61609_50282# a_61400_50300# a_60945_49953# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X2709 a_67431_60339# a_67105_59971# a_67310_60020# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2710 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2711 a_66666_51977# a_65861_51977# a_66368_52081# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X2712 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2713 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X2714 a_67509_61671# a_67445_61451# a_67431_61671# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2715 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2716 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2717 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2718 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2719 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2720 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2721 a_67371_49579# sar10b_0.net34 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X2722 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2723 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2724 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X2725 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2726 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2727 a_66789_58100# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X2728 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2729 sar10b_0.net16 a_66785_50875# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2730 VSSD a_62181_56768# a_62139_56646# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X2731 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2732 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2733 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2734 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2735 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2736 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2737 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2738 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2739 a_63918_50969# a_64199_50761# a_64154_50645# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.09975 ps=0.895 w=0.42 l=0.15
X2740 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2741 c1_45456_73332# m3_45124_73292# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2742 a_60945_60609# a_61400_60956# a_61349_61054# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X2743 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2744 VSSR sar10b_0.SWP[6] a_15533_113041# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2745 a_25137_112201# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2746 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[5] a_22076_8700# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X2747 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2748 a_63509_62783# a_63374_62684# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X2749 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2750 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2751 VSSA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2752 a_29061_5788# sar10b_0.SWN[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2753 VSSD a_68421_54964# a_68379_55068# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X2754 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2755 a_62185_52707# a_61400_52964# a_61677_52854# VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X2756 a_66375_57675# a_66049_57307# a_66254_57356# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2757 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2758 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2759 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2760 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2761 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2762 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2763 VSSD a_68767_54656# sar10b_0.net18 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2764 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2765 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2766 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2767 a_61448_51694# a_60969_51311# a_61358_51694# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X2768 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2769 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2770 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2771 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2772 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2773 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2774 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2775 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2776 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2777 a_64907_50292# sar10b_0.net17 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.21 pd=1.42 as=0.295 ps=2.59 w=1 l=0.15
X2778 a_64149_64635# sar10b_0.net2 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X2779 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2780 VDDD a_60690_49683# sar10b_0.net3 VDDD sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.196 ps=1.47 w=1.12 l=0.15
X2781 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X2782 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X2783 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2784 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2785 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2786 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2787 sar10b_0.net1 a_60690_54641# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X2788 a_60780_51315# sar10b_0.net1 a_60693_51315# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X2789 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2790 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2791 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2792 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2793 VDDD a_60747_57571# sar10b_0.CF[1] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X2794 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2795 VDDD a_66255_50749# a_66210_50650# VDDD sky130_fd_pr__pfet_01v8 ad=0.23985 pd=1.735 as=0.0504 ps=0.66 w=0.42 l=0.15
X2796 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2797 a_14655_111306# sar10b_0.SWP[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2798 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2799 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2800 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2801 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2802 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X2803 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2804 VSSR sar10b_0.SWN[8] a_5929_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2805 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2806 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2807 a_68379_55068# a_67209_55011# a_68169_55011# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2808 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2809 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2810 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2811 VSSD sar10b_0.net16 a_61557_56703# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X2812 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2813 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2814 a_67733_65447# a_67598_65348# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X2815 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2816 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2817 VSSA tdc_0.phase_detector_0.pd_out_0.B a_55121_59650# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.12607 pd=1.1 as=0.17738 ps=1.195 w=0.55 l=0.15
X2818 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2819 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2820 VSSD a_65577_51311# sar10b_0.clknet_0_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X2821 VSSD sar10b_0.net13 a_65577_57971# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2822 VSSD a_60945_52617# a_60747_52617# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X2823 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2824 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2825 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X2826 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2827 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2828 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2829 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2830 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2831 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2832 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X2833 a_64238_67295# a_63457_67583# a_63804_67580# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.12025 ps=1.065 w=0.74 l=0.15
X2834 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2835 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2836 VSSR sar10b_0.SWP[4] a_25137_112201# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2837 c1_n1140_42898# m3_n1472_42858# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2838 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2839 a_51861_59345# th_dif_sw_0.VCN VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X2840 a_62319_51318# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X2841 a_67733_58787# a_67598_58688# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X2842 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2843 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2844 a_67598_62684# a_67393_62635# a_66933_63063# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X2845 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2846 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2847 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2848 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2849 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X2850 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2851 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2852 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2853 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2854 a_67423_57320# a_66825_57675# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X2855 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2856 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2857 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2858 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2859 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2860 a_61395_63280# sar10b_0.net4 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2861 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2862 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2863 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2864 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2865 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2866 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2867 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2868 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2869 VDDD sar10b_0.net3 a_66933_68391# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X2870 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2871 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2872 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2873 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2874 VSSD a_61035_48621# sar10b_0.SWN[1] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X2875 a_61557_56703# a_61493_56924# a_61479_56703# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X2876 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2877 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2878 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X2879 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2880 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2881 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2882 a_62134_52028# a_61705_51992# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X2883 a_5929_113881# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2884 a_66255_50749# a_66103_50668# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.099 pd=0.985 as=0.19715 ps=1.365 w=0.55 l=0.15
X2885 a_61461_56403# sar10b_0.net2 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X2886 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2887 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2888 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2889 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2890 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2891 VDDD sar10b_0.net20 a_68946_52411# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X2892 a_66101_58256# a_65966_58354# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X2893 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2894 VDDA th_dif_sw_0.th_sw_1.CKB a_n9133_63315# VDDA sky130_fd_pr__pfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.15
X2895 VSSA CLK a_52504_60961# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1376 ps=1.14 w=0.64 l=0.15
X2896 a_66254_57356# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X2897 VDDD sar10b_0.cyclic_flag_0.FINAL a_66921_60339# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2898 c1_272_97972# m3_n60_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2899 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2900 c1_n1140_65492# m3_n1472_65452# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2901 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X2902 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2903 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2904 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X2905 VSSA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2906 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2907 DATA[5] a_68946_59303# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X2908 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2909 VDDD a_66865_52076# a_66773_51977# VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.09975 ps=0.895 w=0.42 l=0.15
X2910 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2911 VDDR sar10b_0.CF[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2912 a_68091_60396# a_66921_60339# a_67881_60339# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2913 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X2914 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X2915 VSSR sar10b_0.SWN[4] a_25137_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2916 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2917 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X2918 a_64448_67302# a_63273_67295# a_64238_67295# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X2919 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2920 a_67297_55975# a_67113_56343# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X2921 VSSD sar10b_0.net14 a_65673_56639# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X2922 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2923 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2924 VDDD sar10b_0._07_ a_64667_51628# VDDD sky130_fd_pr__pfet_01v8 ad=0.2382 pd=1.555 as=0.135 ps=1.27 w=1 l=0.15
X2925 a_61173_61974# a_60945_61941# a_61086_61974# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X2926 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2927 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X2928 VSSD a_61677_60846# a_61609_60938# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X2929 a_10731_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2930 a_61479_56703# a_61153_56931# a_61358_57022# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X2931 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2932 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2933 VSSD a_63967_58652# sar10b_0.net32 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X2934 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2935 VDDD sar10b_0.clk_div_0.COUNT\[1\] a_68178_51635# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.24 as=0.2478 ps=2.27 w=0.84 l=0.15
X2936 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X2937 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2938 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X2939 VSSD sar10b_0.net3 a_67020_65727# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X2940 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X2941 VDDD tdc_0.RDY a_60690_53975# VDDD sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3304 ps=2.83 w=1.12 l=0.15
X2942 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2943 a_25137_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2944 a_15533_113041# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2945 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2946 c1_n1140_57458# m3_n1472_57418# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2947 c1_45456_90132# m3_45124_90092# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2948 a_65637_64760# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X2949 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X2950 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X2951 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2952 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2953 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2954 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2955 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2956 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2957 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2958 VDDD sar10b_0.net4 a_61065_53679# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X2959 a_65390_69010# a_65185_68919# a_64725_68631# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X2960 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2961 c1_22864_21618# m3_22532_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2962 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X2963 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2964 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2965 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2966 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2967 a_60945_61941# a_61395_61948# a_61347_61974# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X2968 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X2969 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X2970 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X2971 VDDD sar10b_0.net3 a_66645_60399# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X2972 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2973 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2974 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2975 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X2976 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2977 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2978 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2979 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 a_9853_112162# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X2980 a_61086_65970# a_60945_65937# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X2981 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2982 a_62181_58100# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X2983 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2984 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X2985 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2986 a_67502_56024# a_67297_55975# a_66837_56403# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X2987 VSSD sar10b_0.net16 a_61173_52650# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X2988 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2989 a_66197_56924# a_66062_57022# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X2990 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2991 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2992 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2993 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2994 c1_45456_35058# m3_45124_35018# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2995 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X2996 a_61395_60616# sar10b_0.net4 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X2997 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2998 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X2999 VDDD a_68133_60292# a_68083_59984# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X3000 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3001 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3002 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3003 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3004 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3005 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3006 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3007 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3008 a_62185_64695# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X3009 a_68073_56343# a_67297_55975# a_67637_56123# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X3010 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3011 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3012 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3013 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3014 a_63369_59007# a_62409_59007# a_62933_58787# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X3015 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3016 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3017 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3018 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3019 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3020 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3021 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3022 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3023 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3024 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3025 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3026 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3027 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3028 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3029 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3030 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3031 a_10731_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3032 VSSA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3033 a_67598_54692# a_67209_55011# a_66933_55071# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X3034 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3035 VDDD a_62527_51646# sar10b_0.net28 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X3036 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3037 VSSR sar10b_0.SWN[3] a_29939_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3038 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3039 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3040 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3041 VSSD a_60690_49683# sar10b_0.net3 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.10545 ps=1.025 w=0.74 l=0.15
X3042 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3043 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3044 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X3045 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3046 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3047 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3048 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3049 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X3050 a_62181_67424# a_61929_67295# a_62319_67302# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X3051 VSSD sar10b_0.net11 a_64425_64631# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X3052 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3053 VDDD a_68421_66952# a_68371_66644# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X3054 VSSD a_68767_63980# sar10b_0.net23 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3055 VDDD sar10b_0.net3 a_66837_56403# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X3056 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3057 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3058 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3059 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3060 VSSD sar10b_0.net6 a_61737_56343# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X3061 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3062 a_67526_50041# sar10b_0.net3 a_67439_50041# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.1824 ps=1.85 w=0.64 l=0.15
X3063 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3064 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3065 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3066 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3067 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3068 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3069 a_25137_112201# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3070 a_36482_8700# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X3071 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3072 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3073 a_62187_71265# sar10b_0.net40 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3074 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3075 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3076 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3077 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3078 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X3079 a_68331_52243# sar10b_0._13_ VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3080 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3081 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3082 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3083 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3084 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3085 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3086 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y a_25842_8706# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3087 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3088 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3089 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3090 VDDD a_60747_61567# sar10b_0.CF[4] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3091 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3092 a_67297_55975# a_67113_56343# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3093 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3094 a_62623_50660# a_62025_51015# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X3095 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3096 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3097 a_68371_65312# a_67393_65299# a_68169_65667# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X3098 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3099 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 a_9853_112162# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3100 VDDD sar10b_0.net16 a_60693_51315# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X3101 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3102 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3103 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3104 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3105 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3106 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3107 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3108 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3109 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X3110 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3111 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3112 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3113 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3114 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3115 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3116 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3117 a_64609_64923# a_64425_64631# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3118 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3119 c1_n1140_82292# m3_n1472_82252# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3120 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3121 VSSD a_60945_61941# a_60747_61941# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3122 VSSR sar10b_0.SWP[5] a_20335_112621# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3123 a_66062_57022# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X3124 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3125 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3126 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3127 a_64949_64916# a_64814_65014# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X3128 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3129 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3130 a_52417_59293# tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.252 ps=2.28 w=0.84 l=0.15
X3131 a_61454_50696# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X3132 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3133 a_66109_49318# sar10b_0._02_ VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
X3134 c1_45456_52978# m3_45124_52938# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3135 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3136 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3137 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3138 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X3139 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3140 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3141 a_n4470_65264# th_dif_sw_0.CK VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3142 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3143 VSSD sar10b_0.net17 a_64818_49979# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.1824 ps=1.85 w=0.64 l=0.15
X3144 a_65061_63428# a_64809_63299# a_65199_63306# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X3145 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3146 a_61929_67295# a_61153_67587# a_61493_67580# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X3147 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3148 a_67733_62783# a_67598_62684# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X3149 c1_n1140_97972# m3_n1472_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3150 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3151 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3152 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3153 a_68559_67056# sar10b_0.net3 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X3154 a_62139_51318# a_60969_51311# a_61929_51311# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X3155 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3156 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3157 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3158 a_11436_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X3159 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3160 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3161 a_64888_67630# a_64238_67295# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1638 ps=1.275 w=0.84 l=0.15
X3162 sar10b_0.net15 a_67890_69727# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3163 VSSD sar10b_0.net15 a_68562_71291# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X3164 a_63663_67678# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.1393 ps=1.17 w=0.42 l=0.15
X3165 VSSR sar10b_0.SWP[4] a_25137_112201# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3166 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3167 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3168 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3169 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3170 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3171 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3172 VSSD sar10b_0._15_ sar10b_0._04_ VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X3173 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3174 c1_32748_97972# m3_32416_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3175 sar10b_0._13_ a_67439_50041# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X3176 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3177 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3178 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3179 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3180 c1_45456_75572# m3_45124_75532# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3181 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 a_9853_112162# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3182 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3183 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3184 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3185 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3186 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3187 VSSD a_63810_50901# sar10b_0.net17 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.2109 ps=2.05 w=0.74 l=0.15
X3188 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3189 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3190 a_19457_5788# sar10b_0.SWN[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3191 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X3192 c1_18628_21618# m3_18296_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3193 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3194 a_61349_61054# a_61086_60642# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X3195 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3196 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X3197 DATA[7] a_68946_63299# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3198 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3199 a_61609_50282# a_61395_49960# a_60945_49953# VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X3200 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3201 VDDD a_68767_54656# sar10b_0.net18 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X3202 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3203 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3204 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3205 VDDA CLK a_51345_58977# VDDA sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X3206 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3207 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3208 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3209 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3210 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3211 a_67445_61451# a_67310_61352# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X3212 tdc_0.phase_detector_0.INN a_52417_59293# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1988 ps=1.505 w=1.12 l=0.15
X3213 c1_44044_21618# m3_43712_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3214 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3215 VSSD sar10b_0.clk_div_0.COUNT\[3\] a_67798_52206# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1155 pd=0.97 as=0.15675 ps=1.67 w=0.55 l=0.15
X3216 VDDD a_62933_58787# a_62888_58688# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X3217 a_64085_60119# a_63950_60020# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X3218 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X3219 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3220 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3221 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3222 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3223 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3224 VSSD sar10b_0.net20 a_68946_52411# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X3225 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3226 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3227 VDDD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3228 VDDD sar10b_0.net21 a_68946_53975# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3229 a_61358_51694# a_60969_51311# a_60693_51315# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X3230 a_62025_52347# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X3231 a_68479_61316# a_67881_61671# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X3232 a_64809_63299# a_64033_63591# a_64373_63584# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X3233 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3234 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3235 VDDD EN a_60690_49683# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3236 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3237 th_dif_sw_0.VCN th_dif_sw_0.th_sw_0.th_sw_main_0.VGS VINN VSSA sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=0.15
X3238 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3239 VDDD sar10b_0.cyclic_flag_0.FINAL a_67209_65667# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X3240 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3241 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3242 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3243 a_67105_59971# a_66921_60339# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3244 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3245 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3246 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3247 VSSD sar10b_0.net16 a_63372_60399# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3248 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3249 a_66593_50645# a_65765_50645# a_66255_50749# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1076 pd=0.985 as=0.099 ps=0.985 w=0.55 l=0.15
X3250 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3251 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3252 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3253 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3254 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3255 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3256 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3257 a_65957_50273# a_65778_49979# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3258 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X3259 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3260 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3261 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3262 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3263 a_9853_5788# sar10b_0.SWN[7] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3264 VSSD a_60690_53975# sar10b_0.net4 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0672 ps=0.74 w=0.42 l=0.15
X3265 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3266 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3267 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3268 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3269 VSSD sar10b_0.net16 a_61173_61974# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X3270 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3271 VDDD a_60945_61941# a_60747_61941# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X3272 VDDD sar10b_0.net15 a_68562_71291# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3273 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3274 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3275 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3276 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3277 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3278 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3279 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3280 a_62888_58688# a_62409_59007# a_62798_58688# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X3281 a_1127_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3282 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3283 VSSD a_67423_57320# sar10b_0.net35 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3284 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3285 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3286 a_66885_56768# a_66633_56639# a_67023_56646# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X3287 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3288 a_60945_49953# a_61400_50300# a_61349_50398# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X3289 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3290 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3291 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3292 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3293 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3294 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3295 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3296 w_n9655_56533# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS VDDA w_n9655_56533# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X3297 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3298 VDDD a_68073_56343# a_68325_56296# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X3299 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3300 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3301 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3302 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3303 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3304 a_67393_66631# a_67209_66999# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3305 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3306 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X3307 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X3308 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3309 a_63372_60399# sar10b_0.net1 a_63285_60399# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3310 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3311 a_60747_56239# sar10b_0.net5 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3312 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3313 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3314 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3315 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3316 a_65019_63306# a_63849_63299# a_64809_63299# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X3317 VDDD a_60690_49683# sar10b_0.net3 VDDD sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3318 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y sar10b_0.CF[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3319 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3320 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3321 a_66153_48647# sar10b_0.clknet_0_CLK VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.063 ps=0.72 w=0.42 l=0.15
X3322 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3323 a_67598_64016# a_67209_64335# a_66933_64395# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X3324 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3325 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3326 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3327 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3328 VDDD a_61677_62178# a_61609_62270# VDDD sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X3329 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3330 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3331 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3332 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3333 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3334 a_62997_59007# a_62933_58787# a_62919_59007# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X3335 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3336 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3337 VSSR sar10b_0.SWP[3] a_29939_111781# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3338 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3339 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X3340 VDDD a_66762_50329# a_66961_50219# VDDD sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X3341 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3342 a_20335_112621# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3343 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3344 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3345 a_64238_67295# a_63273_67295# a_63804_67580# VDDD sky130_fd_pr__pfet_01v8 ad=0.22695 pd=1.83 as=0.18405 ps=1.43 w=1 l=0.15
X3346 sar10b_0._02_ sar10b_0._08_ VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3347 a_n9133_57045# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS a_n8277_54249# VSSA sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X3348 sar10b_0.clknet_0_CLK a_65577_51311# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3349 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X3350 a_9853_5788# sar10b_0.SWN[7] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3351 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3352 a_67733_54791# a_67598_54692# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X3353 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3354 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3355 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3356 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3357 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3358 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3359 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3360 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3361 a_64154_50645# a_63810_50901# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1239 ps=1.43 w=0.42 l=0.15
X3362 a_61395_60616# sar10b_0.net4 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3363 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3364 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3365 VSSR sar10b_0.SWN[3] a_29939_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3366 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3367 VDDD a_63967_58652# sar10b_0.net32 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X3368 sar10b_0.net5 a_60747_52617# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X3369 a_62421_57675# a_62357_57455# a_62343_57675# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X3370 VDDD sar10b_0.net16 a_61677_62178# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X3371 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3372 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3373 sar10b_0.net3 a_60690_49683# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.10545 pd=1.025 as=0.1554 ps=1.16 w=0.74 l=0.15
X3374 VDDD sar10b_0.net16 a_65188_51977# VDDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.15 ps=1.3 w=1 l=0.15
X3375 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3376 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3377 a_66823_52361# a_65682_51977# a_66666_51977# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X3378 a_64667_51628# sar10b_0.net16 a_64583_51628# VDDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3379 VDDD a_63804_67580# a_63753_67678# VDDD sky130_fd_pr__pfet_01v8 ad=0.1393 pd=1.17 as=0.0567 ps=0.69 w=0.42 l=0.15
X3380 a_20335_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3381 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[7] a_12472_8700# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3382 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3383 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3384 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3385 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3386 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3387 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3388 VSSR sar10b_0.CF[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3389 a_62919_59007# a_62593_58639# a_62798_58688# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X3390 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3391 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3392 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3393 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3394 c1_45456_92372# m3_45124_92332# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3395 a_29061_5788# sar10b_0.SWN[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3396 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3397 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3398 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3399 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3400 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3401 sar10b_0._01_ a_64338_52411# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3402 a_25137_112201# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3403 a_63457_67583# a_63273_67295# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1554 ps=1.16 w=0.74 l=0.15
X3404 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3405 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3406 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3407 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3408 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3409 a_61803_48621# sar10b_0.net28 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3410 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3411 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3412 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3413 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3414 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3415 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3416 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3417 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3418 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3419 VDDA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VDDA sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3420 VSSD sar10b_0.net25 a_68946_63299# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X3421 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3422 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3423 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3424 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3425 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3426 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3427 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3428 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3429 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3430 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3431 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3432 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3433 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3434 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3435 a_61358_57022# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X3436 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3437 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X3438 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3439 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3440 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3441 c1_45456_37298# m3_45124_37258# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3442 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3443 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3444 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3445 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X3446 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3447 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3448 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3449 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3450 a_67611_50645# a_67564_50907# sar10b_0._12_ VDDD sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.3864 ps=2.93 w=1.12 l=0.15
X3451 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3452 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3453 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3454 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3455 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3456 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X3457 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3458 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3459 VDDD a_60690_53975# sar10b_0.net4 VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3460 VINN th_dif_sw_0.th_sw_1.CK VINN VSSA sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=18.56 ps=130.32001 w=20 l=0.15
X3461 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3462 VDDA th_dif_sw_0.CK a_n4470_65264# VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3463 a_61086_63306# a_60945_63273# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X3464 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X3465 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3466 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3467 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3468 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3469 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3470 a_61677_60846# a_61395_60616# a_62038_61018# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X3471 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3472 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3473 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3474 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3475 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3476 VDDD a_68767_63980# sar10b_0.net23 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X3477 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3478 a_67310_60020# a_66921_60339# a_66645_60399# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X3479 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3480 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3481 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3482 VSSR sar10b_0.SWP[4] a_25137_112201# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3483 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3484 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3485 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3486 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3487 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3488 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3489 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3490 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3491 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3492 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3493 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3494 VSSR sar10b_0.SWP[6] a_15533_113041# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3495 VSSD a_62187_48621# sar10b_0.SWN[2] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X3496 VSSD sar10b_0.net24 a_68946_61735# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X3497 a_61249_53311# a_61065_53679# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3498 c1_8744_97972# m3_8412_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3499 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3500 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3501 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3502 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3503 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3504 a_n4470_53722# th_dif_sw_0.CKB VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3505 a_67215_57732# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X3506 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3507 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3508 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X3509 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3510 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3511 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3512 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3513 a_68133_61624# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X3514 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3515 c1_42632_21618# m3_42300_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3516 a_66368_52081# a_66216_52022# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X3517 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3518 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X3519 a_62527_56974# a_61929_56639# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3520 a_67431_61671# a_67105_61303# a_67310_61352# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X3521 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3522 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3523 VDDD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3524 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_110450# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3525 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3526 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3527 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3528 a_64761_51028# a_64199_50761# a_64428_50947# VDDD sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X3529 a_66785_50875# a_66593_50645# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.14 as=0.1302 ps=1.195 w=0.84 l=0.15
X3530 a_62527_51646# a_61929_51311# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3531 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3532 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3533 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3534 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3535 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3536 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3537 a_66773_51977# a_65861_51977# a_66666_51977# VDDD sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X3538 VDDD a_66795_71265# sar10b_0.SWP[6] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3539 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3540 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3541 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3542 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3543 a_66254_57356# a_65865_57675# a_65589_57735# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X3544 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3545 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3546 a_62185_66027# sar10b_0.net12 a_62706_65967# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3547 sar10b_0._16_ a_67372_52833# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2997 ps=2.29 w=0.74 l=0.15
X3548 sar10b_0._13_ a_67439_50041# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1988 ps=1.505 w=1.12 l=0.15
X3549 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3550 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3551 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3552 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3553 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3554 sar10b_0.clknet_0_CLK a_65577_51311# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X3555 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3556 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3557 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3558 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3559 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3560 a_62222_57356# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X3561 a_61153_58263# a_60969_57971# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3562 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3563 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3564 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3565 sar10b_0.net3 a_60690_49683# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3566 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3567 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X3568 VSSR sar10b_0.SWN[4] a_25137_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3569 VDDD sar10b_0.net5 a_60969_56639# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X3570 a_64238_63682# a_64033_63591# a_63573_63303# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X3571 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3572 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3573 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3574 VSSD tdc_0.OUTN a_60690_54641# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X3575 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3576 a_31680_111642# sar10b_0.CF[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X3577 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3578 c1_n1140_27218# m3_n1472_27178# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3579 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3580 a_62181_56768# a_61929_56639# a_62319_56646# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X3581 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3582 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3583 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3584 VSSA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3585 VDDA tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.pd_out_0.B VDDA sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X3586 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3587 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3588 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3589 VDDD sar10b_0.net16 a_62997_67299# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X3590 a_66159_65970# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X3591 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3592 VSSD sar10b_0.net16 a_65676_69723# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3593 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3594 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3595 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3596 a_15533_113041# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3597 a_60780_57975# sar10b_0.net7 a_60693_57975# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3598 a_67598_58688# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X3599 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X3600 a_62706_65967# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3601 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3602 VSSD a_66079_59638# sar10b_0.net34 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3603 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3604 VDDD a_67881_60339# a_68133_60292# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X3605 VDDD a_65983_64966# sar10b_0.net44 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X3606 VDDD sar10b_0.net16 a_65397_56643# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X3607 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3608 a_n4470_53722# th_dif_sw_0.CKB VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X3609 a_68421_54964# a_68169_55011# a_68559_55068# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X3610 VDDA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VDDA sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3611 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3612 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3613 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3614 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3615 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X3616 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3617 VSSD sar10b_0.net23 a_68946_59303# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X3618 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3619 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X3620 VSSD sar10b_0.clk_div_0.COUNT\[2\] a_68384_51373# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.111 ps=1.045 w=0.64 l=0.15
X3621 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3622 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3623 a_68169_59007# a_67209_59007# a_67733_58787# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X3624 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3625 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3626 a_61347_49986# a_61086_49986# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X3627 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X3628 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3629 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X3630 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3631 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3632 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3633 a_68371_54656# a_67393_54643# a_68169_55011# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X3634 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3635 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3636 VDDD sar10b_0.net4 a_63273_67295# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X3637 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3638 a_61153_56931# a_60969_56639# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3639 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3640 a_5929_113881# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3641 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3642 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3643 c1_45456_54098# m3_45124_54058# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3644 VDDA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3645 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_110450# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3646 a_61153_51603# a_60969_51311# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3647 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3648 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3649 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3650 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3651 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3652 a_65676_69723# sar10b_0.net2 a_65589_69723# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X3653 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3654 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3655 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3656 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3657 a_62319_57978# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X3658 a_9853_112162# sar10b_0.SWP[7] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3659 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3660 VDDD a_68169_66999# a_68421_66952# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X3661 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3662 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3663 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X3664 a_62185_62031# a_61395_61948# a_61677_62178# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X3665 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3666 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3667 VDDA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3668 a_6634_111636# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X3669 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3670 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3671 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3672 VDDD a_69003_71265# sar10b_0.SWP[8] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3673 VSSR sar10b_0.SWN[5] a_20335_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3674 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3675 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X3676 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3677 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3678 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3679 DATA[9] a_68946_68627# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3680 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3681 VSSD sar10b_0._11_ a_64338_52411# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X3682 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3683 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3684 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3685 a_66216_49358# a_65861_49313# a_66109_49318# VDDD sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X3686 th_dif_sw_0.VCP th_dif_sw_0.th_sw_1.CK th_dif_sw_0.VCP VSSA sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=17.4 ps=121.74 w=20 l=0.15
X3687 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3688 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X3689 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_109594# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3690 a_61448_57022# a_60969_56639# a_61358_57022# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X3691 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3692 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3693 VSSR sar10b_0.SWN[3] a_29939_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3694 a_66035_53072# a_65394_52643# a_65928_53032# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X3695 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3696 VDDA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3697 a_65198_66346# a_64993_66255# a_64533_65967# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X3698 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3699 VSSD a_66762_50329# a_66961_50219# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1229 pd=1.085 as=0.1824 ps=1.85 w=0.64 l=0.15
X3700 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3701 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3702 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3703 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3704 a_63339_71265# sar10b_0.net41 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3705 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3706 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3707 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3708 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3709 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3710 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3711 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3712 a_61609_63602# a_61400_63620# a_60945_63273# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X3713 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3714 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3715 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3716 VDDD a_63509_62783# a_63464_62684# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X3717 a_61358_57022# a_60969_56639# a_60693_56643# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X3718 a_61493_58256# a_61358_58354# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X3719 VDDD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3720 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3721 VSSD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3722 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3723 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3724 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3725 c1_20040_97972# m3_19708_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3726 a_25137_112201# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3727 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3728 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3729 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3730 VSSD sar10b_0.net3 a_66732_61731# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X3731 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3732 a_61349_50398# a_61086_49986# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X3733 a_62007_63363# a_61609_63602# a_61929_63363# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X3734 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3735 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_110450# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3736 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3737 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3738 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3739 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3740 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X3741 VSSA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3742 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3743 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3744 VDDD sar10b_0.net13 a_65001_68627# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X3745 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3746 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3747 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3748 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3749 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3750 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3751 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3752 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3753 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3754 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3755 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3756 c1_45456_22738# m3_45124_22698# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3757 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X3758 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3759 a_68767_66644# a_68169_66999# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X3760 a_19457_110450# sar10b_0.SWP[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3761 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3762 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3763 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3764 a_65000_59686# a_64521_59303# a_64910_59686# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X3765 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3766 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3767 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3768 a_n8277_65767# VDDA th_dif_sw_0.th_sw_1.th_sw_main_0.VGS VSSA sky130_fd_pr__nfet_01v8 ad=2.175 pd=15.58 as=2.175 ps=15.58 w=7.5 l=0.15
X3769 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3770 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3771 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3772 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3773 a_16238_111636# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X3774 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3775 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3776 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3777 a_63464_62684# a_62985_63003# a_63374_62684# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X3778 a_67598_68012# a_67393_67963# a_66933_68391# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X3779 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3780 c1_n1140_67732# m3_n1472_67692# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3781 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3782 VDDD sar10b_0.clk_div_0.COUNT\[1\] a_68035_50645# VDDD sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X3783 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X3784 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3785 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3786 VSSD a_61395_60616# a_61400_60956# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X3787 VSSD sar10b_0.net16 a_63573_63003# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X3788 sar10b_0.clknet_0_CLK a_65577_51311# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3789 a_9853_112162# sar10b_0.SWP[7] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3790 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3791 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3792 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3793 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A a_7670_111642# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3794 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3795 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_109594# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3796 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3797 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3798 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3799 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3800 c1_n1140_44018# m3_n1472_43978# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3801 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3802 sar10b_0.clknet_0_CLK a_65577_51311# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3803 a_61929_63363# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X3804 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3805 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3806 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3807 a_68169_68331# a_67393_67963# a_67733_68111# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X3808 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3809 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3810 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3811 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3812 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3813 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3814 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3815 sar10b_0.net4 a_60690_53975# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3816 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3817 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3818 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3819 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3820 VSSD a_68235_71265# sar10b_0.SWP[7] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X3821 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3822 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3823 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3824 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3825 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3826 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3827 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3828 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3829 a_68767_65312# a_68169_65667# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X3830 a_67035_57732# a_65865_57675# a_66825_57675# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X3831 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3832 VDDD a_67733_58787# a_67688_58688# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X3833 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3834 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3835 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3836 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3837 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X3838 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y sar10b_0.CF[2] VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3839 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3840 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3841 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3842 c1_3096_21618# m3_2764_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3843 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3844 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3845 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3846 a_29061_5788# sar10b_0.SWN[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3847 sar10b_0.net13 a_60747_65937# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X3848 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3849 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3850 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3851 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3852 a_19457_5788# sar10b_0.SWN[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3853 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3854 VDDD sar10b_0.net16 a_61182_52404# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X3855 a_63573_63003# a_63509_62783# a_63495_63003# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X3856 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3857 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3858 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3859 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3860 c1_14392_21618# m3_14060_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3861 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X3862 VDDD a_60690_49683# sar10b_0.net3 VDDD sky130_fd_pr__pfet_01v8 ad=0.1876 pd=1.455 as=0.168 ps=1.42 w=1.12 l=0.15
X3863 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3864 a_64188_51135# sar10b_0.clknet_1_0__leaf_CLK VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3865 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3866 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3867 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3868 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3869 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X3870 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3871 VDDD a_67077_57628# a_67027_57320# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X3872 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3873 a_61153_67587# a_60969_67295# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X3874 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3875 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X3876 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3877 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3878 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3879 VSSD a_61131_70891# sar10b_0.SWP[0] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X3880 a_67077_57628# a_66825_57675# a_67215_57732# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X3881 VSSD a_60747_64231# sar10b_0.CF[6] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X3882 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3883 a_62185_63363# a_61400_63620# a_61677_63510# VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X3884 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3885 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3886 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y sar10b_0.CF[9] VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3887 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3888 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3889 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3890 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3891 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3892 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3893 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3894 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3895 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X3896 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3897 a_n9133_57045# th_dif_sw_0.th_sw_1.CKB a_n8277_54249# VSSA sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X3898 a_9853_112162# sar10b_0.SWP[7] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3899 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3900 VSSD sar10b_0.cyclic_flag_0.FINAL a_67113_56343# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X3901 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3902 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3903 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X3904 a_67688_58688# a_67209_59007# a_67598_58688# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X3905 a_19457_110450# sar10b_0.SWP[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3906 VDDA th_dif_sw_0.CK a_n4470_65264# VDDA sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3907 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3908 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3909 a_65683_59722# a_64705_59595# a_65481_59303# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X3910 VSSD sar10b_0.net3 a_67797_59007# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X3911 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A a_17274_111642# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X3912 a_67393_67963# a_67209_68331# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X3913 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3914 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3915 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X3916 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3917 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X3918 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3919 a_66163_69046# a_65185_68919# a_65961_68627# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X3920 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X3921 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3922 a_63495_63003# a_63169_62635# a_63374_62684# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X3923 a_n4470_65264# th_dif_sw_0.CK VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3924 VSSA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3925 a_63573_63303# sar10b_0.net2 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X3926 VSSR sar10b_0.SWN[8] a_5929_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3927 a_67598_62684# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X3928 VSSD sar10b_0.net27 a_68946_68627# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X3929 VDDD a_60747_68227# sar10b_0.CF[8] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X3930 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3931 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3932 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X3933 a_68169_68331# a_67209_68331# a_67733_68111# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X3934 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3935 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3936 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3937 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3938 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X3939 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3940 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3941 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3942 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3943 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3944 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3945 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3946 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3947 a_67023_56646# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X3948 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 a_9853_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3949 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3950 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3951 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3952 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3953 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3954 VSSD sar10b_0._07_ a_64454_51311# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.19013 pd=1.345 as=0.08663 ps=0.865 w=0.55 l=0.15
X3955 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3956 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3957 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X3958 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3959 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3960 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3961 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X3962 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3963 a_24259_109594# sar10b_0.SWP[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3964 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3965 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3966 a_19457_5788# sar10b_0.SWN[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3967 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3968 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X3969 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3970 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3971 a_1127_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3972 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3973 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3974 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3975 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3976 VDDA th_dif_sw_0.CKB a_n4470_53722# VDDA sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X3977 a_68235_48621# sar10b_0.net35 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X3978 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X3979 a_67797_59007# a_67733_58787# a_67719_59007# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X3980 a_62901_61671# a_62837_61451# a_62823_61671# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X3981 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3982 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3983 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3984 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3985 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X3986 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3987 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X3988 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3989 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X3990 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X3991 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X3992 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3993 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X3994 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3995 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3996 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X3997 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X3998 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X3999 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4000 a_n4470_53722# th_dif_sw_0.CKB VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4001 VDDD a_64238_67295# a_64492_67433# VDDD sky130_fd_pr__pfet_01v8 ad=0.1638 pd=1.275 as=0.1176 ps=0.98 w=0.42 l=0.15
X4002 VDDR sar10b_0.CF[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4003 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4004 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4005 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4006 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y sar10b_0.CF[7] VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4007 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4008 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4009 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4010 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4011 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4012 VDDA th_dif_sw_0.CKB a_n4470_53722# VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4013 VSSD sar10b_0.clknet_0_CLK a_65355_53949# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X4014 a_62139_57978# a_60969_57971# a_61929_57971# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X4015 a_64245_59307# sar10b_0.net1 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X4016 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4017 a_66079_59638# a_65481_59303# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X4018 a_19457_110450# sar10b_0.SWP[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4019 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4020 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4021 a_61609_64934# a_61395_64612# a_60945_64605# VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X4022 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4023 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4024 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4025 a_n4470_53722# th_dif_sw_0.CKB VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4026 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4027 VSSD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X4028 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4029 c1_n1140_84532# m3_n1472_84492# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4030 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4031 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4032 a_64935_64695# a_64609_64923# a_64814_65014# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4033 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X4034 a_67719_59007# a_67393_58639# a_67598_58688# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4035 a_62823_61671# a_62497_61303# a_62702_61352# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4036 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4037 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4038 VDDA th_dif_sw_0.CKB a_n4470_53722# VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4039 VSSR sar10b_0.SWP[3] a_29939_111781# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4040 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4041 a_61493_67580# a_61358_67678# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X4042 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_111306# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4043 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4044 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4045 VSSR sar10b_0.SWN[5] a_20335_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4046 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4047 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4048 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X4049 a_n4470_53722# th_dif_sw_0.CKB VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4050 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4051 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4052 a_24259_109594# sar10b_0.SWP[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4053 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4054 a_60747_65563# sar10b_0.net12 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X4055 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4056 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4057 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4058 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4059 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4060 VDDR sar10b_0.CF[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X4061 c1_45456_62132# m3_45124_62092# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4062 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4063 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4064 c1_n1140_29458# m3_n1472_29418# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4065 VSSR sar10b_0.SWN[3] a_29939_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4066 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4067 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X4068 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4069 VSSA th_dif_sw_0.VCP a_51603_58977# VSSA sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X4070 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4071 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4072 a_29061_5788# sar10b_0.SWN[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4073 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4074 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4075 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4076 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4077 a_20335_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4078 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4079 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4080 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4081 VDDD a_66785_50875# sar10b_0.net16 VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4082 a_24259_5788# sar10b_0.SWN[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4083 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4084 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4085 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4086 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4087 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y a_45050_8706# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X4088 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4089 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4090 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4091 c1_24276_97972# m3_23944_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4092 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X4093 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4094 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4095 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4096 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4097 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4098 c1_45456_77812# m3_45124_77772# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4099 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4100 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4101 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4102 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4103 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4104 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4105 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4106 a_66482_50006# a_65957_50273# a_66312_50368# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X4107 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4108 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X4109 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4110 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4111 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4112 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4113 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4114 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4115 VDDD a_62277_50968# a_62227_50660# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X4116 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4117 VDDD a_61773_52237# a_61705_51992# VDDD sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X4118 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4119 a_61041_52340# a_61496_52091# a_61445_51992# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X4120 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4121 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4122 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4123 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4124 VDDD sar10b_0._06_ a_67890_69727# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X4125 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4126 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4127 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4128 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4129 VDDD tdc_0.OUTP a_60690_70625# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3528 ps=2.87 w=1.12 l=0.15
X4130 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4131 VDDA tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.pd_out_0.A VDDA sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.15
X4132 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4133 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4134 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4135 VDDD sar10b_0.net24 a_68946_61735# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X4136 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4137 a_68421_65620# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X4138 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4139 a_66559_68962# a_65961_68627# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4140 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X4141 a_66825_69663# a_66049_69295# a_66389_69443# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X4142 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4143 a_65769_65963# a_64809_65963# a_65333_66248# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X4144 a_65983_64966# a_65385_64631# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4145 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4146 VDDD a_67733_62783# a_67688_62684# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X4147 VDDA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VDDA sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4148 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4149 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4150 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4151 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4152 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4153 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4154 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4155 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4156 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4157 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4158 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 a_9853_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4159 VDDD sar10b_0.cyclic_flag_0.FINAL a_66921_61671# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4160 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4161 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4162 VDDD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.1736 pd=1.43 as=0.168 ps=1.42 w=1.12 l=0.15
X4163 VDDD a_64485_56768# a_64435_57058# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X4164 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X4165 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4166 c1_n1140_31698# m3_n1472_31658# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4167 VSSD a_66080_53027# a_66098_52670# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X4168 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4169 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4170 a_62702_61352# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X4171 c1_1684_21618# m3_1352_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4172 a_66027_53575# sar10b_0._17_ VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X4173 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4174 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4175 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4176 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4177 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4178 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4179 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4180 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4181 VDDA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4182 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4183 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X4184 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4185 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4186 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4187 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4188 c1_12980_21618# m3_12648_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4189 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4190 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4191 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4192 VSSD a_69003_48621# sar10b_0.SWN[8] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4193 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4194 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4195 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4196 VSSD sar10b_0.net16 a_62325_56343# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X4197 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4198 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4199 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4200 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4201 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4202 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4203 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4204 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4205 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4206 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4207 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4208 DATA[3] a_68946_53975# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4209 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4210 a_67688_62684# a_67209_63003# a_67598_62684# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X4211 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4212 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4213 VDDA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4214 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4215 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4216 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4217 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4218 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4219 VSSD sar10b_0.net3 a_67797_63003# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X4220 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4221 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4222 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4223 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4224 a_62415_51072# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X4225 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4226 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4227 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4228 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4229 a_62798_58688# a_62409_59007# a_62133_59067# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4230 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4231 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X4232 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4233 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4234 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4235 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4236 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4237 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4238 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4239 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4240 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4241 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4242 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4243 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4244 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4245 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4246 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4247 a_64780_52239# a_64924_52385# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1248 pd=1.03 as=0.1696 ps=1.81 w=0.64 l=0.15
X4248 VDDD sar10b_0.net16 a_61461_56403# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X4249 c1_45456_24978# m3_45124_24938# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4250 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4251 VDDA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4252 VSSR sar10b_0.SWP[5] a_20335_112621# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4253 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X4254 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4255 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4256 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4257 a_66843_56646# a_65673_56639# a_66633_56639# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X4258 a_62325_56343# a_62261_56123# a_62247_56343# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4259 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4260 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4261 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4262 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4263 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4264 VDDD a_68133_61624# a_68083_61316# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X4265 c1_n1140_69972# m3_n1472_69932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4266 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4267 VSSD sar10b_0.net47 a_68946_71059# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X4268 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4269 VDDD sar10b_0._10_ a_67084_53565# VDDD sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.147 ps=1.19 w=0.84 l=0.15
X4270 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4271 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4272 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4273 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4274 a_67797_63003# a_67733_62783# a_67719_63003# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4275 VSSR sar10b_0.SWN[4] a_25137_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4276 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4277 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4278 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4279 a_14655_111306# sar10b_0.SWP[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4280 c1_n1140_46258# m3_n1472_46218# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4281 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4282 VDDD a_67637_56123# a_67592_56024# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X4283 VDDD sar10b_0.net14 a_65673_56639# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4284 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4285 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4286 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4287 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4288 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4289 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4290 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4291 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4292 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4293 a_24259_5788# sar10b_0.SWN[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4294 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4295 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4296 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X4297 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4298 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4299 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4300 VSSR sar10b_0.SWP[4] a_25137_112201# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4301 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4302 VSSD a_61773_52237# a_61705_51992# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X4303 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4304 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4305 a_15533_113041# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4306 VDDD a_65385_64631# a_65637_64760# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X4307 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4308 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4309 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4310 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4311 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4312 c1_45456_94612# m3_45124_94572# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4313 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4314 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4315 a_61249_53311# a_61065_53679# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X4316 VDDD sar10b_0.cyclic_flag_0.FINAL a_67209_55011# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4317 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4318 a_65480_69010# a_65001_68627# a_65390_69010# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X4319 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4320 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4321 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4322 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4323 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4324 VDDD a_62527_58306# sar10b_0.net8 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X4325 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4326 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4327 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4328 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4329 a_67719_63003# a_67393_62635# a_67598_62684# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4330 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4331 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4332 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4333 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4334 VDDD sar10b_0.net16 a_61086_65970# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X4335 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4336 sar10b_0.net3 a_60690_49683# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4337 a_65188_51977# sar10b_0._10_ VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0.165 ps=1.33 w=1 l=0.15
X4338 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4339 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4340 a_67592_56024# a_67113_56343# a_67502_56024# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X4341 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4342 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4343 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4344 VSSD sar10b_0.net4 a_61065_53679# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X4345 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4346 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4347 a_61677_62178# a_61395_61948# a_62038_62350# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X4348 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4349 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4350 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4351 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4352 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[4] a_26878_8700# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X4353 VDDD a_61589_53459# a_61544_53360# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X4354 c1_45456_39538# m3_45124_39498# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4355 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4356 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4357 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4358 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4359 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4360 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4361 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4362 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4363 a_67310_61352# a_66921_61671# a_66645_61731# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4364 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4365 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4366 VSSD a_65643_71265# sar10b_0.SWP[5] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4367 VSSA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4368 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4369 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4370 a_60780_67299# sar10b_0.net13 a_60693_67299# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X4371 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X4372 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4373 a_65765_50645# a_65586_50645# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2516 pd=2.16 as=0.17575 ps=1.215 w=0.74 l=0.15
X4374 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4375 a_61491_52222# sar10b_0.net4 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X4376 VDDD sar10b_0.net11 a_62185_64695# VDDD sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X4377 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4378 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4379 VSSR sar10b_0.SWP[3] a_29939_111781# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4380 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4381 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4382 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4383 a_68331_52243# sar10b_0._13_ VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4384 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4385 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X4386 a_62185_63363# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X4387 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4388 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4389 VSSR sar10b_0.SWN[5] a_20335_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4390 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4391 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4392 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4393 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4394 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4395 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4396 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4397 VSSD a_65577_51311# sar10b_0.clknet_0_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X4398 a_62527_58306# a_61929_57971# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4399 VSSD a_60747_69559# sar10b_0.CF[9] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4400 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4401 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4402 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=3.48 ps=37.92 w=0.5 l=0.5
X4403 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4404 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4405 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4406 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4407 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4408 VDDD a_66961_50219# a_66869_50413# VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.09975 ps=0.895 w=0.42 l=0.15
X4409 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4410 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4411 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4412 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4413 a_68767_54656# a_68169_55011# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X4414 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4415 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4416 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4417 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4418 VDDD a_66389_69443# a_66344_69344# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X4419 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 a_5051_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4420 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4421 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4422 c1_22864_97972# m3_22532_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4423 sar10b_0._09_ a_64454_51311# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.2382 ps=1.555 w=1.12 l=0.15
X4424 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4425 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4426 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4427 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4428 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4429 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4430 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4431 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4432 a_51861_60437# th_dif_sw_0.VCP VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X4433 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4434 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4435 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4436 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4437 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4438 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4439 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4440 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4441 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4442 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4443 VDDD sar10b_0.net47 a_68946_71059# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X4444 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4445 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4446 a_64356_51029# a_64199_50761# a_63918_50969# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1181 ps=1.035 w=0.55 l=0.15
X4447 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4448 a_51603_58977# CLK a_51345_58977# VSSA sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X4449 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4450 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4451 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X4452 c1_n1140_71092# m3_n1472_71052# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4453 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4454 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X4455 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4456 a_65775_64638# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X4457 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4458 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4459 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4460 c1_34160_21618# m3_33828_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4461 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4462 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4463 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4464 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4465 a_65119_59984# a_64521_60339# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4466 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4467 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4468 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4469 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4470 a_62126_56024# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X4471 a_63662_57022# a_63457_56931# a_62997_56643# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X4472 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=3.48 ps=28.64 w=1.5 l=0.5
X4473 c1_45456_41778# m3_45124_41738# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4474 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4475 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4476 VSSD a_66464_50363# a_66482_50006# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.0441 ps=0.63 w=0.42 l=0.15
X4477 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y a_16238_8706# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X4478 VSSD a_64543_62648# sar10b_0.net42 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4479 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4480 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4481 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4482 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4483 VSSD sar10b_0.net5 a_60969_56639# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X4484 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4485 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X4486 c1_n1140_86772# m3_n1472_86732# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4487 a_62038_53026# a_61609_52946# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X4488 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4489 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4490 a_20335_112621# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4491 VDDA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VDDA sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4492 VSSD sar10b_0.net5 a_60969_51311# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X4493 VSSD a_63045_57628# a_63003_57732# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X4494 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4495 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4496 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4497 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4498 a_65643_48621# sar10b_0.net33 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X4499 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4500 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4501 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4502 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4503 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4504 a_1832_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4505 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4506 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4507 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4508 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4509 a_61677_62178# a_61400_62288# a_62007_62031# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X4510 a_63871_61316# a_63273_61671# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X4511 a_61419_48621# sar10b_0.net17 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4512 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4513 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4514 a_67105_61303# a_66921_61671# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X4515 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X4516 a_61153_58263# a_60969_57971# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X4517 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4518 a_62025_53679# a_61065_53679# a_61589_53459# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X4519 VDDA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4520 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4521 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4522 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4523 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4524 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4525 c1_45456_64372# m3_45124_64332# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4526 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4527 a_68559_65724# sar10b_0.net3 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X4528 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4529 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4530 a_66109_51982# sar10b_0._04_ VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X4531 a_62235_51072# a_61065_51015# a_62025_51015# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X4532 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4533 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X4534 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4535 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4536 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4537 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4538 VDDD a_64428_50947# a_64356_51029# VDDD sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.2331 ps=1.395 w=0.84 l=0.15
X4539 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4540 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4541 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4542 a_25137_112201# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4543 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4544 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4545 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X4546 a_9853_5788# sar10b_0.SWN[7] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4547 a_62185_60699# a_61395_60616# a_61677_60846# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X4548 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4549 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4550 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4551 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4552 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4553 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4554 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X4555 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4556 VDDD a_63871_61316# sar10b_0.net41 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X4557 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4558 a_64437_63363# a_64373_63584# a_64359_63363# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4559 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4560 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4561 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4562 VSSD a_64428_50947# a_64356_51029# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1648 pd=1.245 as=0.10905 ps=1.025 w=0.55 l=0.15
X4563 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4564 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4565 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4566 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4567 VSSD a_68767_58652# sar10b_0.net19 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4568 VSSD sar10b_0.net16 a_65109_59367# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X4569 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A a_2868_111642# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X4570 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4571 a_62277_50968# a_62025_51015# a_62415_51072# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X4572 c1_45456_56338# m3_45124_56298# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4573 VSSA th_dif_sw_0.VCN a_51603_61205# VSSA sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=1
X4574 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4575 a_63339_71265# sar10b_0.net41 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4576 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4577 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4578 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4579 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_111306# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4580 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4581 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_109594# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4582 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4583 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X4584 a_62227_50660# a_61249_50647# a_62025_51015# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X4585 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4586 sar10b_0.clknet_0_CLK a_65577_51311# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4587 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4588 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4589 VDDD a_61491_52222# a_61496_52091# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4590 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4591 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X4592 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4593 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X4594 a_61493_51596# a_61358_51694# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X4595 a_67393_65299# a_67209_65667# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X4596 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4597 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4598 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4599 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4600 VSSD a_62277_53632# a_62235_53736# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X4601 VSSD a_67135_58306# sar10b_0.net36 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4602 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X4603 VDDD sar10b_0.cyclic_flag_0.FINAL a_67209_64335# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X4604 a_62793_57675# a_61833_57675# a_62357_57455# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X4605 a_64359_63363# a_64033_63591# a_64238_63682# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4606 a_65481_59303# a_64705_59595# a_65045_59588# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X4607 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4608 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4609 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4610 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4611 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4612 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4613 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4614 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4615 VDDD a_62527_67630# sar10b_0.net14 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X4616 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4617 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4618 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4619 a_65109_59367# a_65045_59588# a_65031_59367# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4620 VSSD sar10b_0.net16 a_65397_66027# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X4621 a_67733_64115# a_67598_64016# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X4622 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4623 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4624 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4625 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4626 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y sar10b_0.CF[0] VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4627 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4628 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4629 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4630 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4631 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X4632 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4633 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X4634 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4635 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4636 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4637 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4638 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4639 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4640 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4641 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4642 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4643 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4644 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4645 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4646 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4647 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4648 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4649 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4650 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X4651 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4652 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4653 VSSD CLK a_65577_51311# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.063 pd=0.72 as=0.0588 ps=0.7 w=0.42 l=0.15
X4654 c1_18628_97972# m3_18296_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4655 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4656 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4657 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4658 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4659 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4660 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4661 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4662 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4663 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4664 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4665 c1_44044_97972# m3_43712_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4666 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4667 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4668 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4669 a_64238_63682# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X4670 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4671 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4672 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4673 a_29061_5788# sar10b_0.SWN[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4674 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4675 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4676 a_68169_66999# a_67393_66631# a_67733_66779# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X4677 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4678 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4679 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4680 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4681 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4682 a_65397_66027# a_65333_66248# a_65319_66027# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4683 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4684 a_53652_61050# tdc_0.phase_detector_0.INN VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.15
X4685 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4686 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4687 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4688 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4689 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4690 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4691 VSSD sar10b_0._08_ sar10b_0._04_ VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4692 tdc_0.RDY tdc_0.phase_detector_0.pd_out_0.B a_55382_59612# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.0888 ps=0.98 w=0.74 l=0.15
X4693 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4694 a_68421_54964# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X4695 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4696 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4697 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4698 VSSD a_67231_56974# sar10b_0.net37 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4699 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4700 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4701 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4702 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4703 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4704 sar10b_0.clk_div_0.COUNT\[3\] a_66577_52883# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X4705 VSSR sar10b_0.SWP[3] a_29939_111781# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4706 a_65957_50273# a_65778_49979# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X4707 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4708 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4709 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4710 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=10.44 ps=85.92 w=1.5 l=0.5
X4711 a_5051_113018# sar10b_0.SWP[8] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4712 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4713 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4714 VSSR sar10b_0.SWN[5] a_20335_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4715 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4716 VSSD sar10b_0.cyclic_flag_0.FINAL a_67209_68331# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X4717 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4718 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4719 a_65021_50292# sar10b_0._08_ a_64907_50292# VDDD sky130_fd_pr__pfet_01v8 ad=0.1703 pd=1.355 as=0.21 ps=1.42 w=1 l=0.15
X4720 a_66109_51982# sar10b_0._04_ VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
X4721 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4722 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4723 VDDD a_62187_48621# sar10b_0.SWN[2] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X4724 a_61173_60642# a_60945_60609# a_61086_60642# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X4725 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X4726 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4727 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4728 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4729 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4730 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4731 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4732 c1_45456_81172# m3_45124_81132# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4733 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4734 a_63374_62684# a_62985_63003# a_62709_63063# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4735 c1_n1140_48498# m3_n1472_48458# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4736 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4737 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X4738 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4739 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4740 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4741 a_14655_5788# sar10b_0.SWN[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4742 VSSR sar10b_0.SWN[3] a_29939_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4743 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4744 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4745 a_65319_66027# a_64993_66255# a_65198_66346# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X4746 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4747 VSSR sar10b_0.CF[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4748 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4749 a_64910_59686# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X4750 DATA[2] a_68946_52411# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4751 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X4752 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4753 a_20335_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4754 a_66294_51051# a_65765_50645# a_66103_50668# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07568 ps=0.83 w=0.42 l=0.15
X4755 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4756 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4757 a_55382_59612# tdc_0.phase_detector_0.pd_out_0.A VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.12607 ps=1.1 w=0.74 l=0.15
X4758 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X4759 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4760 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4761 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4762 a_67393_66631# a_67209_66999# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X4763 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4764 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4765 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4766 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4767 a_62261_56123# a_62126_56024# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X4768 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4769 c1_45456_96852# m3_45124_96812# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4770 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y sar10b_0.CF[5] VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X4771 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4772 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4773 a_60945_60609# a_61395_60616# a_61347_60642# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X4774 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4775 c1_45456_26098# m3_45124_26058# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4776 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X4777 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4778 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4779 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4780 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4781 a_66197_56924# a_66062_57022# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X4782 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4783 a_66485_53077# a_65573_52937# a_66378_52993# VDDD sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X4784 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4785 a_61086_64638# a_60945_64605# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X4786 VDDA CLK a_51345_60437# VDDA sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=1
X4787 c1_38396_21618# m3_38064_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4788 VSSA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4789 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4790 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4791 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4792 VDDD a_64233_56639# a_64485_56768# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X4793 a_65637_64760# a_65385_64631# a_65775_64638# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X4794 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4795 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4796 a_29061_108738# sar10b_0.SWP[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4797 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4798 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4799 a_65198_66346# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X4800 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4801 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X4802 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X4803 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4804 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4805 a_61609_52946# a_61400_52964# a_60945_52617# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X4806 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4807 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4808 a_21040_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X4809 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4810 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4811 VSSD a_64485_56768# a_64443_56646# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X4812 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4813 a_14655_111306# sar10b_0.SWP[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4814 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4815 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS VDDA a_n8277_54565# VSSA sky130_fd_pr__nfet_01v8 ad=2.175 pd=15.58 as=2.175 ps=15.58 w=7.5 l=0.15
X4816 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4817 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4818 a_67423_69308# a_66825_69663# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4819 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4820 a_24259_109594# sar10b_0.SWP[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4821 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4822 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4823 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4824 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4825 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4826 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4827 a_64814_65014# a_64425_64631# a_64149_64635# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4828 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4829 a_60693_56643# sar10b_0.net2 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X4830 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X4831 a_67598_58688# a_67209_59007# a_66933_59067# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4832 a_62702_61352# a_62313_61671# a_62037_61731# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X4833 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4834 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4835 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4836 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4837 VSSR sar10b_0.SWN[3] a_29939_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4838 VDDD sar10b_0.net16 a_61086_63306# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X4839 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4840 a_62185_60699# a_61400_60956# a_61677_60846# VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X4841 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4842 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4843 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X4844 VSSD a_66027_53575# sar10b_0._05_ VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X4845 a_52504_59293# tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A a_52417_59293# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.1824 ps=1.85 w=0.64 l=0.15
X4846 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4847 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4848 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4849 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4850 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4851 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4852 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4853 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4854 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4855 sar10b_0.net7 a_60843_52216# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X4856 sar10b_0.cyclic_flag_0.FINAL a_64888_67630# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3584 ps=2.88 w=1.12 l=0.15
X4857 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4858 VDDD a_68421_65620# a_68371_65312# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X4859 VSSD a_68767_62648# sar10b_0.net24 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4860 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4861 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4862 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4863 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4864 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4865 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4866 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4867 a_67598_68012# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X4868 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X4869 a_64521_60339# a_63561_60339# a_64085_60119# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X4870 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4871 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4872 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4873 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4874 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4875 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4876 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4877 VDDD a_67881_61671# a_68133_61624# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X4878 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4879 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X4880 a_5929_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4881 a_60747_65563# sar10b_0.net12 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4882 VSSD tdc_0.RDY a_60690_53975# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0798 pd=0.8 as=0.126 ps=1.44 w=0.42 l=0.15
X4883 a_29061_108738# sar10b_0.SWP[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4884 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4885 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X4886 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4887 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X4888 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X4889 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4890 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4891 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4892 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4893 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4894 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X4895 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4896 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4897 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4898 VDDD a_66593_50645# a_66785_50875# VDDD sky130_fd_pr__pfet_01v8 ad=0.203 pd=1.505 as=0.126 ps=1.14 w=0.84 l=0.15
X4899 VDDD a_64543_62648# sar10b_0.net42 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X4900 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4901 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X4902 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4903 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4904 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4905 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X4906 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4907 a_65643_48621# sar10b_0.net33 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4908 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4909 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4910 VSSR sar10b_0.SWP[5] a_20335_112621# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4911 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4912 a_64924_52385# sar10b_0._09_ VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.231 pd=2.23 as=0.203 ps=1.505 w=0.84 l=0.15
X4913 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4914 VSSD a_60945_60609# a_60747_60609# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4915 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4916 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4917 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4918 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4919 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4920 a_62319_67302# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X4921 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4922 VDDR sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X4923 a_51603_61205# CLK a_51345_60437# VSSA sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X4924 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4925 DATA[7] a_68946_63299# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X4926 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4927 VDDD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4928 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4929 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 a_249_113874# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4930 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4931 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X4932 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4933 VSSR sar10b_0.SWN[4] a_25137_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4934 a_61153_56931# a_60969_56639# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X4935 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4936 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4937 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4938 a_14655_5788# sar10b_0.SWN[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4939 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4940 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X4941 a_65733_59432# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X4942 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X4943 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X4944 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4945 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X4946 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4947 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X4948 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4949 VSSD a_66593_50645# a_66785_50875# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1147 pd=1.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X4950 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4951 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4952 VDDD a_66666_49313# a_66865_49412# VDDD sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X4953 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4954 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4955 a_63861_56703# a_63797_56924# a_63783_56703# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X4956 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4957 a_66213_68756# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X4958 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X4959 VSSD sar10b_0.net16 a_60780_51315# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4960 VDDD a_65045_59588# a_65000_59686# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X4961 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X4962 a_63660_63303# sar10b_0.net2 a_63573_63303# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X4963 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4964 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4965 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4966 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4967 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4968 tdc_0.phase_detector_0.INN a_52417_59293# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X4969 sar10b_0.net11 a_60747_63273# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X4970 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4971 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X4972 a_67637_56123# a_67502_56024# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X4973 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4974 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X4975 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4976 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4977 a_15533_113041# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4978 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4979 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4980 VSSD sar10b_0.net16 a_64332_59307# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X4981 c1_42632_97972# m3_42300_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4982 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X4983 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X4984 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4985 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4986 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X4987 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4988 a_63295_55988# a_62697_56343# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X4989 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4990 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4991 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X4992 VSSD sar10b_0.clknet_0_CLK a_66153_48647# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.063 pd=0.72 as=0.0588 ps=0.7 w=0.42 l=0.15
X4993 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X4994 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X4995 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4996 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4997 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X4998 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X4999 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5000 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5001 c1_28512_21618# m3_28180_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5002 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5003 a_7670_111642# sar10b_0.CF[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5004 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5005 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5006 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5007 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5008 sar10b_0.net3 a_60690_49683# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5009 VDDD a_68767_58652# sar10b_0.net19 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5010 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5011 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5012 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5013 VSSD a_66795_71265# sar10b_0.SWP[6] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X5014 a_63457_67583# a_63273_67295# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5015 VSSD sar10b_0.clknet_1_1__leaf_CLK a_65586_50645# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.17575 pd=1.215 as=0.2109 ps=2.05 w=0.74 l=0.15
X5016 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5017 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5018 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X5019 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5020 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5021 a_63783_56703# a_63457_56931# a_63662_57022# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X5022 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5023 VDDD a_65333_66248# a_65288_66346# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X5024 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5025 a_67445_60119# a_67310_60020# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5026 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5027 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5028 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5029 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5030 a_65199_63306# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X5031 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5032 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X5033 VSSD sar10b_0.net37 a_68562_49747# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X5034 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5035 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5036 DATA[6] a_68946_61735# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5037 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5038 tdc_0.phase_detector_0.INP a_52417_60961# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1988 ps=1.505 w=1.12 l=0.15
X5039 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5040 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5041 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5042 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5043 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5044 a_62025_51015# a_61249_50647# a_61589_50795# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X5045 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X5046 VSSR sar10b_0.SWP[3] a_29939_111781# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5047 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5048 VSSD sar10b_0.net3 a_66732_60399# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5049 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5050 VSSD sar10b_0.net16 a_65484_56643# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5051 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5052 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5053 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5054 a_68035_50645# sar10b_0.clk_div_0.COUNT\[0\] a_67564_50907# VDDD sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X5055 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5056 VSSR sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5057 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5058 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5059 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5060 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5061 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5062 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5063 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5064 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5065 c1_n1140_33938# m3_n1472_33898# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5066 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5067 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5068 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5069 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5070 VSSR sar10b_0.SWN[7] a_10731_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5071 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5072 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5073 VDDD a_68479_61316# sar10b_0.net22 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5074 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5075 a_67084_53565# sar10b_0._16_ VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.1988 ps=1.505 w=0.84 l=0.15
X5076 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5077 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5078 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5079 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5080 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5081 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5082 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5083 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5084 a_55085_59917# tdc_0.phase_detector_0.pd_out_0.A VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.27 as=0.295 ps=2.59 w=1 l=0.15
X5085 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_109594# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5086 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5087 VSSD sar10b_0.net16 a_61173_60642# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X5088 a_65288_66346# a_64809_65963# a_65198_66346# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X5089 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5090 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5091 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5092 VSSD a_68133_60292# a_68091_60396# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X5093 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5094 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5095 sar10b_0.cyclic_flag_0.FINAL a_64888_67630# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5096 sar10b_0.clknet_0_CLK a_65577_51311# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X5097 VDDD a_67733_68111# a_67688_68012# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X5098 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5099 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5100 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5101 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5102 a_61609_62270# a_61400_62288# a_60945_61941# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X5103 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5104 a_17274_8700# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5105 c1_36984_21618# m3_36652_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5106 a_17274_111642# sar10b_0.CF[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5107 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5108 a_61493_56924# a_61358_57022# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5109 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5110 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5111 VSSD a_66255_50749# a_66294_51051# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.19715 pd=1.365 as=0.0441 ps=0.63 w=0.42 l=0.15
X5112 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5113 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=3.48 ps=28.64 w=1.5 l=0.5
X5114 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5115 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5116 a_29061_108738# sar10b_0.SWP[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5117 a_65484_56643# sar10b_0.net1 a_65397_56643# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5118 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5119 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5120 a_60747_60235# sar10b_0.net8 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X5121 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5122 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5123 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5124 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5125 VDDD a_61395_65944# a_61400_66284# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5126 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5127 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5128 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5129 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5130 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5131 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5132 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5133 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5134 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X5135 a_65185_68919# a_65001_68627# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5136 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5137 a_62527_67630# a_61929_67295# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5138 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X5139 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X5140 VDDD a_61677_66174# a_61609_66266# VDDD sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X5141 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5142 VDDD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5143 a_67598_62684# a_67209_63003# a_66933_63063# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X5144 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5145 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5146 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5147 a_68767_65312# a_68169_65667# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5148 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5149 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5150 DATA[5] a_68946_59303# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5151 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5152 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5153 a_n8277_66083# th_dif_sw_0.th_sw_1.CKB a_n9133_63315# VSSA sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.15
X5154 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5155 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5156 a_67688_68012# a_67209_68331# a_67598_68012# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X5157 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5158 a_20335_112621# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5159 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5160 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 a_249_113874# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5161 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5162 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5163 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X5164 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5165 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5166 VDDD a_65577_51311# sar10b_0.clknet_0_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5167 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5168 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5169 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5170 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5171 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5172 a_65961_68627# a_65001_68627# a_65525_68912# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5173 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5174 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5175 a_61035_48621# sar10b_0.net29 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5176 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5177 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5178 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5179 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5180 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5181 a_63663_61728# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X5182 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5183 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5184 VSSD a_61491_52222# a_61496_52091# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X5185 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5186 a_65961_68627# a_65185_68919# a_65525_68912# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X5187 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5188 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5189 a_249_113874# sar10b_0.SWP[9] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5190 VDDD sar10b_0.net16 a_61677_66174# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X5191 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5192 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5193 VDDD a_60690_53975# sar10b_0.net4 VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5194 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X5195 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5196 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5197 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5198 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5199 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5200 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X5201 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_109594# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5202 a_9853_5788# sar10b_0.SWN[7] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5203 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5204 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5205 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5206 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5207 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5208 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5209 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5210 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5211 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5212 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5213 a_25137_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5214 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5215 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5216 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5217 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5218 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5219 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5220 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5221 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5222 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5223 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X5224 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5225 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5226 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5227 a_65407_63634# a_64809_63299# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5228 a_64491_71265# sar10b_0.net42 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5229 a_19457_5788# sar10b_0.SWN[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5230 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5231 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5232 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5233 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5234 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5235 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5236 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5237 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5238 a_5929_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5239 a_66216_49358# a_65682_49313# a_66109_49318# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.15563 ps=1.215 w=0.42 l=0.15
X5240 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5241 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5242 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5243 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5244 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5245 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5246 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5247 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5248 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5249 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5250 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5251 a_61153_67587# a_60969_67295# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X5252 a_62139_67302# a_60969_67295# a_61929_67295# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X5253 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5254 VDDR sar10b_0.CF[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X5255 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5256 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5257 VDDD a_65119_59984# sar10b_0.net33 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5258 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5259 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5260 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X5261 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5262 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5263 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5264 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5265 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5266 VSSD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X5267 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5268 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X5269 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 a_5051_113018# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5270 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5271 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5272 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5273 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5274 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5275 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5276 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5277 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5278 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5279 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5280 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5281 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5282 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5283 VDDD sar10b_0.net16 a_63573_63303# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X5284 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5285 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5286 c1_n1140_50738# m3_n1472_50698# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5287 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5288 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5289 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5290 c1_11568_21618# m3_11236_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5291 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X5292 a_62357_57455# a_62222_57356# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X5293 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5294 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_109594# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5295 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5296 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5297 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5298 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5299 a_68235_71265# sar10b_0.net45 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X5300 a_65589_69723# sar10b_0.net2 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X5301 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5302 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A a_46086_111642# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5303 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5304 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5305 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5306 c1_3096_97972# m3_2764_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5307 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5308 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5309 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5310 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5311 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5312 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5313 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5314 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5315 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5316 VDDD a_68767_62648# sar10b_0.net24 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5317 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5318 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5319 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5320 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5321 c1_14392_97972# m3_14060_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5322 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5323 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5324 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5325 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5326 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5327 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5328 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5329 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5330 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5331 a_24259_109594# sar10b_0.SWP[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5332 VSSD sar10b_0.net4 a_60969_57971# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X5333 a_15533_113041# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5334 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5335 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5336 a_68479_61316# a_67881_61671# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5337 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5338 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5339 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5340 a_54660_59599# tdc_0.phase_detector_0.pd_out_0.A VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5341 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5342 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5343 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5344 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5345 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5346 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5347 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5348 a_29061_5788# sar10b_0.SWN[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5349 a_64033_63591# a_63849_63299# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X5350 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5351 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[0] a_46086_8700# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5352 c1_n1140_73332# m3_n1472_73292# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5353 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5354 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5355 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5356 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5357 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5358 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5359 a_68073_56343# a_67113_56343# a_67637_56123# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5360 a_61677_60846# a_61400_60956# a_62007_60699# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X5361 VDDD sar10b_0.net16 a_64245_59307# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X5362 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_108738# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5363 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5364 a_67027_57320# a_66049_57307# a_66825_57675# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X5365 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5366 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5367 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5368 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5369 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5370 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5371 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5372 VDDD a_67371_49579# sar10b_0.SWN[6] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X5373 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5374 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5375 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5376 VDDD a_67231_56974# sar10b_0.net37 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5377 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5378 a_64339_51661# sar10b_0.net3 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1595 pd=1.68 as=0.1925 ps=1.8 w=0.55 l=0.15
X5379 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5380 a_62185_52707# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X5381 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5382 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5383 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5384 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5385 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5386 a_62185_64695# sar10b_0.net11 a_62706_64635# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5387 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5388 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5389 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5390 VDDD a_63339_48621# sar10b_0.SWN[3] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X5391 a_61445_51992# a_61182_52404# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X5392 a_60945_65937# a_61400_66284# a_61349_66382# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X5393 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5394 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y sar10b_0.CF[1] VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5395 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5396 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5397 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5398 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5399 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5400 a_67077_57628# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X5401 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5402 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5403 VSSR sar10b_0.SWN[5] a_20335_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5404 a_249_113874# sar10b_0.SWP[9] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5405 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5406 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5407 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5408 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5409 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X5410 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5411 a_67371_49579# sar10b_0.net34 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X5412 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5413 VSSR sar10b_0.SWN[7] a_10731_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5414 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5415 a_61589_53459# a_61454_53360# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X5416 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5417 a_64435_57058# a_63457_56931# a_64233_56639# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X5418 a_60747_64231# sar10b_0.net11 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X5419 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5420 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5421 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5422 c1_45456_66612# m3_45124_66572# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5423 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5424 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5425 VDDD a_68421_54964# a_68371_54656# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X5426 a_64238_63682# a_63849_63299# a_63573_63303# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X5427 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5428 a_249_5788# sar10b_0.SWN[9] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5429 a_67020_55071# sar10b_0.net38 a_66933_55071# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5430 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5431 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5432 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 a_9853_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5433 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5434 a_20335_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5435 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5436 a_60780_56643# sar10b_0.net2 a_60693_56643# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5437 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5438 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5439 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X5440 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5441 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5442 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5443 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5444 a_62706_64635# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5445 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5446 a_24259_109594# sar10b_0.SWP[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5447 a_19457_5788# sar10b_0.SWN[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5448 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5449 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A a_22076_111642# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5450 DATA[9] a_68946_68627# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5451 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5452 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5453 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5454 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5455 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_108738# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5456 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X5457 VDDD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5458 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X5459 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5460 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5461 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5462 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5463 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5464 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5465 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5466 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5467 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5468 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X5469 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5470 VSSD sar10b_0.clk_div_0.COUNT\[3\] a_67552_52656# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.12607 pd=1.1 as=0.0888 ps=0.98 w=0.74 l=0.15
X5471 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5472 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5473 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5474 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5475 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5476 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5477 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5478 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5479 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X5480 a_65031_59367# a_64705_59595# a_64910_59686# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X5481 VSSD sar10b_0.clknet_1_1__leaf_CLK a_65394_52643# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X5482 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5483 CKO a_68562_71291# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5484 VSSD a_68479_59984# sar10b_0.net21 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X5485 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5486 a_67733_62783# a_67598_62684# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5487 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5488 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5489 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X5490 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5491 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5492 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5493 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X5494 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5495 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5496 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5497 sar10b_0.net9 a_60747_60609# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X5498 VDDD sar10b_0.net9 a_62409_59007# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5499 sar10b_0.net2 a_60690_70625# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5500 a_62185_66027# a_61395_65944# a_61677_66174# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X5501 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5502 a_62319_56646# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X5503 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5504 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5505 VDDD a_68169_65667# a_68421_65620# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X5506 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X5507 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5508 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5509 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5510 VSSR sar10b_0.SWN[5] a_20335_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5511 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5512 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5513 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5514 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5515 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5516 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5517 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5518 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5519 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5520 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5521 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5522 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5523 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5524 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 a_9853_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5525 a_67552_52656# sar10b_0._14_ sar10b_0._16_ VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.1554 ps=1.16 w=0.74 l=0.15
X5526 a_68559_55068# sar10b_0.net3 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X5527 a_65589_57735# sar10b_0.net1 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X5528 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5529 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5530 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5531 a_63525_61624# a_63273_61671# a_63663_61728# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X5532 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X5533 a_66645_61731# sar10b_0.net42 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X5534 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5535 a_24259_109594# sar10b_0.SWP[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5536 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5537 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5538 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5539 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5540 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5541 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5542 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5543 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5544 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5545 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5546 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5547 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5548 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5549 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5550 a_66080_53027# a_65928_53032# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X5551 a_61493_56924# a_61358_57022# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X5552 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5553 a_25137_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5554 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X5555 a_63003_57732# a_61833_57675# a_62793_57675# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X5556 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5557 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X5558 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5559 a_61493_51596# a_61358_51694# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X5560 a_65198_66346# a_64809_65963# a_64533_65967# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X5561 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5562 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5563 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5564 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5565 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5566 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5567 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5568 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5569 c1_n1140_90132# m3_n1472_90092# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5570 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5571 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5572 a_24259_5788# sar10b_0.SWN[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5573 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5574 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X5575 a_62007_62031# a_61609_62270# a_61929_62031# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X5576 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5577 VSSD sar10b_0.net16 a_62421_57675# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X5578 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5579 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5580 VSSD sar10b_0.cyclic_flag_0.FINAL a_67209_66999# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X5581 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5582 VSSD a_61677_66174# a_61609_66266# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X5583 a_5929_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5584 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y sar10b_0.CF[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5585 a_66825_69663# a_65865_69663# a_66389_69443# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5586 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5587 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5588 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5589 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5590 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5591 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5592 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5593 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5594 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5595 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5596 a_65068_49569# sar10b_0.net3 a_65236_49657# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1376 ps=1.14 w=0.64 l=0.15
X5597 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5598 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5599 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5600 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5601 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5602 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5603 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5604 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5605 a_62220_59067# sar10b_0.net1 a_62133_59067# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5606 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5607 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5608 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5609 VDDR sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X5610 VSSR sar10b_0.SWP[5] a_20335_112621# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5611 VDDD a_66368_52081# a_66323_51982# VDDD sky130_fd_pr__pfet_01v8 ad=0.18985 pd=1.545 as=0.0504 ps=0.66 w=0.42 l=0.15
X5612 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5613 VDDD a_67372_52243# sar10b_0._07_ VDDD sky130_fd_pr__pfet_01v8 ad=0.2362 pd=1.555 as=0.3304 ps=2.83 w=1.12 l=0.15
X5614 c1_n1140_35058# m3_n1472_35018# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5615 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5616 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5617 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5618 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5619 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5620 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X5621 a_64236_64635# sar10b_0.net2 a_64149_64635# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5622 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5623 VDDD sar10b_0.net7 a_61065_51015# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5624 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5625 VSSD a_64491_48621# sar10b_0.SWN[4] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X5626 a_62038_63682# a_61609_63602# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X5627 c1_1684_97972# m3_1352_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5628 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5629 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5630 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5631 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5632 a_68271_60396# sar10b_0.net3 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X5633 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5634 a_66933_65727# sar10b_0.net45 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X5635 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5636 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5637 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5638 a_61929_62031# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X5639 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X5640 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5641 a_62277_50968# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X5642 a_67419_52937# sar10b_0.clk_div_0.COUNT\[3\] VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3752 pd=2.91 as=0.2352 ps=1.54 w=1.12 l=0.15
X5643 c1_12980_97972# m3_12648_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5644 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5645 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5646 a_249_5788# sar10b_0.SWN[9] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5647 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5648 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5649 a_65857_56931# a_65673_56639# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5650 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5651 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5652 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5653 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5654 c1_45456_83412# m3_45124_83372# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5655 a_64831_56974# a_64233_56639# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X5656 a_61395_65944# sar10b_0.net4 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X5657 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5658 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5659 VDDD a_60945_49953# a_60747_49953# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X5660 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5661 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X5662 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5663 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5664 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5665 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5666 VDDD sar10b_0.net37 a_68562_49747# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X5667 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5668 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5669 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5670 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5671 a_24259_5788# sar10b_0.SWN[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5672 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5673 a_66323_51982# a_65682_51977# a_66216_52022# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.09835 ps=1.005 w=0.42 l=0.15
X5674 a_64233_56639# a_63273_56639# a_63797_56924# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5675 a_15533_113041# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5676 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5677 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5678 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_108738# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5679 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5680 sar10b_0.net12 a_60747_64605# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X5681 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X5682 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5683 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5684 a_65511_68691# a_65185_68919# a_65390_69010# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X5685 a_67393_54643# a_67209_55011# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5686 a_64233_56639# a_63457_56931# a_63797_56924# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X5687 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5688 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5689 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5690 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5691 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5692 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5693 VDDD a_65733_59432# a_65683_59722# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X5694 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5695 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5696 c1_45456_28338# m3_45124_28298# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5697 a_67543_51991# sar10b_0.clk_div_0.COUNT\[1\] VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.195 pd=1.39 as=0.2362 ps=1.555 w=1 l=0.15
X5698 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5699 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5700 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5701 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5702 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5703 VDDD a_61395_49960# a_61400_50300# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X5704 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5705 VDDD a_66213_68756# a_66163_69046# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X5706 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5707 VDDD a_62527_56974# sar10b_0.net38 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5708 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5709 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5710 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5711 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5712 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5713 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5714 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5715 VSSD a_60747_62899# sar10b_0.CF[5] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X5716 VSSD a_68421_64288# a_68379_64392# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X5717 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5718 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5719 a_62185_62031# a_61400_62288# a_61677_62178# VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X5720 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5721 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5722 VDDD a_61677_50190# a_61609_50282# VDDD sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X5723 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5724 a_69003_48621# sar10b_0.net36 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5725 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5726 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5727 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5728 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5729 a_62837_61451# a_62702_61352# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5730 a_67020_64395# sar10b_0.net43 a_66933_64395# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X5731 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5732 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5733 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5734 VSSD a_66865_49412# a_66823_49697# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05565 ps=0.685 w=0.42 l=0.15
X5735 sar10b_0._14_ a_68178_51635# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.15535 ps=1.17 w=0.74 l=0.15
X5736 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5737 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5738 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5739 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5740 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5741 VDDD sar10b_0.net10 a_62185_63363# VDDD sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X5742 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5743 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X5744 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5745 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5746 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5747 VDDD sar10b_0.clknet_1_1__leaf_CLK a_65394_52643# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5748 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5749 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5750 a_68169_66999# a_67209_66999# a_67733_66779# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X5751 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5752 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5753 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5754 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5755 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5756 c1_n1140_52978# m3_n1472_52938# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5757 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5758 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5759 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5760 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5761 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X5762 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5763 a_64594_51052# a_64356_51029# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1648 ps=1.245 w=0.42 l=0.15
X5764 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5765 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5766 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5767 VSSR sar10b_0.SWN[7] a_10731_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5768 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X5769 a_63457_56931# a_63273_56639# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X5770 VDDD a_63797_56924# a_63752_57022# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X5771 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5772 VDDD sar10b_0.net16 a_61677_50190# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X5773 a_61347_52650# a_61086_52650# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X5774 a_68371_62648# a_67393_62635# a_68169_63003# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X5775 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5776 a_60789_51075# sar10b_0.net1 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X5777 a_68379_64392# a_67209_64335# a_68169_64335# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X5778 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5779 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5780 a_63374_62684# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X5781 a_29061_108738# sar10b_0.SWP[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5782 a_2868_111642# sar10b_0.CF[9] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5783 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5784 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5785 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5786 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5787 a_35446_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X5788 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5789 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5790 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5791 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5792 VSSR sar10b_0.SWP[8] a_5929_113881# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5793 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5794 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5795 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5796 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5797 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5798 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5799 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5800 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5801 sar10b_0.SWP[9] a_68946_71059# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5802 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5803 c1_45456_30578# m3_45124_30538# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5804 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5805 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X5806 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5807 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X5808 a_62037_61731# sar10b_0.net2 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X5809 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X5810 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5811 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X5812 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5813 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5814 a_67733_68111# a_67598_68012# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X5815 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y a_6634_8706# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X5816 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5817 a_60690_49683# EN VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.12025 ps=1.065 w=0.74 l=0.15
X5818 c1_n1140_75572# m3_n1472_75532# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5819 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5820 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5821 a_62139_56646# a_60969_56639# a_61929_56639# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X5822 VSSD sar10b_0.net16 a_60780_57975# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5823 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5824 a_63752_57022# a_63273_56639# a_63662_57022# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X5825 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5826 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5827 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5828 a_61609_63602# a_61395_63280# a_60945_63273# VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X5829 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5830 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5831 a_65577_51311# CLK VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5832 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5833 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5834 a_n8277_66083# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS a_n9133_63315# VSSA sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X5835 a_65643_71265# sar10b_0.net43 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X5836 a_66216_52022# a_65861_51977# a_66109_51982# VDDD sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X5837 a_62187_48621# sar10b_0.net30 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X5838 VSSD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X5839 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5840 VSSR sar10b_0.SWP[3] a_29939_111781# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5841 a_63662_57022# a_63273_56639# a_62997_56643# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X5842 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5843 a_20335_112621# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5844 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5845 tdc_0.phase_detector_0.pd_out_0.B tdc_0.phase_detector_0.INN a_53564_60302# VDDA sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X5846 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5847 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5848 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5849 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X5850 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5851 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5852 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5853 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X5854 a_61349_66382# a_61086_65970# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X5855 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5856 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5857 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5858 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5859 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X5860 a_66389_57455# a_66254_57356# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X5861 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5862 VSSR sar10b_0.SWN[3] a_29939_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5863 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5864 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5865 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5866 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5867 a_15533_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5868 c1_31336_21618# m3_31004_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5869 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5870 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5871 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5872 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5873 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5874 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5875 c1_45456_68852# m3_45124_68812# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5876 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5877 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5878 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5879 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5880 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5881 VDDD a_62623_53324# sar10b_0.net6 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X5882 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5883 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5884 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5885 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5886 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X5887 VDDD sar10b_0.net23 a_68946_59303# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X5888 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5889 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5890 a_25137_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5891 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X5892 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5893 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5894 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5895 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5896 VSSD sar10b_0.net16 a_64149_60339# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X5897 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5898 c1_34160_97972# m3_33828_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5899 c1_45456_45138# m3_45124_45098# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5900 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5901 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5902 a_60945_63273# a_61400_63620# a_61349_63718# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X5903 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=3.48 ps=37.92 w=0.5 l=0.5
X5904 VSSD a_60690_54641# sar10b_0.net1 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X5905 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5906 a_63804_67580# a_63663_67678# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.12025 pd=1.065 as=0.35328 ps=1.84 w=0.74 l=0.15
X5907 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5908 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5909 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5910 sar10b_0.clknet_0_CLK a_65577_51311# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1736 ps=1.43 w=1.12 l=0.15
X5911 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5912 VDDD a_63810_50901# sar10b_0.net17 VDDD sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.3304 ps=2.83 w=1.12 l=0.15
X5913 VSSD a_65577_51311# sar10b_0.clknet_0_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X5914 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X5915 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5916 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X5917 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5918 VDDA CLK a_52417_60961# VDDA sky130_fd_pr__pfet_01v8 ad=0.1988 pd=1.505 as=0.147 ps=1.19 w=0.84 l=0.15
X5919 sar10b_0.net4 a_60690_53975# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.74 as=0.0798 ps=0.8 w=0.42 l=0.15
X5920 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5921 sar10b_0.clk_div_0.COUNT\[0\] a_66865_49412# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X5922 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X5923 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5924 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5925 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5926 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X5927 sar10b_0.net29 a_60747_49953# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X5928 a_62997_56643# sar10b_0.net1 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X5929 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5930 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5931 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5932 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5933 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5934 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X5935 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5936 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5937 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5938 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5939 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5940 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5941 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X5942 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5943 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X5944 VDDD a_65577_51311# sar10b_0.clknet_0_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5945 a_61491_52222# sar10b_0.net4 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5946 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5947 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5948 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5949 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X5950 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5951 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5952 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X5953 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X5954 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5955 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X5956 a_67393_63967# a_67209_64335# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X5957 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_111306# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5958 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X5959 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5960 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5961 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5962 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5963 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5964 VDDD sar10b_0.net3 a_66933_65727# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X5965 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5966 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X5967 a_68133_60292# a_67881_60339# a_68271_60396# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X5968 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5969 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5970 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5971 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5972 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5973 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5974 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5975 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5976 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5977 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5978 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5979 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5980 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5981 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5982 VSSD sar10b_0.net16 a_65676_57735# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X5983 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5984 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5985 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5986 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X5987 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5988 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X5989 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5990 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5991 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5992 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5993 a_63475_61316# a_62497_61303# a_63273_61671# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X5994 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5995 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5996 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5997 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X5998 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X5999 tdc_0.OUTN tdc_0.phase_detector_0.pd_out_0.A VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X6000 a_15533_113041# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6001 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6002 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X6003 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[2] a_36482_8700# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X6004 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6005 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X6006 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X6007 a_65577_51311# CLK VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.063 ps=0.72 w=0.42 l=0.15
X6008 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6009 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6010 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6011 VSSR sar10b_0.CF[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X6012 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6013 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6014 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6015 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X6016 sar10b_0._01_ a_64338_52411# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X6017 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6018 c1_n1140_92372# m3_n1472_92332# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6019 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6020 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6021 sar10b_0._12_ a_67564_50907# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2997 ps=2.29 w=0.74 l=0.15
X6022 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X6023 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6024 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6025 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6026 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6027 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6028 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6029 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6030 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6031 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X6032 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6033 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X6034 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6035 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6036 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6037 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6038 VSSA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6039 a_65676_57735# sar10b_0.net1 a_65589_57735# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X6040 a_66919_50029# a_65778_49979# a_66762_50329# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X6041 a_61347_61974# a_61086_61974# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X6042 a_66098_52670# a_65573_52937# a_65928_53032# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.07875 ps=0.865 w=0.42 l=0.15
X6043 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6044 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6045 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6046 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6047 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6048 VDDD a_68169_55011# a_68421_54964# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X6049 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6050 a_62185_50043# a_61395_49960# a_61677_50190# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0735 ps=0.77 w=0.42 l=0.15
X6051 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y a_40248_8706# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X6052 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6053 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6054 VDDD a_62187_71265# sar10b_0.SWP[2] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X6055 VSSD sar10b_0.net4 a_60969_67295# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X6056 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_111306# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6057 c1_n1140_37298# m3_n1472_37258# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6058 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X6059 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6060 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6061 VDDD a_68331_52243# sar10b_0._03_ VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X6062 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6063 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6064 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6065 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X6066 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X6067 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X6068 a_65119_59984# a_64521_60339# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X6069 VSSR sar10b_0.SWN[4] a_25137_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6070 a_63509_62783# a_63374_62684# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X6071 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6072 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X6073 a_61454_53360# a_61249_53311# a_60789_53739# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X6074 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6075 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X6076 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6077 DATA[4] a_68946_56639# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X6078 a_5051_5788# sar10b_0.SWN[8] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6079 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X6080 a_64491_48621# sar10b_0.net32 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X6081 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6082 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6083 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6084 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6085 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6086 VDDR sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X6087 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X6088 VSSR sar10b_0.SWN[7] a_10731_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6089 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6090 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6091 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X6092 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6093 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6094 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6095 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6096 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6097 a_66205_50408# sar10b_0._03_ VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X6098 a_64188_51135# sar10b_0.clknet_1_0__leaf_CLK VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1739 ps=1.21 w=0.74 l=0.15
X6099 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6100 c1_45456_85652# m3_45124_85612# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6101 a_64543_62648# a_63945_63003# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X6102 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y sar10b_0.CF[4] VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X6103 a_61589_50795# a_61454_50696# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X6104 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6105 a_67701_56343# a_67637_56123# a_67623_56343# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X6106 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=1.16 ps=12.64 w=0.5 l=0.5
X6107 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6108 a_64428_50947# a_64199_50761# a_64594_51052# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.0441 ps=0.63 w=0.42 l=0.15
X6109 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6110 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6111 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6112 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6113 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6114 a_65971_66382# a_64993_66255# a_65769_65963# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X6115 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6116 VDDD sar10b_0.cyclic_flag_0.FINAL a_67209_59007# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X6117 VSSR sar10b_0.SWP[8] a_5929_113881# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6118 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6119 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6120 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6121 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6122 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6123 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X6124 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X6125 VSSD a_61041_52340# a_60843_52216# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X6126 a_64492_67433# a_64238_67295# a_64630_67302# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1176 pd=1.4 as=0.0504 ps=0.66 w=0.42 l=0.15
X6127 a_66254_69344# a_66049_69295# a_65589_69723# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X6128 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6129 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6130 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6131 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X6132 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X6133 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6134 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6135 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6136 a_68235_71265# sar10b_0.net45 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X6137 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6138 a_61677_66174# a_61395_65944# a_62038_66346# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X6139 VDDD sar10b_0.net16 a_61086_64638# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X6140 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X6141 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6142 a_68767_54656# a_68169_55011# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X6143 VSSD sar10b_0.net16 a_62901_61671# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X6144 a_66021_66092# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X6145 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6146 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6147 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6148 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6149 a_62261_56123# a_62126_56024# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X6150 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6151 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6152 a_65485_50273# sar10b_0._08_ sar10b_0._02_ VDDD sky130_fd_pr__pfet_01v8 ad=0.1512 pd=1.39 as=0.3304 ps=2.83 w=1.12 l=0.15
X6153 sar10b_0.clknet_0_CLK a_65577_51311# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1792 ps=1.44 w=1.12 l=0.15
X6154 a_67623_56343# a_67297_55975# a_67502_56024# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X6155 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6156 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6157 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6158 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6159 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X6160 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6161 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6162 VDDD sar10b_0.net14 a_65865_69663# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X6163 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X6164 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6165 a_65861_51977# a_65682_51977# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X6166 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X6167 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X6168 a_65385_64631# a_64425_64631# a_64949_64916# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X6169 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X6170 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6171 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6172 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X6173 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6174 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6175 a_62185_62031# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X6176 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6177 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6178 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6179 VDDD sar10b_0.net25 a_68946_63299# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X6180 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6181 a_60747_64231# sar10b_0.net11 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X6182 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6183 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X6184 VDDD sar10b_0.net16 a_60693_56643# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X6185 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6186 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6187 VSSD a_61419_71265# th_dif_sw_0.CK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X6188 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6189 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X6190 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6191 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6192 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6193 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6194 a_5051_113018# sar10b_0.SWP[8] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6195 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6196 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6197 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X6198 a_64533_65967# sar10b_0.net2 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X6199 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6200 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6201 a_66367_66298# a_65769_65963# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X6202 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6203 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6204 a_14655_111306# sar10b_0.SWP[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6205 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6206 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6207 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6208 a_15533_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6209 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X6210 sar10b_0.clknet_0_CLK a_65577_51311# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6211 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6212 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6213 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6214 c1_7332_21618# m3_7000_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6215 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6216 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6217 VDDD a_64888_67630# sar10b_0.cyclic_flag_0.FINAL VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X6218 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6219 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6220 a_14655_5788# sar10b_0.SWN[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6221 VSSR sar10b_0.SWP[4] a_25137_112201# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6222 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6223 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6224 a_25137_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6225 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X6226 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X6227 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X6228 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6229 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6230 c1_38396_97972# m3_38064_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6231 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6232 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6233 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6234 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6235 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A a_35446_111636# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X6236 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6237 a_66049_69295# a_65865_69663# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X6238 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6239 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6240 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X6241 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6242 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X6243 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6244 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X6245 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6246 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6247 VSSD a_66785_50875# sar10b_0.net16 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.04 as=0.1184 ps=1.06 w=0.74 l=0.15
X6248 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6249 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X6250 a_64818_49979# sar10b_0._08_ VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0896 pd=0.92 as=0.0896 ps=0.92 w=0.64 l=0.15
X6251 VSSD sar10b_0.net16 a_62124_61731# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X6252 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6253 VDDD a_65577_51311# sar10b_0.clknet_0_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6254 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6255 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6256 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6257 a_67310_61352# a_67105_61303# a_66645_61731# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X6258 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6259 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6260 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X6261 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6262 a_65390_69010# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X6263 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6264 VSSR sar10b_0.SWP[5] a_20335_112621# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6265 c1_n1140_54098# m3_n1472_54058# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6266 VDDD sar10b_0.net10 a_63849_63299# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X6267 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X6268 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6269 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6270 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A a_1832_111636# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X6271 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X6272 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6273 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6274 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6275 a_29061_108738# sar10b_0.SWP[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6276 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6277 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6278 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6279 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X6280 a_5051_5788# sar10b_0.SWN[8] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6281 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6282 VSSD sar10b_0.net22 a_68946_56639# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X6283 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6284 VDDD a_60747_56239# sar10b_0.CF[0] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X6285 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6286 a_14655_111306# sar10b_0.SWP[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6287 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6288 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6289 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6290 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6291 a_67502_56024# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X6292 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6293 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6294 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6295 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6296 a_65301_57975# sar10b_0.net1 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X6297 a_66666_49313# a_65682_49313# a_66368_49417# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X6298 a_67135_58306# a_66537_57971# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X6299 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X6300 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6301 a_61677_66174# a_61400_66284# a_62007_66027# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X6302 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6303 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6304 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6305 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X6306 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6307 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6308 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6309 VDDD a_65481_59303# a_65733_59432# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X6310 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6311 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_108738# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6312 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6313 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X6314 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X6315 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6316 VSSD a_64188_51135# a_64199_50761# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2553 ps=2.17 w=0.74 l=0.15
X6317 a_62124_61731# sar10b_0.net2 a_62037_61731# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X6318 a_14655_5788# sar10b_0.SWN[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6319 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6320 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6321 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6322 VDDD a_65961_68627# a_66213_68756# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X6323 VSSD a_68479_61316# sar10b_0.net22 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X6324 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6325 a_61419_48621# sar10b_0.net17 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X6326 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6327 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6328 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6329 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6330 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X6331 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X6332 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6333 a_64723_59984# a_63745_59971# a_64521_60339# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X6334 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6335 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6336 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6337 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6338 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6339 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6340 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6341 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6342 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6343 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6344 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X6345 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6346 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6347 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6348 a_68364_51015# sar10b_0.clk_div_0.COUNT\[0\] VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.95 as=0.1961 ps=2.01 w=0.74 l=0.15
X6349 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6350 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6351 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X6352 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6353 VDDD sar10b_0.net11 a_64521_59303# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X6354 c1_45456_47378# m3_45124_47338# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6355 a_68272_51373# sar10b_0.clk_div_0.COUNT\[1\] a_68178_51635# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1312 pd=1.05 as=0.1824 ps=1.85 w=0.64 l=0.15
X6356 VSSD a_62949_56296# a_62907_56400# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X6357 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X6358 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X6359 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6360 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X6361 tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.INP a_53564_59480# VDDA sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.15
X6362 a_61349_63718# a_61086_63306# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X6363 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=2.32 ps=25.28 w=0.5 l=0.5
X6364 a_61609_52946# a_61395_52624# a_60945_52617# VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X6365 a_66312_50368# a_65957_50273# a_66205_50408# VDDD sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X6366 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6367 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6368 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6369 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X6370 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6371 a_29061_108738# sar10b_0.SWP[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6372 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A a_11436_111636# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X6373 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X6374 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6375 VDDD sar10b_0.net12 a_65865_57675# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X6376 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6377 a_66537_57971# a_65577_57971# a_66101_58256# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X6378 sar10b_0.clknet_0_CLK a_65577_51311# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X6379 VSSD sar10b_0.clknet_1_1__leaf_CLK a_65682_51977# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X6380 c1_n1140_22738# m3_n1472_22698# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6381 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X6382 a_61493_58256# a_61358_58354# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X6383 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6384 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6385 VDDD sar10b_0._11_ a_64338_52411# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X6386 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6387 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6388 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6389 VDDD a_61803_48621# sar10b_0.SWN[0] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X6390 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6391 VDDD a_61041_52340# a_60843_52216# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X6392 a_66171_68634# a_65001_68627# a_65961_68627# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X6393 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6394 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6395 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X6396 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6397 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6398 VSSR sar10b_0.SWN[9] a_1127_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6399 VDDD sar10b_0.net12 a_64809_65963# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X6400 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6401 a_62907_56400# a_61737_56343# a_62697_56343# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X6402 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X6403 VSSD a_64339_51661# a_64454_51311# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1155 pd=0.97 as=0.15675 ps=1.67 w=0.55 l=0.15
X6404 VDDD sar10b_0.cyclic_flag_0.FINAL a_67209_63003# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X6405 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6406 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6407 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6408 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6409 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6410 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X6411 a_62007_60699# a_61609_60938# a_61929_60699# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X6412 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X6413 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6414 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6415 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6416 a_25842_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X6417 a_67733_68111# a_67598_68012# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X6418 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6419 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6420 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6421 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6422 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6423 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6424 VSSA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X6425 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6426 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6427 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6428 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6429 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6430 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6431 VSSD sar10b_0.clknet_0_CLK a_66153_48647# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X6432 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6433 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6434 a_7670_8700# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X6435 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6436 a_66213_68756# a_65961_68627# a_66351_68634# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X6437 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X6438 a_64428_50947# a_64188_51135# a_64651_50650# VDDD sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.0504 ps=0.66 w=0.42 l=0.15
X6439 VSSD a_61395_65944# a_61400_66284# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X6440 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X6441 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X6442 VSSA a_n4470_65264# th_dif_sw_0.th_sw_1.CK VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X6443 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6444 c1_28512_97972# m3_28180_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6445 VSSR sar10b_0.SWP[8] a_5929_113881# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6446 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6447 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X6448 a_67881_60339# a_67105_59971# a_67445_60119# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X6449 a_67598_65348# a_67393_65299# a_66933_65727# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X6450 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6451 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X6452 a_64485_56768# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X6453 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X6454 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X6455 a_25137_112201# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6456 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6457 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X6458 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6459 a_62343_57675# a_62017_57307# a_62222_57356# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X6460 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6461 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6462 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6463 a_61395_65944# sar10b_0.net4 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X6464 VSSD sar10b_0.net16 a_61653_53679# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X6465 a_61929_60699# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X6466 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6467 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6468 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6469 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X6470 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6471 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6472 a_65390_69010# a_65001_68627# a_64725_68631# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X6473 VDDD a_61395_64612# a_61400_64952# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X6474 a_64831_56974# a_64233_56639# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X6475 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6476 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6477 a_63295_55988# a_62697_56343# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X6478 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6479 a_68169_65667# a_67393_65299# a_67733_65447# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X6480 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6481 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6482 a_46086_111642# sar10b_0.CF[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X6483 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6484 VDDD a_65525_68912# a_65480_69010# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X6485 a_65185_68919# a_65001_68627# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X6486 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6487 VDDD a_61677_64842# a_61609_64934# VDDD sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X6488 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6489 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X6490 a_68767_62648# a_68169_63003# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X6491 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6492 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6493 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X6494 a_66368_49417# a_66216_49358# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X6495 a_66825_57675# a_66049_57307# a_66389_57455# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X6496 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X6497 a_66049_69295# a_65865_69663# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X6498 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6499 a_20335_112621# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6500 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6501 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X6502 sar10b_0.clknet_0_CLK a_65577_51311# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6503 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X6504 VSSR sar10b_0.SWN[5] a_20335_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6505 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6506 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6507 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6508 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6509 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X6510 c1_5920_21618# m3_5588_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6511 a_61173_64638# a_60945_64605# a_61086_64638# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X6512 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6513 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6514 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6515 a_61653_53679# a_61589_53459# a_61575_53679# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X6516 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6517 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6518 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6519 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6520 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6521 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X6522 VSSR sar10b_0.SWN[3] a_29939_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6523 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6524 VSSD sar10b_0.net16 a_60780_67299# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X6525 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6526 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6527 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6528 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6529 a_15533_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6530 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6531 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X6532 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6533 c1_36984_97972# m3_36652_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6534 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6535 c1_45456_87892# m3_45124_87852# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6536 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6537 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6538 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6539 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6540 VDDD a_65577_51311# sar10b_0.clknet_0_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.1792 pd=1.44 as=0.168 ps=1.42 w=1.12 l=0.15
X6541 VSSD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X6542 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6543 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6544 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X6545 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6546 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6547 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6548 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6549 VSSD sar10b_0.net8 a_63273_56639# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X6550 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6551 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X6552 a_67393_65299# a_67209_65667# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X6553 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6554 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6555 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6556 a_60945_64605# a_61395_64612# a_61347_64638# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X6557 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6558 VDDD sar10b_0.net3 a_65068_49569# VDDD sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.28 as=0.147 ps=1.19 w=0.84 l=0.15
X6559 a_62038_61018# a_61609_60938# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X6560 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6561 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6562 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6563 a_63391_57320# a_62793_57675# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X6564 VSSD a_63871_61316# sar10b_0.net41 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X6565 VSSD a_63621_58960# a_63579_59064# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X6566 a_68421_64288# a_68169_64335# a_68559_64392# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X6567 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6568 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6569 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6570 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6571 VSSA th_dif_sw_0.CKB a_n4470_53722# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6572 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6573 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6574 VDDR sar10b_0.CF[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X6575 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6576 a_61575_53679# a_61249_53311# a_61454_53360# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X6577 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6578 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6579 a_66079_59638# a_65481_59303# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X6580 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6581 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6582 VSSD sar10b_0.net3 a_67020_55071# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X6583 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6584 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6585 a_68371_63980# a_67393_63967# a_68169_64335# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X6586 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6587 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6588 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6589 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X6590 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6591 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X6592 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6593 a_67696_52265# sar10b_0.clk_div_0.COUNT\[2\] VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.147 ps=1.19 w=0.84 l=0.15
X6594 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6595 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6596 VSSR sar10b_0.SWP[5] a_20335_112621# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6597 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6598 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X6599 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6600 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6601 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6602 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6603 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X6604 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6605 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6606 a_64033_63591# a_63849_63299# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X6607 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6608 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6609 a_63797_56924# a_63662_57022# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X6610 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6611 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6612 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6613 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X6614 sar10b_0.net3 a_60690_49683# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X6615 a_22076_111642# sar10b_0.CF[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X6616 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6617 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X6618 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X6619 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6620 a_63579_59064# a_62409_59007# a_63369_59007# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X6621 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6622 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6623 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X6624 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6625 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6626 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6627 a_67733_66779# a_67598_66680# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X6628 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6629 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6630 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6631 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6632 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6633 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6634 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6635 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6636 sar10b_0.net16 a_66785_50875# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1147 ps=1.05 w=0.74 l=0.15
X6637 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6638 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6639 VDDD sar10b_0.net16 a_65589_69723# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X6640 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6641 VDDD sar10b_0.net8 a_62313_61671# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X6642 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6643 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6644 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6645 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6646 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6647 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6648 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6649 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6650 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6651 VSSD sar10b_0.net16 a_60876_51075# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X6652 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X6653 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6654 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6655 VSSR sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X6656 c1_n1140_62132# m3_n1472_62092# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6657 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6658 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6659 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6660 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6661 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6662 VSSD sar10b_0.net16 a_61644_57735# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X6663 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6664 VSSR sar10b_0.SWN[6] a_15533_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6665 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6666 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6667 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6668 c1_45456_32818# m3_45124_32778# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6669 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X6670 a_67881_60339# a_66921_60339# a_67445_60119# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X6671 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X6672 VDDD sar10b_0.net27 a_68946_68627# VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X6673 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X6674 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6675 VSSA th_dif_sw_0.CK a_n4470_65264# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X6676 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6677 a_60747_69559# sar10b_0.net14 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X6678 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 a_9853_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6679 a_66933_55071# sar10b_0.net38 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X6680 a_5929_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6681 a_41284_8700# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X6682 sar10b_0._15_ sar10b_0.clk_div_0.COUNT\[1\] a_68364_51015# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1443 pd=1.13 as=0.0777 ps=0.95 w=0.74 l=0.15
X6683 a_62623_53324# a_62025_53679# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X6684 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6685 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6686 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6687 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6688 c1_n1140_77812# m3_n1472_77772# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6689 a_19457_5788# sar10b_0.SWN[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6690 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6691 a_61677_50190# a_61395_49960# a_62038_50362# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X6692 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6693 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6694 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6695 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6696 VDDD a_63339_71265# sar10b_0.SWP[3] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X6697 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X6698 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6699 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6700 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6701 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X6702 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y a_30644_8706# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X6703 a_65861_49313# a_65682_49313# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X6704 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6705 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6706 a_52417_60961# tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.252 ps=2.28 w=0.84 l=0.15
X6707 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X6708 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6709 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6710 a_60876_51075# sar10b_0.net1 a_60789_51075# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X6711 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X6712 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6713 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X6714 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6715 VDDD sar10b_0.net16 a_62185_52707# VDDD sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X6716 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6717 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6718 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6719 a_66049_57307# a_65865_57675# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X6720 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6721 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X6722 c1_11568_97972# m3_11236_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6723 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6724 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6725 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6726 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6727 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6728 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6729 VDDR sar10b_0.CF[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X6730 VSSA th_dif_sw_0.CKB a_n4470_53722# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6731 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6732 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6733 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6734 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6735 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6736 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 a_5051_113018# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6737 VDDD a_66825_57675# a_67077_57628# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X6738 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6739 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6740 VSSD a_60747_57571# sar10b_0.CF[1] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X6741 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6742 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6743 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X6744 a_67423_69308# a_66825_69663# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X6745 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6746 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6747 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6748 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6749 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6750 VSSR sar10b_0.SWN[7] a_10731_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6751 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A a_26878_111642# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X6752 VDDD a_66389_57455# a_66344_57356# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X6753 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6754 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6755 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6756 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6757 a_66103_50668# a_65586_50645# a_65996_50650# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.07568 pd=0.83 as=0.0588 ps=0.7 w=0.42 l=0.15
X6758 VDDD a_60945_60609# a_60747_60609# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X6759 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6760 a_62527_58306# a_61929_57971# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X6761 a_64373_63584# a_64238_63682# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X6762 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6763 sar10b_0.net10 a_60747_61941# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X6764 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6765 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6766 a_15533_113041# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6767 VDDD a_64085_60119# a_64040_60020# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X6768 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X6769 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X6770 a_64071_60339# a_63745_59971# a_63950_60020# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X6771 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X6772 VDDD sar10b_0.clk_div_0.COUNT\[0\] a_68276_50645# VDDD sky130_fd_pr__pfet_01v8 ad=0.1848 pd=1.45 as=0.308 ps=2.79 w=1.12 l=0.15
X6773 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X6774 a_64620_65967# sar10b_0.net2 a_64533_65967# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X6775 a_68421_62956# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X6776 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X6777 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6778 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6779 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6780 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6781 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6782 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6783 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6784 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6785 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6786 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X6787 DATA[8] a_68946_65963# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X6788 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6789 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6790 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6791 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6792 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6793 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6794 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6795 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6796 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6797 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X6798 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6799 a_24259_5788# sar10b_0.SWN[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6800 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6801 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X6802 a_67611_50645# sar10b_0.clk_div_0.COUNT\[1\] VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3752 pd=2.91 as=0.2352 ps=1.54 w=1.12 l=0.15
X6803 a_68671_55988# a_68073_56343# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X6804 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_108738# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6805 a_65691_59310# a_64521_59303# a_65481_59303# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X6806 a_66732_61731# sar10b_0.net42 a_66645_61731# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X6807 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X6808 VSSD sar10b_0.clk_div_0.COUNT\[3\] a_67372_52833# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.33275 pd=2.31 as=0.17738 ps=1.195 w=0.55 l=0.15
X6809 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X6810 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6811 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6812 a_62593_58639# a_62409_59007# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X6813 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6814 VDDD a_60690_70625# sar10b_0.net2 VDDD sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X6815 a_55121_59650# tdc_0.phase_detector_0.pd_out_0.B a_55085_59917# VDDA sky130_fd_pr__pfet_01v8 ad=0.295 pd=2.59 as=0.135 ps=1.27 w=1 l=0.15
X6816 c1_n1140_24978# m3_n1472_24938# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6817 a_20335_112621# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6818 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6819 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X6820 a_65045_59588# a_64910_59686# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X6821 VSSD sar10b_0.net3 a_67797_68331# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X6822 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6823 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6824 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6825 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6826 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6827 VSSD a_61035_71265# sar10b_0.SWP[1] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X6828 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6829 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X6830 VSSA th_dif_sw_0.CK a_n4470_65264# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6831 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6832 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6833 a_62133_59067# sar10b_0.net1 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X6834 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X6835 VSSD sar10b_0.net16 a_66165_58035# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X6836 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6837 a_61677_50190# a_61400_50300# a_62007_50043# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0504 ps=0.66 w=0.42 l=0.15
X6838 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6839 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6840 VDDD a_66021_66092# a_65971_66382# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X6841 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6842 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6843 VSSR sar10b_0.SWN[7] a_10731_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6844 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6845 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6846 VDDD sar10b_0.net16 a_65589_57735# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X6847 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6848 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6849 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6850 VSSD sar10b_0.net16 a_61173_64638# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X6851 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6852 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6853 a_15533_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6854 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6855 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6856 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X6857 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6858 VDDD sar10b_0.net3 a_66645_61731# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X6859 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6860 VSSD sar10b_0.net3 a_67020_64395# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X6861 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6862 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X6863 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6864 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6865 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6866 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6867 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X6868 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6869 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6870 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6871 VSSR sar10b_0.SWP[4] a_25137_112201# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6872 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6873 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6874 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6875 a_25137_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6876 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6877 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6878 a_61609_60938# a_61400_60956# a_60945_60609# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X6879 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6880 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6881 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6882 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6883 a_65333_66248# a_65198_66346# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X6884 a_67797_68331# a_67733_68111# a_67719_68331# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X6885 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6886 a_29061_108738# sar10b_0.SWP[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6887 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6888 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6889 a_60747_58903# sar10b_0.net7 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X6890 c1_n1140_94612# m3_n1472_94572# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6891 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6892 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6893 a_66165_58035# a_66101_58256# a_66087_58035# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X6894 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X6895 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X6896 a_64705_59595# a_64521_59303# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X6897 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_108738# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6898 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6899 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X6900 VSSD sar10b_0.clknet_1_0__leaf_CLK a_65682_49313# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1739 pd=1.21 as=0.2109 ps=2.05 w=0.74 l=0.15
X6901 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X6902 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X6903 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X6904 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6905 VDDD a_68235_48621# sar10b_0.SWN[7] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X6906 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6907 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6908 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6909 VSSD sar10b_0._10_ a_65299_52305# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1696 pd=1.81 as=0.0672 ps=0.85 w=0.64 l=0.15
X6910 a_64924_52385# sar10b_0._09_ VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.11312 ps=1.065 w=0.55 l=0.15
X6911 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6912 VSSR sar10b_0.SWP[5] a_20335_112621# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6913 a_68384_51373# sar10b_0.clk_div_0.COUNT\[0\] a_68272_51373# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.111 pd=1.045 as=0.1312 ps=1.05 w=0.64 l=0.15
X6914 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6915 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6916 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6917 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6918 sar10b_0.net11 a_60747_63273# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X6919 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6920 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X6921 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6922 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y sar10b_0.CF[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X6923 c1_45456_72212# m3_45124_72172# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6924 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6925 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6926 c1_n1140_39538# m3_n1472_39498# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6927 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6928 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X6929 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6930 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6931 a_67502_56024# a_67113_56343# a_66837_56403# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X6932 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6933 a_61249_50647# a_61065_51015# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X6934 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6935 a_64630_67302# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0777 ps=0.79 w=0.42 l=0.15
X6936 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6937 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6938 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6939 a_67719_68331# a_67393_67963# a_67598_68012# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X6940 a_63745_59971# a_63561_60339# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X6941 a_65966_58354# a_65761_58263# a_65301_57975# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X6942 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6943 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6944 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X6945 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6946 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6947 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6948 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6949 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6950 a_66087_58035# a_65761_58263# a_65966_58354# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X6951 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X6952 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6953 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6954 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X6955 sar10b_0.net2 a_60690_70625# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X6956 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6957 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6958 VDDD a_62025_51015# a_62277_50968# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X6959 a_66933_64395# sar10b_0.net43 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X6960 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6961 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X6962 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6963 a_61035_48621# sar10b_0.net29 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X6964 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6965 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6966 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6967 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6968 VDDD sar10b_0.net16 a_61677_64842# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X6969 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X6970 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X6971 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6972 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6973 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6974 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6975 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6976 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6977 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6978 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6979 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6980 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6981 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6982 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X6983 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X6984 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6985 VDDD a_61589_50795# a_61544_50696# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X6986 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X6987 VSSD a_63391_57320# sar10b_0.net40 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X6988 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6989 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X6990 a_25137_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6991 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X6992 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X6993 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A a_45050_111636# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X6994 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6995 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X6996 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X6997 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6998 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X6999 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7000 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7001 VSSR sar10b_0.SWN[6] a_15533_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7002 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7003 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7004 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X7005 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7006 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7007 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X7008 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7009 VDDD a_66785_50875# a_66700_50645# VDDD sky130_fd_pr__pfet_01v8 ad=0.1302 pd=1.195 as=0.09975 ps=0.895 w=0.42 l=0.15
X7010 VDDD a_60747_65563# sar10b_0.CF[7] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X7011 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7012 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7013 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7014 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7015 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7016 a_61395_49960# sar10b_0.net6 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X7017 a_63525_61624# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X7018 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7019 VDDD sar10b_0.net3 a_66933_55071# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X7020 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7021 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7022 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7023 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7024 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7025 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X7026 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7027 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X7028 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7029 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7030 VSSD a_60747_61567# sar10b_0.CF[4] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X7031 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7032 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7033 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7034 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7035 sar10b_0.clk_div_0.COUNT\[2\] a_66865_52076# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X7036 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7037 c1_n1140_41778# m3_n1472_41738# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7038 VDDD a_66666_51977# a_66865_52076# VDDD sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X7039 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7040 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7041 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7042 a_65011_63718# a_64033_63591# a_64809_63299# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X7043 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7044 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7045 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X7046 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X7047 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X7048 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X7049 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7050 VDDD sar10b_0.net7 a_61833_57675# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X7051 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X7052 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7053 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7054 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X7055 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X7056 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7057 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7058 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7059 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X7060 VSSR sar10b_0.SWN[9] a_1127_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7061 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7062 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7063 c1_21452_21618# m3_21120_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7064 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7065 a_65573_52937# a_65394_52643# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X7066 VSSD a_67371_49579# sar10b_0.SWN[6] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X7067 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7068 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7069 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7070 VDDD a_66789_58100# a_66739_58390# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X7071 VSSD a_64197_62956# a_64155_63060# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X7072 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7073 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7074 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7075 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7076 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7077 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7078 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7079 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7080 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7081 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y sar10b_0.CF[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X7082 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7083 tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.pd_out_0.B a_53652_59132# VSSA sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.15
X7084 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X7085 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7086 VDDD sar10b_0.net16 a_60789_51075# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X7087 VDDD a_68767_66644# sar10b_0.net26 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X7088 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7089 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X7090 VDDD a_64197_62956# a_64147_62648# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X7091 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7092 a_65061_63428# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X7093 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7094 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7095 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7096 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7097 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7098 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7099 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7100 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7101 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X7102 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7103 VSSD sar10b_0.clk_div_0.COUNT\[1\] a_67744_51002# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.12607 pd=1.1 as=0.0888 ps=0.98 w=0.74 l=0.15
X7104 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7105 c1_n1140_64372# m3_n1472_64332# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7106 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7107 VSSD a_62623_53324# sar10b_0.net6 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X7108 a_65355_53949# sar10b_0.clknet_0_CLK VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X7109 a_61493_67580# a_61358_67678# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X7110 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7111 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X7112 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7113 th_dif_sw_0.th_sw_1.CKB a_n4470_53722# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7114 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7115 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[8] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X7116 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7117 a_25137_112201# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7118 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7119 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7120 VSSD sar10b_0.net16 a_63861_56703# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X7121 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7122 a_61249_50647# a_61065_51015# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X7123 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X7124 VDDD sar10b_0.net16 a_62037_61731# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X7125 VDDD a_66027_53575# sar10b_0._05_ VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X7126 VSSD sar10b_0.net16 a_63660_63303# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X7127 a_61086_52650# a_60945_52617# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X7128 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7129 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7130 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7131 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7132 a_66027_53575# sar10b_0._17_ VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X7133 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7134 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7135 VSSD sar10b_0.net10 a_63849_63299# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X7136 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7137 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7138 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7139 sar10b_0._08_ sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X7140 a_64155_63060# a_62985_63003# a_63945_63003# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X7141 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A a_21040_111636# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X7142 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7143 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7144 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7145 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X7146 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7147 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7148 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7149 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7150 VDDD CLK a_65577_51311# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7151 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7152 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7153 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X7154 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7155 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7156 c1_n1140_56338# m3_n1472_56298# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7157 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X7158 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7159 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7160 a_67423_57320# a_66825_57675# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X7161 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7162 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7163 a_62185_63363# sar10b_0.net10 a_62706_63303# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X7164 a_60945_64605# a_61400_64952# a_61349_65050# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.0567 ps=0.69 w=0.42 l=0.15
X7165 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7166 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X7167 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7168 VSSD a_68325_56296# a_68283_56400# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X7169 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7170 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7171 a_20335_112621# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7172 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7173 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7174 VDDR sar10b_0.CF[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X7175 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7176 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7177 a_64197_62956# a_63945_63003# a_64335_63060# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X7178 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7179 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7180 VSSR sar10b_0.SWN[5] a_20335_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7181 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7182 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7183 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7184 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7185 VSSD a_63339_48621# sar10b_0.SWN[3] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X7186 VSSD a_65577_51311# sar10b_0.clknet_0_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X7187 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7188 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7189 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7190 VSSD a_68421_58960# a_68379_59064# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X7191 a_62933_58787# a_62798_58688# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X7192 a_64814_65014# a_64609_64923# a_64149_64635# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X7193 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7194 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7195 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X7196 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7197 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7198 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7199 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7200 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7201 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X7202 VDDD a_60945_65937# a_60747_65937# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X7203 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7204 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7205 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7206 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7207 VSSR sar10b_0.SWN[3] a_29939_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7208 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7209 a_64373_63584# a_64238_63682# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X7210 a_67020_59067# sar10b_0.net39 a_66933_59067# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X7211 a_60747_62899# sar10b_0.net10 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X7212 a_66559_68962# a_65961_68627# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X7213 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X7214 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7215 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7216 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7217 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7218 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X7219 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7220 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7221 VSSR sar10b_0.SWP[8] a_5929_113881# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7222 VDDD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7223 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7224 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7225 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7226 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7227 a_62706_63303# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X7228 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7229 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7230 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7231 a_68283_56400# a_67113_56343# a_68073_56343# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X7232 a_65821_53072# sar10b_0._05_ VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.2972 ps=2.41 w=0.42 l=0.15
X7233 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7234 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X7235 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7236 a_63183_57732# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X7237 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X7238 c1_45456_49618# m3_45124_49578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7239 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X7240 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X7241 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7242 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7243 VSSD a_62527_56974# sar10b_0.net38 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X7244 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7245 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7246 a_68379_59064# a_67209_59007# a_68169_59007# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X7247 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X7248 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7249 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7250 VDDD a_66101_58256# a_66056_58354# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X7251 VSSD a_62527_51646# sar10b_0.net28 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X7252 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7253 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7254 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7255 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7256 VDDD sar10b_0.net16 a_62997_56643# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X7257 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7258 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7259 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7260 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7261 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X7262 a_63950_60020# a_63745_59971# a_63285_60399# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X7263 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7264 a_62222_57356# a_61833_57675# a_61557_57735# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X7265 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X7266 a_64910_59686# a_64521_59303# a_64245_59307# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X7267 a_66869_50413# a_65957_50273# a_66762_50329# VDDD sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X7268 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7269 a_64651_50650# a_64356_51029# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.18985 ps=1.545 w=0.42 l=0.15
X7270 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7271 VSSR sar10b_0.SWP[5] a_20335_112621# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7272 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7273 a_62281_52347# sar10b_0.net6 a_62802_52407# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X7274 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7275 sar10b_0.clknet_0_CLK a_65577_51311# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7276 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7277 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7278 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7279 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7280 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7281 a_67881_61671# a_67105_61303# a_67445_61451# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X7282 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7283 a_67598_66680# a_67393_66631# a_66933_67059# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X7284 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7285 VSSD sar10b_0.net13 a_65001_68627# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X7286 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7287 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X7288 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7289 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7290 a_66795_71265# sar10b_0.net44 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X7291 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X7292 c1_31336_97972# m3_31004_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7293 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7294 VSSD a_67077_69616# a_67035_69720# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X7295 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7296 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7297 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7298 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7299 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7300 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7301 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7302 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7303 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7304 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7305 a_66056_58354# a_65577_57971# a_65966_58354# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X7306 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_111306# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7307 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X7308 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7309 sar10b_0.SWN[9] a_68562_49747# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X7310 c1_17216_21618# m3_16884_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7311 a_62247_56343# a_61921_55975# a_62126_56024# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X7312 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7313 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7314 VDDD sar10b_0.net3 a_66933_64395# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X7315 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X7316 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7317 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7318 VSSD a_66789_58100# a_66747_57978# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X7319 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7320 VSSD a_60690_49683# sar10b_0.net3 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X7321 a_66216_52022# a_65682_51977# a_66109_51982# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.15563 ps=1.215 w=0.42 l=0.15
X7322 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7323 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7324 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7325 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7326 c1_n1140_81172# m3_n1472_81132# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7327 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7328 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7329 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7330 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7331 a_68767_63980# a_68169_64335# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X7332 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X7333 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X7334 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 a_9853_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7335 VDDA tdc_0.OUTP tdc_0.OUTN VDDA sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X7336 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7337 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7338 a_62802_52407# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X7339 c1_45456_51858# m3_45124_51818# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7340 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7341 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7342 a_31680_8700# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X7343 VSSR sar10b_0.SWN[6] a_15533_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7344 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7345 VDDD a_65407_63634# sar10b_0.net43 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X7346 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X7347 a_62007_66027# a_61609_66266# a_61929_66027# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X7348 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7349 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X7350 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7351 a_62415_53736# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X7352 a_64773_60292# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X7353 a_61173_65970# a_60945_65937# a_61086_65970# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X7354 VSSD sar10b_0.cyclic_flag_0.FINAL a_67209_65667# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X7355 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7356 VSSD a_61677_64842# a_61609_64934# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X7357 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X7358 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7359 c1_n1140_96852# m3_n1472_96812# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7360 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7361 c1_n1140_26098# m3_n1472_26058# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7362 a_65068_49569# sar10b_0._07_ VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.1988 ps=1.505 w=0.84 l=0.15
X7363 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7364 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7365 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7366 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7367 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7368 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7369 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7370 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7371 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7372 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_107026# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7373 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7374 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7375 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7376 a_61454_53360# a_61065_53679# a_60789_53739# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X7377 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7378 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7379 a_64491_71265# sar10b_0.net42 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X7380 a_67696_52265# sar10b_0.clk_div_0.COUNT\[2\] VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.1155 ps=0.97 w=0.55 l=0.15
X7381 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X7382 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7383 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7384 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7385 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7386 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7387 a_60945_65937# a_61395_65944# a_61347_65970# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X7388 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7389 a_45050_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X7390 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7391 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7392 c1_45456_74452# m3_45124_74412# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7393 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7394 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7395 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7396 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7397 VDDD sar10b_0.clk_div_0.COUNT\[3\] a_67798_52206# VDDD sky130_fd_pr__pfet_01v8 ad=0.147 pd=1.19 as=0.43785 ps=2.97 w=0.84 l=0.15
X7398 a_62038_62350# a_61609_62270# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.13713 ps=1.155 w=0.42 l=0.15
X7399 a_61929_66027# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X7400 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7401 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7402 a_63810_50901# a_63918_50969# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1862 ps=1.475 w=0.84 l=0.15
X7403 a_61544_53360# a_61065_53679# a_61454_53360# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X7404 VDDD sar10b_0.clknet_0_CLK a_65355_53949# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7405 a_35446_111636# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X7406 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7407 c1_25688_21618# m3_25356_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7408 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X7409 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7410 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X7411 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7412 a_61086_61974# a_60945_61941# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1428 ps=1.225 w=0.42 l=0.15
X7413 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7414 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_111306# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7415 a_61395_64612# sar10b_0.net4 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X7416 VSSD a_60690_49683# sar10b_0.net3 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X7417 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7418 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7419 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7420 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7421 a_66666_51977# a_65682_51977# a_66368_52081# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2331 ps=1.395 w=0.84 l=0.15
X7422 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7423 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7424 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7425 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7426 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7427 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7428 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7429 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7430 a_5051_113018# sar10b_0.SWP[8] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7431 a_63621_58960# a_63369_59007# a_63759_59064# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X7432 a_67393_58639# a_67209_59007# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X7433 VDDD a_65643_48621# sar10b_0.SWN[5] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X7434 a_67252_53653# sar10b_0._16_ VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1376 pd=1.14 as=0.15535 ps=1.17 w=0.64 l=0.15
X7435 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_108738# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7436 sar10b_0._09_ a_64454_51311# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.19013 ps=1.345 w=0.74 l=0.15
X7437 a_1832_111636# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X7438 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7439 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7440 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7441 a_62185_60699# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X7442 VDDA tdc_0.phase_detector_0.pd_out_0.A a_55282_59893# VDDA sky130_fd_pr__pfet_01v8 ad=0.2352 pd=1.54 as=0.3752 ps=2.91 w=1.12 l=0.15
X7443 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X7444 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7445 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7446 a_63571_58652# a_62593_58639# a_63369_59007# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X7447 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7448 a_65573_52937# a_65394_52643# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2553 pd=2.17 as=0.1739 ps=1.21 w=0.74 l=0.15
X7449 a_66344_69344# a_65865_69663# a_66254_69344# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X7450 a_14655_5788# sar10b_0.SWN[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7451 a_24259_5788# sar10b_0.SWN[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7452 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7453 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X7454 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X7455 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X7456 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7457 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7458 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7459 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X7460 VSSD a_68421_68284# a_68379_68388# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X7461 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7462 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7463 a_62185_66027# a_61400_66284# a_61677_66174# VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X7464 VDDD a_66367_66298# sar10b_0.net45 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X7465 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7466 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7467 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7468 VSSD a_68421_62956# a_68379_63060# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X7469 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7470 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X7471 VDDD a_65769_65963# a_66021_66092# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X7472 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7473 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7474 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7475 VSSD a_68767_67976# sar10b_0.net27 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X7476 tdc_0.OUTN tdc_0.OUTP a_54660_59599# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X7477 VDDD a_65577_51311# sar10b_0.clknet_0_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X7478 VSSD a_62187_71265# sar10b_0.SWP[2] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X7479 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X7480 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X7481 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X7482 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7483 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7484 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7485 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7486 VDDD a_68421_62956# a_68371_62648# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X7487 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7488 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7489 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7490 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7491 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7492 a_67020_63063# sar10b_0.net44 a_66933_63063# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X7493 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X7494 a_20335_112621# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7495 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7496 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X7497 a_67598_65348# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X7498 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7499 c1_45456_89012# m3_45124_88972# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7500 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X7501 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7502 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7503 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X7504 VDDD sar10b_0.net9 a_62185_62031# VDDD sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X7505 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7506 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7507 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7508 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_111306# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7509 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7510 a_66378_52993# a_65573_52937# a_66080_53027# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X7511 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X7512 VSSD sar10b_0.net16 a_61548_56403# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X7513 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A a_36482_111642# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X7514 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7515 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7516 a_68169_65667# a_67209_65667# a_67733_65447# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X7517 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7518 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X7519 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X7520 a_68379_68388# a_67209_68331# a_68169_68331# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X7521 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7522 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X7523 VDDD sar10b_0.net16 a_64533_65967# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X7524 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7525 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7526 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X7527 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7528 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X7529 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7530 a_5051_5788# sar10b_0.SWN[8] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7531 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7532 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7533 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7534 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7535 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7536 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7537 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7538 a_15533_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7539 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7540 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7541 a_68379_63060# a_67209_63003# a_68169_63003# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X7542 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7543 a_14655_111306# sar10b_0.SWP[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7544 a_66367_66298# a_65769_65963# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X7545 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X7546 VSSD a_60945_65937# a_60747_65937# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X7547 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7548 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X7549 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7550 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X7551 a_11436_111636# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X7552 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7553 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7554 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7555 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7556 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7557 VSSR sar10b_0.SWP[4] a_25137_112201# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7558 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7559 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7560 a_24259_5788# sar10b_0.SWN[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7561 a_64147_62648# a_63169_62635# a_63945_63003# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X7562 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X7563 a_64623_56646# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X7564 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7565 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7566 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7567 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7568 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X7569 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7570 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X7571 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7572 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7573 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7574 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X7575 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7576 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X7577 a_63045_57628# a_62793_57675# a_63183_57732# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X7578 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7579 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7580 sar10b_0.net16 a_66785_50875# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.111 ps=1.04 w=0.74 l=0.15
X7581 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7582 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7583 VSSD sar10b_0.net16 a_60780_56643# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X7584 sar10b_0.net4 a_60690_53975# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X7585 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X7586 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7587 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7588 th_dif_sw_0.VCP th_dif_sw_0.th_sw_1.th_sw_main_0.VGS VINP VSSA sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=5.8 ps=40.58 w=20 l=0.15
X7589 a_67400_61352# a_66921_61671# a_67310_61352# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X7590 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7591 a_65928_53032# a_65573_52937# a_65821_53072# VDDD sky130_fd_pr__pfet_01v8 ad=0.09835 pd=1.005 as=0.09835 ps=1.005 w=0.42 l=0.15
X7592 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7593 VSSD sar10b_0.net16 a_63084_67299# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X7594 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y sar10b_0.CF[3] VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X7595 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7596 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7597 a_64040_60020# a_63561_60339# a_63950_60020# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X7598 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X7599 c1_4508_21618# m3_4176_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7600 VSSD a_61677_50190# a_61609_50282# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X7601 a_38665_107026# sar10b_0.SWP[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7602 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7603 c1_45456_91252# m3_45124_91212# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7604 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X7605 a_62527_51646# a_61929_51311# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X7606 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X7607 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7608 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7609 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7610 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7611 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7612 a_68421_64288# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X7613 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7614 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7615 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7616 c1_15804_21618# m3_15472_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7617 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7618 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7619 a_61131_70891# sar10b_0.net38 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X7620 VDDD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7621 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7622 a_61419_71265# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X7623 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7624 VDDD sar10b_0.net16 a_65301_57975# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X7625 a_66368_52081# a_66216_52022# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.18985 ps=1.545 w=0.84 l=0.15
X7626 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X7627 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X7628 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7629 a_61349_65050# a_61086_64638# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.08925 ps=0.845 w=0.42 l=0.15
X7630 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X7631 VSSD a_67372_52243# sar10b_0._07_ VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.14887 pd=1.195 as=0.2109 ps=2.05 w=0.74 l=0.15
X7632 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7633 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7634 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7635 c1_7332_97972# m3_7000_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7636 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7637 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7638 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X7639 VSSR sar10b_0.CF[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X7640 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X7641 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7642 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7643 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X7644 c1_41220_21618# m3_40888_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7645 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7646 a_64725_68631# sar10b_0.net2 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X7647 a_15533_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7648 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7649 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7650 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7651 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7652 c1_45456_36178# m3_45124_36138# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7653 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7654 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7655 DATA[1] a_68946_49747# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X7656 a_5051_113018# sar10b_0.SWP[8] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7657 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X7658 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7659 a_66700_50645# a_65765_50645# a_66593_50645# VDDD sky130_fd_pr__pfet_01v8 ad=0.09975 pd=0.895 as=0.1428 ps=1.225 w=0.42 l=0.15
X7660 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7661 a_14655_111306# sar10b_0.SWP[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7662 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7663 a_62235_53736# a_61065_53679# a_62025_53679# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X7664 a_29061_108738# sar10b_0.SWP[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7665 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7666 a_63084_67299# sar10b_0.net14 a_62997_67299# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X7667 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7668 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A a_12472_111642# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X7669 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7670 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7671 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7672 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_110450# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7673 a_33863_5788# sar10b_0.SWN[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7674 VSSR sar10b_0.SWN[6] a_15533_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7675 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7676 a_61395_49960# sar10b_0.net6 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X7677 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7678 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X7679 VSSD sar10b_0.net3 a_67797_66999# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X7680 a_64705_59595# a_64521_59303# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X7681 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X7682 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7683 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7684 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7685 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X7686 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X7687 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X7688 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7689 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7690 VDDD a_62277_53632# a_62227_53324# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X7691 a_66464_50363# a_66312_50368# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.10905 pd=1.025 as=0.1648 ps=1.245 w=0.55 l=0.15
X7692 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7693 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7694 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7695 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X7696 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7697 a_62277_53632# a_62025_53679# a_62415_53736# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X7698 VSSD sar10b_0.net16 a_61173_65970# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X7699 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7700 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7701 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7702 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7703 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7704 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X7705 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7706 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7707 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7708 tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A a_51345_58977# a_51861_59345# VDDA sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=1
X7709 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X7710 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X7711 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X7712 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7713 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7714 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X7715 a_62185_52707# sar10b_0.net16 a_62706_52647# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X7716 VSSD sar10b_0.net11 a_64521_59303# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X7717 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7718 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X7719 VDDD a_62181_67424# a_62131_67714# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X7720 VDDD a_61493_58256# a_61448_58354# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X7721 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7722 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7723 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7724 VDDD a_67733_65447# a_67688_65348# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X7725 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7726 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7727 VSSR sar10b_0.SWP[3] a_29939_111781# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7728 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X7729 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7730 a_64356_51029# a_64188_51135# a_63918_50969# VDDD sky130_fd_pr__pfet_01v8 ad=0.2331 pd=1.395 as=0.1428 ps=1.225 w=0.84 l=0.15
X7731 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7732 VDDD sar10b_0.net16 a_61773_52237# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.1239 ps=1.43 w=0.42 l=0.15
X7733 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7734 VDDD a_63525_61624# a_63475_61316# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X7735 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7736 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7737 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7738 a_67797_66999# a_67733_66779# a_67719_66999# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X7739 th_dif_sw_0.VCN VCM sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7740 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7741 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7742 a_64993_66255# a_64809_65963# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X7743 a_63662_57022# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X7744 a_67105_59971# a_66921_60339# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X7745 a_67393_62635# a_67209_63003# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X7746 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A a_40248_111636# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X7747 VSSD sar10b_0.net16 a_62220_59067# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X7748 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7749 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7750 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7751 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7752 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7753 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7754 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7755 VDDD a_67077_69616# a_67027_69308# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X7756 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X7757 a_14655_111306# sar10b_0.SWP[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7758 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7759 VSSD sar10b_0._12_ a_67526_50041# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1376 ps=1.14 w=0.64 l=0.15
X7760 VSSD sar10b_0.net10 a_63561_60339# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X7761 a_67598_68012# a_67209_68331# a_66933_68391# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X7762 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7763 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7764 VSSD sar10b_0.net16 a_65589_68691# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X7765 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7766 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7767 a_16238_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X7768 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7769 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7770 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7771 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X7772 VSSD tdc_0.OUTP a_60690_70625# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X7773 a_62706_52647# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X7774 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X7775 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7776 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7777 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X7778 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7779 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X7780 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7781 DATA[4] a_68946_56639# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.119 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X7782 a_65045_59588# a_64910_59686# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X7783 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X7784 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7785 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7786 a_67688_65348# a_67209_65667# a_67598_65348# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X7787 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.2331 ps=2.11 w=0.74 l=0.15
X7788 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7789 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7790 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7791 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7792 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7793 a_25137_112201# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7794 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7795 sar10b_0.clk_div_0.COUNT\[1\] a_66961_50219# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1229 ps=1.085 w=0.74 l=0.15
X7796 a_67719_66999# a_67393_66631# a_67598_66680# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0735 ps=0.77 w=0.42 l=0.15
X7797 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7798 VSSD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X7799 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7800 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7801 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X7802 a_67733_58787# a_67598_58688# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X7803 VSSD a_66865_52076# a_66823_52361# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05565 ps=0.685 w=0.42 l=0.15
X7804 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7805 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7806 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7807 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7808 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7809 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7810 a_61395_64612# sar10b_0.net4 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X7811 VDDD a_65061_63428# a_65011_63718# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X7812 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7813 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X7814 a_65928_53032# a_65394_52643# a_65821_53072# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.07875 pd=0.865 as=0.15563 ps=1.215 w=0.42 l=0.15
X7815 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7816 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X7817 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7818 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7819 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7820 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X7821 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X7822 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7823 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7824 a_65589_68691# a_65525_68912# a_65511_68691# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X7825 VDDD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7826 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X7827 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7828 a_64085_60119# a_63950_60020# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X7829 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7830 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7831 a_61347_60642# a_61086_60642# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0756 ps=0.78 w=0.42 l=0.15
X7832 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X7833 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7834 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X7835 VSSD a_65983_64966# sar10b_0.net44 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X7836 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7837 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7838 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X7839 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7840 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X7841 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7842 a_62623_50660# a_62025_51015# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X7843 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7844 th_dif_sw_0.VCP VCM sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7845 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7846 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7847 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7848 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7849 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X7850 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7851 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7852 VSSD a_63295_55988# sar10b_0.net39 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X7853 VINP th_dif_sw_0.th_sw_1.CK VINP VSSA sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=18.56 ps=130.32001 w=20 l=0.15
X7854 VDDD a_65577_51311# sar10b_0.clknet_0_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7855 a_24259_5788# sar10b_0.SWN[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7856 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7857 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7858 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7859 VSSR sar10b_0.SWN[5] a_20335_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7860 c1_45456_76692# m3_45124_76652# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7861 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7862 a_68091_61728# a_66921_61671# a_67881_61671# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X7863 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X7864 DATA[0] a_68562_48647# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X7865 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7866 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7867 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7868 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7869 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7870 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7871 a_64443_56646# a_63273_56639# a_64233_56639# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.229 ps=1.64 w=0.42 l=0.15
X7872 VSSR sar10b_0.SWN[3] a_29939_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7873 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7874 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7875 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X7876 sar10b_0.clknet_0_CLK a_65577_51311# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X7877 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7878 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7879 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7880 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7881 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7882 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7883 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7884 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7885 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_110450# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7886 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7887 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7888 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7889 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7890 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7891 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7892 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7893 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7894 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7895 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X7896 VDDD sar10b_0.clk_div_0.COUNT\[0\] a_65485_50273# VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1512 ps=1.39 w=1.12 l=0.15
X7897 VDDD sar10b_0.net8 a_63273_56639# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X7898 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1792 ps=1.44 w=1.12 l=0.15
X7899 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7900 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X7901 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7902 a_62007_50043# a_61609_50282# a_61929_50043# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.0504 ps=0.66 w=0.42 l=0.15
X7903 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7904 a_19457_110450# sar10b_0.SWP[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7905 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7906 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7907 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7908 a_64485_56768# a_64233_56639# a_64623_56646# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X7909 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7910 a_65525_68912# a_65390_69010# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X7911 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7912 VSSD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X7913 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7914 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7915 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X7916 VDDD sar10b_0.clknet_1_0__leaf_CLK a_65682_49313# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7917 a_67881_61671# a_66921_61671# a_67445_61451# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X7918 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7919 a_61677_64842# a_61395_64612# a_62038_65014# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X7920 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7921 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7922 VSSD sar10b_0.net7 a_61065_51015# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X7923 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7924 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7925 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7926 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7927 VDDD a_68767_67976# sar10b_0.net27 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X7928 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7929 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7930 a_26878_111642# sar10b_0.CF[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X7931 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7932 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7933 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7934 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7935 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7936 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7937 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7938 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X7939 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7940 c1_5920_97972# m3_5588_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7941 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7942 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7943 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7944 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7945 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7946 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7947 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7948 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7949 a_61929_50043# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.21123 ps=1.45 w=0.42 l=0.15
X7950 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X7951 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X7952 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7953 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7954 a_60747_62899# sar10b_0.net10 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X7955 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X7956 VDDD a_63391_57320# sar10b_0.net40 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X7957 a_68169_55011# a_67393_54643# a_67733_54791# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X7958 a_29061_5788# sar10b_0.SWN[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7959 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X7960 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7961 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7962 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7963 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7964 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7965 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7966 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7967 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7968 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7969 c1_45456_21618# m3_45124_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7970 a_62497_61303# a_62313_61671# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X7971 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X7972 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7973 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X7974 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7975 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7976 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 a_5051_113018# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7977 VSSD a_67798_52206# a_67372_52243# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.165 pd=1.7 as=0.09212 ps=0.885 w=0.55 l=0.15
X7978 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7979 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7980 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7981 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7982 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X7983 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7984 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7985 a_25137_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7986 sar10b_0.net5 a_60747_52617# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X7987 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X7988 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[6] a_17274_8700# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X7989 c1_n1140_66612# m3_n1472_66572# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7990 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X7991 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7992 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7993 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7994 a_67651_51991# sar10b_0.clk_div_0.COUNT\[0\] a_67543_51991# VDDD sky130_fd_pr__pfet_01v8 ad=0.165 pd=1.33 as=0.195 ps=1.39 w=1 l=0.15
X7995 VSSR sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X7996 VDDD a_61493_67580# a_61448_67678# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X7997 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X7998 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X7999 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X8000 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X8001 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8002 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X8003 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8004 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8005 VSSD a_60747_58903# sar10b_0.CF[2] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X8006 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X8007 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8008 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X8009 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8010 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8011 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8012 VSSD sar10b_0.net14 a_65865_69663# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2109 ps=2.05 w=0.74 l=0.15
X8013 a_62185_50043# a_61400_50300# a_61677_50190# VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.063 ps=0.72 w=0.42 l=0.15
X8014 a_53564_60302# tdc_0.phase_detector_0.INP VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X8015 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8016 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8017 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X8018 a_64332_59307# sar10b_0.net1 a_64245_59307# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X8019 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8020 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8021 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X8022 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X8023 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8024 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8025 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8026 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8027 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X8028 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8029 a_67310_60020# a_67105_59971# a_66645_60399# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X8030 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8031 VSSR sar10b_0.SWP[5] a_20335_112621# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8032 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8033 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 a_14655_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8034 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8035 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8036 a_10731_113461# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8037 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8038 a_67393_54643# a_67209_55011# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X8039 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8040 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8041 a_68421_58960# a_68169_59007# a_68559_59064# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X8042 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8043 VDDD a_60747_60235# sar10b_0.CF[3] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X8044 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8045 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8046 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X8047 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8048 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8049 VSSR sar10b_0.SWP[3] a_29939_111781# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8050 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8051 c1_45456_93492# m3_45124_93452# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8052 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X8053 VDDD a_64773_60292# a_64723_59984# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X8054 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8055 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X8056 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8057 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8058 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8059 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8060 VSSD sar10b_0.net18 a_68562_48647# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.1197 ps=1.41 w=0.42 l=0.15
X8061 a_68169_55011# a_67209_55011# a_67733_54791# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X8062 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8063 a_68371_58652# a_67393_58639# a_68169_59007# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X8064 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8065 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8066 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8067 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8068 VSSD a_62527_58306# sar10b_0.net8 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X8069 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8070 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8071 VSSR sar10b_0.SWN[0] a_44345_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8072 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8073 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X8074 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8075 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X8076 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8077 a_63087_56400# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X8078 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8079 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X8080 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8081 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8082 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8083 a_66389_69443# a_66254_69344# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X8084 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8085 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8086 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8087 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8088 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8089 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8090 a_66732_60399# sar10b_0.net41 a_66645_60399# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X8091 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8092 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8093 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X8094 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X8095 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X8096 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8097 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X8098 a_62126_56024# a_61737_56343# a_61461_56403# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X8099 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8100 a_19457_110450# sar10b_0.SWP[5] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8101 a_14655_5788# sar10b_0.SWN[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8102 VSSD sar10b_0.net4 a_63273_67295# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.2109 ps=2.05 w=0.74 l=0.15
X8103 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8104 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8105 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X8106 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X8107 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8108 VDDD a_68169_63003# a_68421_62956# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X8109 a_66103_50668# a_65765_50645# a_65996_50650# VDDD sky130_fd_pr__pfet_01v8 ad=0.08873 pd=0.895 as=0.08873 ps=0.895 w=0.42 l=0.15
X8110 a_61041_52340# a_61491_52222# a_61443_52404# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X8111 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X8112 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8113 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X8114 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8115 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8116 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8117 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8118 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8119 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8120 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8121 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X8122 VSSD a_69003_71265# sar10b_0.SWP[8] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X8123 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8124 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8125 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8126 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8127 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8128 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X8129 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8130 VDDD a_66378_52993# a_66577_52883# VDDD sky130_fd_pr__pfet_01v8 ad=0.1862 pd=1.475 as=0.2478 ps=2.27 w=0.84 l=0.15
X8131 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8132 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X8133 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X8134 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8135 a_62227_53324# a_61249_53311# a_62025_53679# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X8136 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X8137 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X8138 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8139 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8140 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8141 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X8142 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8143 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8144 VSSA a_n4470_53722# th_dif_sw_0.th_sw_1.CKB VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8145 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8146 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X8147 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8148 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8149 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X8150 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8151 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8152 a_45050_111636# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X8153 VSSD sar10b_0.net16 a_64812_68631# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X8154 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8155 a_29061_5788# sar10b_0.SWN[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8156 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8157 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X8158 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X8159 VDDD sar10b_0.net16 a_62133_59067# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X8160 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8161 VSSD a_61803_48621# sar10b_0.SWN[0] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X8162 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8163 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8164 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8165 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8166 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8167 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8168 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8169 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8170 a_64146_51029# a_63810_50901# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1197 ps=1.41 w=0.42 l=0.15
X8171 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8172 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8173 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8174 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 a_5051_113018# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8175 a_63967_58652# a_63369_59007# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X8176 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X8177 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8178 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8179 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8180 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X8181 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_108738# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8182 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8183 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8184 a_14655_5788# sar10b_0.SWN[6] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8185 VSSD a_66961_50219# a_66919_50029# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.05565 ps=0.685 w=0.42 l=0.15
X8186 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8187 VDDD sar10b_0.net9 a_62985_63003# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X8188 c1_n1140_83412# m3_n1472_83372# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8189 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8190 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X8191 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS a_n9133_57045# w_n9655_56533# w_n9655_56533# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
X8192 th_dif_sw_0.VCN th_dif_sw_0.th_sw_1.CK th_dif_sw_0.VCN VSSA sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=17.4 ps=121.74 w=20 l=0.15
X8193 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X8194 a_66762_50329# a_65957_50273# a_66464_50363# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1181 pd=1.035 as=0.10905 ps=1.025 w=0.55 l=0.15
X8195 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8196 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8197 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X8198 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X8199 VSSR sar10b_0.SWP[4] a_25137_112201# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8200 VSSD a_61395_64612# a_61400_64952# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X8201 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X8202 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8203 a_67598_64016# a_67393_63967# a_66933_64395# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X8204 a_64812_68631# sar10b_0.net2 a_64725_68631# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X8205 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8206 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X8207 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8208 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8209 VSSD a_65068_49569# sar10b_0._10_ VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.2109 ps=2.05 w=0.74 l=0.15
X8210 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8211 VDDD a_68235_71265# sar10b_0.SWP[7] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X8212 VSSD sar10b_0.net3 a_67701_56343# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X8213 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8214 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8215 VSSD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8216 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8217 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8218 a_61705_51992# a_61496_52091# a_61041_52340# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.229 ps=1.64 w=0.74 l=0.15
X8219 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8220 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8221 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8222 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8223 a_62185_50043# sar10b_0.net1 a_62706_49983# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X8224 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X8225 c1_n1140_28338# m3_n1472_28298# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8226 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8227 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8228 VINN th_dif_sw_0.th_sw_0.th_sw_main_0.VGS a_n8277_54249# VSSA sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X8229 a_68169_64335# a_67393_63967# a_67733_64115# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X8230 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8231 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8232 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8233 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8234 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8235 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8236 a_29061_108738# sar10b_0.SWP[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8237 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8238 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8239 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0735 ps=0.77 w=0.42 l=0.15
X8240 a_69003_48621# sar10b_0.net36 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X8241 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8242 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X8243 VDDD a_62181_51440# a_62131_51730# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X8244 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8245 a_20335_112621# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8246 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X8247 VDDD a_63295_55988# sar10b_0.net39 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X8248 a_61035_71265# sar10b_0.net39 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X8249 sar10b_0.net10 a_60747_61941# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X8250 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8251 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8252 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8253 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8254 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8255 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8256 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X8257 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8258 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8259 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8260 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8261 a_68671_55988# a_68073_56343# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X8262 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X8263 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8264 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8265 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8266 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8267 VSSR sar10b_0.SWN[4] a_25137_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8268 a_61173_63306# a_60945_63273# a_61086_63306# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.1197 ps=1.41 w=0.42 l=0.15
X8269 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8270 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8271 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8272 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8273 VSSD a_60747_68227# sar10b_0.CF[8] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X8274 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X8275 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8276 VSSD a_64831_56974# sar10b_0.net31 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X8277 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8278 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X8279 a_62706_49983# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X8280 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8281 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8282 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8283 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8284 a_21040_111636# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X8285 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8286 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8287 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8288 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X8289 VSSD a_68767_66644# sar10b_0.net26 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X8290 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8291 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8292 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8293 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8294 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X8295 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8296 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8297 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8298 VDDD a_68421_64288# a_68371_63980# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X8299 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8300 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8301 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8302 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X8303 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8304 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8305 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8306 a_67393_63967# a_67209_64335# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X8307 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X8308 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8309 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8310 VSSR sar10b_0.SWN[6] a_15533_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8311 a_60945_63273# a_61395_63280# a_61347_63306# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.0504 ps=0.66 w=0.42 l=0.15
X8312 a_65525_68912# a_65390_69010# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X8313 VDDD a_61929_67295# a_62181_67424# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X8314 a_67598_66680# sar10b_0.net3 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.1239 pd=1.43 as=0.13713 ps=1.155 w=0.42 l=0.15
X8315 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8316 a_68421_68284# a_68169_68331# a_68559_68388# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X8317 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8318 VDDA th_dif_sw_0.th_sw_1.th_sw_main_0.VGS w_n9655_63119# w_n9655_63119# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.15
X8319 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8320 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8321 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8322 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8323 a_62709_63063# sar10b_0.net2 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X8324 a_68421_62956# a_68169_63003# a_68559_63060# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X8325 c1_n1140_30578# m3_n1472_30538# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8326 VDDD a_60747_64231# sar10b_0.CF[6] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X8327 VDDD a_63273_61671# a_63525_61624# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X8328 VSSD sar10b_0.net3 a_67020_59067# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X8329 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8330 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X8331 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X8332 VSSD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8333 sar10b_0.clknet_1_1__leaf_CLK a_65355_53949# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.1792 ps=1.44 w=1.12 l=0.15
X8334 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8335 a_68371_67976# a_67393_67963# a_68169_68331# VDDD sky130_fd_pr__pfet_01v8 ad=0.0567 pd=0.69 as=0.23015 ps=1.73 w=0.42 l=0.15
X8336 a_29061_108738# sar10b_0.SWP[3] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8337 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8338 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8339 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8340 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8341 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8342 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X8343 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8344 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8345 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8346 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8347 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8348 a_2868_8700# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X8349 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8350 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X8351 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8352 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8353 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X8354 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8355 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8356 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X8357 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8358 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8359 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8360 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8361 a_61131_70891# sar10b_0.net38 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X8362 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8363 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8364 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8365 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8366 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X8367 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8368 a_63797_56924# a_63662_57022# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X8369 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8370 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8371 VSSR sar10b_0.SWP[3] a_29939_111781# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8372 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8373 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8374 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8375 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X8376 a_62017_57307# a_61833_57675# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X8377 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8378 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8379 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8380 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8381 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8382 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8383 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8384 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8385 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X8386 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X8387 a_67733_65447# a_67598_65348# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.24605 pd=1.405 as=0.21123 ps=1.45 w=0.74 l=0.15
X8388 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8389 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X8390 a_43467_106170# sar10b_0.SWP[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8391 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8392 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8393 VSSR sar10b_0.SWP[1] a_39543_110941# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8394 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 a_33863_107882# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8395 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8396 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8397 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8398 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8399 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8400 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8401 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.1036 ps=1.02 w=0.74 l=0.15
X8402 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8403 c1_45456_23858# m3_45124_23818# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8404 a_68559_64392# sar10b_0.net3 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0441 pd=0.63 as=0.0756 ps=0.78 w=0.42 l=0.15
X8405 VSSD sar10b_0.net16 a_61269_52404# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X8406 a_62949_56296# a_62697_56343# a_63087_56400# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0441 ps=0.63 w=0.42 l=0.15
X8407 a_61609_60938# a_61395_60616# a_60945_60609# VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X8408 VDDD a_64809_63299# a_65061_63428# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X8409 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8410 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X8411 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X8412 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8413 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X8414 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8415 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8416 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8417 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A a_25842_111636# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X8418 VSSR sar10b_0.SWN[6] a_15533_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8419 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8420 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8421 c1_n1140_68852# m3_n1472_68812# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8422 VSSR sar10b_0.SWP[2] a_34741_111361# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8423 a_66933_59067# sar10b_0.net39 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X8424 a_61419_71265# sar10b_0.net16 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.1638 ps=1.2 w=0.42 l=0.15
X8425 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X8426 a_66254_57356# a_66049_57307# a_65589_57735# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X8427 a_25137_112201# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8428 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8429 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8430 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8431 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8432 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8433 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8434 VDDD a_64949_64916# a_64904_65014# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X8435 a_63810_50901# a_63918_50969# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1824 pd=1.85 as=0.1229 ps=1.085 w=0.64 l=0.15
X8436 VDDD sar10b_0.net16 a_61086_52650# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X8437 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8438 c1_n1140_45138# m3_n1472_45098# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8439 a_60747_69559# sar10b_0.net14 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X8440 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X8441 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1184 ps=1.06 w=0.74 l=0.15
X8442 VDDD a_62949_56296# a_62899_55988# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X8443 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8444 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X8445 a_n8277_65767# th_dif_sw_0.th_sw_1.CK VSSA VSSA sky130_fd_pr__nfet_01v8 ad=2.175 pd=15.58 as=2.175 ps=15.58 w=7.5 l=0.15
X8446 VSSD a_61395_49960# a_61400_50300# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1295 pd=1.09 as=0.2627 ps=2.19 w=0.74 l=0.15
X8447 VDDD sar10b_0._07_ sar10b_0._08_ VDDD sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X8448 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X8449 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8450 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8451 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X8452 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8453 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X8454 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X8455 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2331 pd=2.11 as=0.1184 ps=1.06 w=0.74 l=0.15
X8456 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8457 VDDD a_66559_68962# sar10b_0.net46 VDDD sky130_fd_pr__pfet_01v8 ad=0.336 pd=2.84 as=0.3808 ps=2.92 w=1.12 l=0.15
X8458 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8459 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8460 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8461 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8462 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8463 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X8464 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8465 a_63621_58960# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X8466 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8467 a_65577_51311# CLK VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8468 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8469 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8470 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8471 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X8472 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X8473 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8474 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8475 c1_21452_97972# m3_21120_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8476 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8477 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X8478 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8479 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8480 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8481 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1184 pd=1.06 as=0.1221 ps=1.07 w=0.74 l=0.15
X8482 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8483 a_62185_50043# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1176 ps=1.4 w=0.42 l=0.15
X8484 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8485 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 a_249_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8486 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8487 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8488 VSSD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X8489 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8490 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8491 VSSR sar10b_0.SWN[5] a_20335_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8492 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X8493 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1295 ps=1.09 w=0.74 l=0.15
X8494 a_64904_65014# a_64425_64631# a_64814_65014# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X8495 a_43467_5788# sar10b_0.SWN[0] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8496 sar10b_0._00_ a_65021_50292# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X8497 a_39543_110941# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8498 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8499 a_66153_48647# sar10b_0.clknet_0_CLK VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.1197 ps=1.41 w=0.42 l=0.15
X8500 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8501 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 a_19457_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8502 VSSD a_60747_56239# sar10b_0.CF[0] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X8503 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8504 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8505 c1_39808_21618# m3_39476_21578# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8506 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8507 a_65355_53949# sar10b_0.clknet_0_CLK VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.063 ps=0.72 w=0.42 l=0.15
X8508 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8509 VSSR sar10b_0.SWN[3] a_29939_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8510 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8511 VDDD a_60945_64605# a_60747_64605# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.2478 ps=2.27 w=0.84 l=0.15
X8512 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8513 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X8514 sar10b_0.net13 a_60747_65937# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3808 pd=2.92 as=0.336 ps=2.84 w=1.12 l=0.15
X8515 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8516 c1_45456_38418# m3_45124_38378# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8517 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8518 VSSD a_66213_68756# a_66171_68634# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0504 ps=0.66 w=0.42 l=0.15
X8519 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8520 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8521 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8522 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8523 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X8524 a_65821_53072# sar10b_0._05_ VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15563 pd=1.215 as=0.23015 ps=2.1 w=0.42 l=0.15
X8525 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8526 a_53564_59480# tdc_0.phase_detector_0.INN VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.15
X8527 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8528 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8529 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8530 a_61705_51992# a_61491_52222# a_61041_52340# VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.23015 ps=1.73 w=1 l=0.15
X8531 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X8532 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8533 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8534 VSSD sar10b_0._00_ a_64761_51028# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.23015 pd=2.1 as=0.15563 ps=1.215 w=0.42 l=0.15
X8535 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X8536 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8537 VDDD a_67733_66779# a_67688_66680# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X8538 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8539 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8540 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8541 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X8542 VSSR sar10b_0.SWP[6] a_15533_113041# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8543 a_65769_65963# a_64993_66255# a_65333_66248# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.229 pd=1.64 as=0.24605 ps=1.405 w=0.74 l=0.15
X8544 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8545 a_61929_51311# a_60969_51311# a_61493_51596# VDDD sky130_fd_pr__pfet_01v8 ad=0.23015 pd=1.73 as=0.19062 ps=1.505 w=1 l=0.15
X8546 VDDD a_61493_51596# a_61448_51694# VDDD sky130_fd_pr__pfet_01v8 ad=0.13713 pd=1.155 as=0.0504 ps=0.66 w=0.42 l=0.15
X8547 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8548 a_66049_57307# a_65865_57675# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X8549 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X8550 a_63950_60020# a_63561_60339# a_63285_60399# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X8551 th_dif_sw_0.th_sw_1.CK a_n4470_65264# VSSA VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8552 tdc_0.RDY a_55121_59650# a_55282_59893# VDDA sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.196 ps=1.47 w=1.12 l=0.15
X8553 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8554 a_67105_61303# a_66921_61671# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X8555 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8556 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8557 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8558 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0 ps=0 w=0.42 l=1
X8559 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X8560 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8561 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8562 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8563 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2627 ps=2.19 w=0.74 l=0.15
X8564 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8565 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8566 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8567 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8568 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8569 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8570 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8571 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8572 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8573 a_64197_62956# sar10b_0.net16 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.08925 ps=0.845 w=0.42 l=0.15
X8574 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8575 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8576 a_67598_66680# a_67209_66999# a_66933_67059# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X8577 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8578 VSSR sar10b_0.SWP[7] a_10731_113461# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8579 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.168 ps=1.42 w=1.12 l=0.15
X8580 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8581 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8582 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8583 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8584 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8585 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8586 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8587 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8588 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8589 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8590 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8591 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8592 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8593 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8594 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.196 ps=1.47 w=1.12 l=0.15
X8595 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8596 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8597 VDDD sar10b_0.net13 a_65577_57971# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X8598 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8599 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8600 VDDD a_65577_51311# sar10b_0.clknet_0_CLK VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8601 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X8602 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8603 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8604 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8605 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8606 a_67688_66680# a_67209_66999# a_67598_66680# VDDD sky130_fd_pr__pfet_01v8 ad=0.0504 pd=0.66 as=0.063 ps=0.72 w=0.42 l=0.15
X8607 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X8608 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8609 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8610 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8611 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.3864 ps=2.93 w=1.12 l=0.15
X8612 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8613 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8614 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8615 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8616 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8617 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8618 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8619 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X8620 VSSR sar10b_0.SWN[4] a_25137_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8621 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8622 VSSD a_61677_63510# a_61609_63602# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.24605 ps=1.405 w=0.74 l=0.15
X8623 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X8624 a_33863_107882# sar10b_0.SWP[2] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8625 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8626 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X8627 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8628 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8629 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8630 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8631 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8632 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X8633 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8634 c1_45456_40658# m3_45124_40618# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8635 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8636 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8637 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8638 a_64993_66255# a_64809_65963# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.1295 ps=1.09 w=0.74 l=0.15
X8639 a_15533_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8640 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8641 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2627 pd=2.19 as=0.2109 ps=2.05 w=0.74 l=0.15
X8642 VDDR sar10b_0.CF[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X8643 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8644 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8645 VSSD sar10b_0.net16 a_61173_63306# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0756 pd=0.78 as=0.0441 ps=0.63 w=0.42 l=0.15
X8646 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X8647 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8648 VSSR sar10b_0.SWN[2] a_34741_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8649 VSSD sar10b_0.net16 a_63084_56643# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X8650 VSSD sar10b_0.net3 a_67020_63063# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1197 pd=1.41 as=0.0504 ps=0.66 w=0.42 l=0.15
X8651 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8652 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X8653 c1_n1140_85652# m3_n1472_85612# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8654 a_25137_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8655 VSSD sar10b_0.clk_div_0.COUNT\[0\] sar10b_0._02_ VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X8656 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8657 VSSD a_65577_51311# sar10b_0.clknet_0_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X8658 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8659 a_61773_52237# a_61491_52222# a_62134_52028# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.0504 ps=0.66 w=0.42 l=0.15
X8660 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8661 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8662 VSSR sar10b_0.SWN[1] a_39543_5779# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8663 a_66062_57022# a_65857_56931# a_65397_56643# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X8664 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8665 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8666 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.285 pd=2.57 as=0 ps=0 w=1 l=1
X8667 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8668 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X8669 a_22076_8700# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X8670 a_60747_57571# sar10b_0.net6 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X8671 a_61454_50696# a_61249_50647# a_60789_51075# VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1239 ps=1.43 w=0.42 l=0.15
X8672 VDDD a_64521_60339# a_64773_60292# VDDD sky130_fd_pr__pfet_01v8 ad=0.1428 pd=1.225 as=0.063 ps=0.72 w=0.42 l=0.15
X8673 a_63285_60399# sar10b_0.net1 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X8674 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8675 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8676 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8677 a_36482_111642# sar10b_0.CF[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.0888 pd=0.98 as=0.2109 ps=2.05 w=0.74 l=0.15
X8678 VSSD a_66153_48647# sar10b_0.clknet_1_0__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8679 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8680 a_61395_63280# sar10b_0.net4 VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1295 ps=1.09 w=0.74 l=0.15
X8681 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.168 ps=1.42 w=1.12 l=0.15
X8682 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8683 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y a_11436_8706# VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.0888 ps=0.98 w=0.74 l=0.15
X8684 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8685 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8686 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8687 c1_45456_63252# m3_45124_63212# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8688 VDDD a_62181_56768# a_62131_57058# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.0567 ps=0.69 w=0.42 l=0.15
X8689 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8690 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8691 VSSD a_68331_52243# sar10b_0._03_ VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X8692 VSSD a_64492_67433# a_64448_67302# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0777 pd=0.79 as=0.0504 ps=0.66 w=0.42 l=0.15
X8693 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 a_38665_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8694 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8695 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8696 a_63084_56643# sar10b_0.net1 a_62997_56643# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0504 pd=0.66 as=0.1197 ps=1.41 w=0.42 l=0.15
X8697 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2109 ps=2.05 w=0.74 l=0.15
X8698 w_n9655_63119# a_n8277_66083# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8699 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8700 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8701 a_61921_55975# a_61737_56343# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3136 pd=2.8 as=0.168 ps=1.42 w=1.12 l=0.15
X8702 a_10731_113461# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8703 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X8704 w_n9655_56533# a_n8277_54249# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8705 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8706 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8707 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 a_249_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8708 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2146 pd=2.06 as=0.1036 ps=1.02 w=0.74 l=0.15
X8709 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8710 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8711 VSSD a_68235_48621# sar10b_0.SWN[7] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X8712 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8713 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8714 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8715 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X8716 VSSR sar10b_0.SWP[3] a_29939_111781# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8717 a_66535_52693# a_65394_52643# a_66378_52993# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.05565 pd=0.685 as=0.1181 ps=1.035 w=0.42 l=0.15
X8718 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.2146 ps=2.06 w=0.74 l=0.15
X8719 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8720 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3864 ps=2.93 w=1.12 l=0.15
X8721 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X8722 c1_45456_78932# m3_45124_78892# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8723 c1_17216_97972# m3_16884_97932# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8724 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8725 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8726 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 a_24259_5788# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8727 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8728 a_65355_53949# sar10b_0.clknet_0_CLK VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8729 a_68841_51605# sar10b_0._15_ sar10b_0._04_ VDDD sky130_fd_pr__pfet_01v8 ad=0.2016 pd=1.48 as=0.3192 ps=2.81 w=1.12 l=0.15
X8730 VSSD sar10b_0.clk_div_0.COUNT\[0\] a_67372_52243# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.11412 pd=0.965 as=0.09625 ps=0.9 w=0.55 l=0.15
X8731 VSSA CLK a_52504_59293# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.15535 pd=1.17 as=0.1376 ps=1.14 w=0.64 l=0.15
X8732 VDDR sar10b_0.CF[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X8733 sar10b_0.clk_div_0.COUNT\[1\] a_66961_50219# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.1862 ps=1.475 w=1.12 l=0.15
X8734 a_66933_63063# sar10b_0.net44 VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.063 pd=0.72 as=0.1197 ps=1.41 w=0.42 l=0.15
X8735 VSSD sar10b_0.net16 a_65013_64695# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.21123 pd=1.45 as=0.0504 ps=0.66 w=0.42 l=0.15
X8736 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8737 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3192 pd=2.81 as=0.168 ps=1.42 w=1.12 l=0.15
X8738 a_62357_57455# a_62222_57356# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X8739 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8740 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.1036 ps=1.02 w=0.74 l=0.15
X8741 VDDD sar10b_0.net16 a_61086_61974# VDDD sky130_fd_pr__pfet_01v8 ad=0.08925 pd=0.845 as=0.063 ps=0.72 w=0.42 l=0.15
X8742 c1_45456_55218# m3_45124_55178# sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8743 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X8744 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8745 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8746 a_65966_58354# a_65577_57971# a_65301_57975# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0735 pd=0.77 as=0.1197 ps=1.41 w=0.42 l=0.15
X8747 VDDD a_65643_71265# sar10b_0.SWP[5] VDDD sky130_fd_pr__pfet_01v8 ad=0.224 pd=1.52 as=0.3304 ps=2.83 w=1.12 l=0.15
X8748 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8749 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1554 pd=1.16 as=0.1036 ps=1.02 w=0.74 l=0.15
X8750 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8751 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1036 ps=1.02 w=0.74 l=0.15
X8752 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8753 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8754 a_39543_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8755 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3192 ps=2.81 w=1.12 l=0.15
X8756 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8757 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8758 VDDD VSSD VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.275 pd=2.55 as=0 ps=0 w=1 l=1
X8759 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8760 a_66153_48647# sar10b_0.clknet_0_CLK VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3304 ps=2.83 w=1.12 l=0.15
X8761 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8762 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8763 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1221 ps=1.07 w=0.74 l=0.15
X8764 a_38665_5788# sar10b_0.SWN[1] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8765 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR sky130_fd_pr__pfet_01v8 ad=0.3864 pd=2.93 as=0.3304 ps=2.83 w=1.12 l=0.15
X8766 a_63871_61316# a_63273_61671# VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.15675 pd=1.67 as=0.15675 ps=1.67 w=0.55 l=0.15
X8767 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8768 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1221 pd=1.07 as=0.1036 ps=1.02 w=0.74 l=0.15
X8769 DATA[2] a_68946_52411# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.3304 pd=2.83 as=0.224 ps=1.52 w=1.12 l=0.15
X8770 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8771 VDDD sar10b_0.net8 a_62185_60699# VDDD sky130_fd_pr__pfet_01v8 ad=0.1197 pd=1.41 as=0.063 ps=0.72 w=0.42 l=0.15
X8772 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8773 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X8774 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8775 a_65299_52305# sar10b_0.net16 a_64780_52239# VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0672 pd=0.85 as=0.1248 ps=1.03 w=0.64 l=0.15
X8776 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 a_43467_106170# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8777 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8778 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VDDR sky130_fd_pr__pfet_01v8 ad=0.196 pd=1.47 as=0.168 ps=1.42 w=1.12 l=0.15
X8779 VSSR sar10b_0.SWP[0] a_44345_110521# VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8780 VDDD sar10b_0.net3 a_66933_59067# VDDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.4 as=0.063 ps=0.72 w=0.42 l=0.15
X8781 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8782 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8783 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8784 VDDD a_61395_52624# a_61400_52964# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3136 ps=2.8 w=1.12 l=0.15
X8785 VSSD a_62527_67630# sar10b_0.net14 VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.2109 pd=2.05 as=0.2109 ps=2.05 w=0.74 l=0.15
X8786 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8787 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8788 VSSA th_dif_sw_0.CK a_n4470_65264# VSSA sky130_fd_pr__nfet_01v8_lvt ad=0.11655 pd=1.055 as=0.1036 ps=1.02 w=0.74 l=0.15
X8789 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X8790 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8791 a_67637_56123# a_67502_56024# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.19062 pd=1.505 as=0.305 ps=2.61 w=1 l=0.15
X8792 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR VSSR sky130_fd_pr__nfet_01v8_lvt ad=0.1036 pd=1.02 as=0.1554 ps=1.16 w=0.74 l=0.15
X8793 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X8794 a_24259_5788# sar10b_0.SWN[4] VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8795 VDDD tdc_0.OUTN a_60690_54641# VDDD sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.3528 ps=2.87 w=1.12 l=0.15
X8796 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8797 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0 ps=0 w=1.5 l=0.5
X8798 a_68767_58652# a_68169_59007# VDDD VDDD sky130_fd_pr__pfet_01v8 ad=0.2478 pd=2.27 as=0.1428 ps=1.225 w=0.84 l=0.15
X8799 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VDDR VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8800 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8801 VSSD a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8802 th_dif_sw_0.VCN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8803 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 a_29061_108738# VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8804 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8805 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8806 VDDD a_61677_52854# a_61609_52946# VDDD sky130_fd_pr__pfet_01v8 ad=0.305 pd=2.61 as=0.19062 ps=1.505 w=1 l=0.15
X8807 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8808 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8809 VSSD a_60747_60235# sar10b_0.CF[3] VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1638 pd=1.2 as=0.119 ps=1.41 w=0.42 l=0.15
X8810 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM VDDR sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.58 as=0.435 ps=3.58 w=1.5 l=0.5
X8811 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sky130_fd_pr__cap_mim_m3_1 l=4 w=4
X8812 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VDDR sky130_fd_pr__pfet_01v8 ad=0.168 pd=1.42 as=0.168 ps=1.42 w=1.12 l=0.15
X8813 VSSD VDDD VSSD VSSD sky130_fd_pr__nfet_01v8_lvt ad=0.1113 pd=1.37 as=0 ps=0 w=0.42 l=1
X8814 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM VSSR sky130_fd_pr__nfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
C0 VSSR m3_n1472_31658# 0.66371f
C1 sar10b_0.net16 a_63804_67580# 0.14209f
C2 sar10b_0.CF[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP 0.166f
C3 sar10b_0.clknet_1_0__leaf_CLK sar10b_0.SWN[7] 0.0242f
C4 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP 2.92166f
C5 c1_45456_47378# VDDR 0.01151f
C6 m3_45124_50698# th_dif_sw_0.VCN 0.17339f
C7 tdc_0.phase_detector_0.pd_out_0.B tdc_0.OUTN 0.19048f
C8 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A 0.11547f
C9 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 a_249_5788# 0.07568f
C10 sar10b_0.CF[3] sar10b_0.SWP[1] 0.12237f
C11 sar10b_0.SWP[2] sar10b_0.CF[2] 2.49372f
C12 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.38989f
C13 VSSR c1_44044_21618# 0.07152f
C14 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.68875f
C15 a_60945_60609# a_61086_60642# 0.27388f
C16 sar10b_0.net16 sar10b_0.net5 0.57378f
C17 a_67055_68689# VSSD 0.15822f
C18 a_66254_57356# a_66389_57455# 0.35559f
C19 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_1684_21618# 0.0106f
C20 c1_10156_21618# th_dif_sw_0.VCN 0.13255f
C21 sar10b_0.CF[9] sar10b_0.SWP[7] 0.16188f
C22 m3_19708_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 0.48426f
C23 VSSR m3_n1472_72172# 0.66316f
C24 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A 0.41861f
C25 c1_n1140_48498# c1_n1140_47378# 0.13255f
C26 a_65996_50650# sar10b_0.net16 0.01523f
C27 a_64197_62956# sar10b_0.net16 0.2125f
C28 sar10b_0.net3 sar10b_0._07_ 0.44943f
C29 a_62697_56343# a_62949_56296# 0.27388f
C30 VSSD a_64485_56768# 0.2612f
C31 sar10b_0.net30 sar10b_0.SWN[2] 0.01009f
C32 m3_n1472_23818# VCM 0.01415f
C33 c1_n1140_74452# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C34 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP 0.02666f
C35 m3_n1472_49578# m3_n1472_48458# 0.29566f
C36 sar10b_0._00_ sar10b_0.net16 0.01749f
C37 sar10b_0.clknet_1_0__leaf_CLK sar10b_0.SWN[6] 0.08154f
C38 sar10b_0.net21 sar10b_0.net20 0.04927f
C39 sar10b_0.cyclic_flag_0.FINAL a_66825_57675# 0.01543f
C40 sar10b_0._04_ a_66865_52076# 0.0314f
C41 VSSA a_n8277_65767# 3.41645f
C42 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN 1.88527f
C43 sar10b_0.net39 sar10b_0.net11 0.02956f
C44 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.19711f
C45 a_65385_64631# sar10b_0.net13 0.0129f
C46 m3_n1472_64332# VCM 0.01412f
C47 sar10b_0.SWN[2] VSSD 0.98519f
C48 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 0.02632f
C49 VDDD sar10b_0.cyclic_flag_0.FINAL 4.48858f
C50 a_67393_66631# a_68421_66952# 0.07826f
C51 a_65061_63428# a_64809_63299# 0.27388f
C52 a_64033_63591# a_64238_63682# 0.09983f
C53 a_65301_57975# sar10b_0.net13 0.04002f
C54 sar10b_0.net2 a_61929_56639# 0.06237f
C55 VDDD a_66205_50408# 0.01232f
C56 c1_n1140_48498# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C57 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VSSR 3.96291f
C58 sar10b_0.net18 a_68562_48647# 0.29272f
C59 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] a_38665_5788# 2.68762f
C60 th_dif_sw_0.CK sar10b_0.CF[3] 0.08543f
C61 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP sar10b_0.SWP[6] 0.22363f
C62 a_65983_64966# sar10b_0.net44 0.27797f
C63 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.95198f
C64 sar10b_0.CF[4] th_dif_sw_0.VCP 0.33063f
C65 VSSD a_62222_57356# 0.12212f
C66 VSSR c1_n1140_38418# 0.04956f
C67 a_61065_51015# a_61249_50647# 0.43491f
C68 sar10b_0.net34 a_65765_50645# 0.03051f
C69 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 sar10b_0.SWN[5] 0.41984f
C70 a_64924_52385# VSSD 0.3354f
C71 sar10b_0.net16 a_61086_49986# 0.17549f
C72 m3_45124_81132# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C73 c1_45456_57458# th_dif_sw_0.VCN 0.03459f
C74 sar10b_0.net4 a_61496_52091# 0.07165f
C75 a_65957_50273# a_65861_49313# 0.12274f
C76 m3_n1472_90092# m3_n1472_88972# 0.29566f
C77 sar10b_0.net40 a_62185_66027# 0.0151f
C78 VSSR m3_8412_97932# 0.53625f
C79 m3_45124_21578# c1_45456_21618# 1.74381f
C80 m3_8412_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.63895f
C81 VDDD a_64491_71265# 0.26997f
C82 sar10b_0.net2 sar10b_0.net16 4.72049f
C83 m3_45124_56298# VDDR 0.0103f
C84 sar10b_0.net1 sar10b_0.net6 0.63077f
C85 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y 0.07183f
C86 a_64485_56768# sar10b_0.net31 0.04494f
C87 a_64233_56639# a_64831_56974# 0.06623f
C88 a_64238_63682# sar10b_0.net42 0.02218f
C89 sar10b_0.net7 a_61065_51015# 0.24406f
C90 m3_n1472_93452# c1_n1140_94612# 0.01078f
C91 m3_45124_94572# c1_45456_94612# 1.74381f
C92 VSSR m3_33828_21578# 0.52359f
C93 sar10b_0.net16 a_61609_66266# 0.15586f
C94 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.2477f
C95 sar10b_0.net18 a_68946_49747# 0.03133f
C96 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A 0.07418f
C97 VDDD a_67393_67963# 0.25559f
C98 c1_45456_52978# m3_45124_52938# 1.74381f
C99 c1_n1140_52978# m3_n1472_51818# 0.01078f
C100 c1_n1140_51858# m3_n1472_52938# 0.01078f
C101 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR 2.42866f
C102 m3_45124_96812# VDDR 0.01034f
C103 m3_45124_93452# th_dif_sw_0.VCP 0.17339f
C104 a_66825_69663# sar10b_0.net45 0.02301f
C105 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN sar10b_0.SWN[0] 0.24496f
C106 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.10847f
C107 m3_28180_97932# VCM 0.13579f
C108 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VDDR 0.83958f
C109 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.27764p
C110 sar10b_0.SWN[2] sar10b_0.CF[8] 0.13034f
C111 a_67445_60119# sar10b_0.cyclic_flag_0.FINAL 0.03175f
C112 sar10b_0.net14 sar10b_0.net43 0.17422f
C113 a_60693_51315# sar10b_0.net1 0.22198f
C114 sar10b_0.clk_div_0.COUNT\[0\] a_66961_50219# 0.05887f
C115 c1_5920_97972# VCM 0.01358f
C116 m3_32416_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C117 a_62185_52707# sar10b_0.net6 0.01556f
C118 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.74879f
C119 sar10b_0.CF[6] sar10b_0.CF[9] 0.11464f
C120 m3_45124_75532# c1_45456_74452# 0.01078f
C121 m3_n1472_74412# c1_n1140_74452# 1.74381f
C122 m3_45124_74412# c1_45456_75572# 0.01078f
C123 VSSR c1_45456_82292# 0.0935f
C124 sar10b_0.SWN[1] sar10b_0.CF[9] 0.31957f
C125 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C126 m3_18296_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.80922f
C127 sar10b_0.SWN[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 0.23954f
C128 c1_10156_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C129 m3_14060_97932# m3_15472_97932# 0.23959f
C130 sar10b_0.clknet_1_0__leaf_CLK sar10b_0.SWN[5] 0.02082f
C131 a_62837_61451# sar10b_0.net11 0.01944f
C132 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VDDR 0.95194f
C133 c1_45456_92372# c1_45456_91252# 0.13255f
C134 c1_1684_21618# m3_1352_21578# 1.74381f
C135 a_61249_53311# sar10b_0.net16 0.10331f
C136 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 2.76306f
C137 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] 1.41359f
C138 VDDD a_61493_56924# 0.20009f
C139 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A VSSR 0.39674f
C140 VDDD a_67598_62684# 0.27382f
C141 m3_4176_97932# c1_3096_97972# 0.15596f
C142 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VDDR 8.23921f
C143 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN sar10b_0.CF[7] 0.12367f
C144 VSSR m3_n1472_47338# 0.66371f
C145 a_67733_68111# a_68169_68331# 0.16939f
C146 sar10b_0.net17 a_63339_48621# 0.05778f
C147 c1_45456_66612# VDDR 0.01153f
C148 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.11339f
C149 m3_18296_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C150 sar10b_0.net33 sar10b_0._03_ 0.03841f
C151 m3_39476_21578# m3_40888_21578# 0.23959f
C152 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] sar10b_0.CF[3] 0.0136f
C153 VSSR c1_17216_21618# 0.04949f
C154 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP sar10b_0.SWP[2] 0.30836f
C155 a_61065_53679# a_61395_52624# 0.19391f
C156 sar10b_0.CF[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17717f
C157 a_62017_57307# a_62793_57675# 0.3578f
C158 VDDD a_68767_66644# 0.21881f
C159 a_62709_63063# sar10b_0.net11 0.01185f
C160 VSSR m3_n1472_87852# 0.66316f
C161 sar10b_0.clknet_0_CLK a_67084_53565# 0.01187f
C162 a_66645_60399# a_67105_59971# 0.26257f
C163 c1_n1140_56338# c1_n1140_55218# 0.13255f
C164 a_66921_60339# a_67310_60020# 0.05462f
C165 sar10b_0.CF[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 0.16034f
C166 a_63810_50901# sar10b_0.net17 0.12004f
C167 m3_n1472_31658# VDDR 0.02681f
C168 a_61249_50647# sar10b_0.net16 0.12232f
C169 a_65682_51977# a_65861_51977# 0.54426f
C170 m3_n1472_39498# VCM 0.01415f
C171 c1_n1140_90132# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C172 VSSR sar10b_0.SWP[2] 5.50483f
C173 a_66255_50749# VSSD 0.14904f
C174 VSSR c1_n1140_96852# 0.04956f
C175 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A 0.11547f
C176 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_39476_21578# 0.03017f
C177 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_22532_21578# 0.53626f
C178 VDDD a_64454_51311# 0.1391f
C179 c1_24276_21618# VCM 0.01358f
C180 a_67209_66999# a_66933_67059# 0.1263f
C181 sar10b_0.net7 sar10b_0.net16 0.65149f
C182 a_67598_58688# sar10b_0.cyclic_flag_0.FINAL 0.01473f
C183 m3_n1472_72172# VDDR 0.02674f
C184 sar10b_0.net34 a_66049_57307# 0.01081f
C185 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A 0.04073f
C186 VDDD a_60747_61567# 0.28538f
C187 m3_26768_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.30253f
C188 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A 0.10815f
C189 m3_n1472_80012# VCM 0.01412f
C190 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A 1.29717f
C191 c1_45456_24978# c1_45456_23858# 0.13255f
C192 sar10b_0.net30 sar10b_0.net1 0.1278f
C193 a_64725_68631# a_65001_68627# 0.1263f
C194 a_63967_58652# sar10b_0.net32 0.28124f
C195 VDDD a_64705_59595# 0.22277f
C196 m3_45124_26058# m3_45124_24938# 0.29566f
C197 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.11339f
C198 a_1832_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A 0.01076f
C199 VSSR c1_n1140_54098# 0.04956f
C200 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP a_44345_110521# 0.01864f
C201 a_65861_51977# sar10b_0._07_ 0.05867f
C202 sar10b_0._08_ a_64454_51311# 0.08209f
C203 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A 0.41861f
C204 a_67077_69616# VSSD 0.27141f
C205 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.40216f
C206 sar10b_0.clk_div_0.COUNT\[3\] a_67696_52265# 0.1154f
C207 m3_45124_96812# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.23379f
C208 m3_23944_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.18853f
C209 sar10b_0.net13 sar10b_0.net43 2.09953f
C210 m3_25356_21578# c1_25688_21618# 1.74381f
C211 a_62025_53679# a_62623_53324# 0.06623f
C212 m3_45124_33898# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C213 VSSA a_51603_61205# 0.06774f
C214 th_dif_sw_0.VCP sar10b_0.CF[8] 0.28586f
C215 VSSR cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 22.8983f
C216 VSSD sar10b_0.net1 4.80907f
C217 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VDDR 4.32668f
C218 VCM sar10b_0.SWP[6] 0.13076f
C219 sar10b_0.clknet_0_CLK a_65577_51311# 1.42127f
C220 m3_33828_97932# c1_34160_97972# 1.74381f
C221 VSSR m3_45124_23818# 0.63261f
C222 VSSD a_61086_61974# 0.27173f
C223 a_61153_51603# a_61358_51694# 0.09983f
C224 sar10b_0.SWN[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 0.3013f
C225 sar10b_0.net1 a_63561_60339# 0.01033f
C226 VDDD a_63745_59971# 0.22133f
C227 a_61395_49960# a_61677_50190# 0.05462f
C228 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP sar10b_0.SWP[8] 0.18137f
C229 VDDD a_65397_56643# 0.27876f
C230 c1_39808_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26825f
C231 a_9853_5788# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 0.28709f
C232 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.80358f
C233 sar10b_0.net43 a_65198_66346# 0.02484f
C234 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 sar10b_0.CF[0] 0.26333f
C235 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A 1.37694f
C236 VSSD a_61400_66284# 0.8561f
C237 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A sar10b_0.CF[2] 0.06369f
C238 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 sar10b_0.CF[8] 0.40665f
C239 c1_n1140_97972# c1_n1140_96852# 0.13255f
C240 VDDA sar10b_0.CF[1] 0.12679f
C241 sar10b_0.net42 a_64533_65967# 0.019f
C242 sar10b_0.net4 a_62185_62031# 0.04114f
C243 sar10b_0.clk_div_0.COUNT\[0\] a_65778_49979# 0.16897f
C244 a_67423_57320# sar10b_0.net35 0.26996f
C245 sar10b_0.net46 sar10b_0.net43 0.08173f
C246 m3_45124_66572# m3_45124_65452# 0.29566f
C247 VSSR m3_45124_64332# 0.63305f
C248 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP a_24259_5788# 0.14286f
C249 sar10b_0.net4 sar10b_0.net12 0.12815f
C250 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y sar10b_0.CF[4] 0.12541f
C251 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM 3.0061f
C252 sar10b_0.clknet_1_1__leaf_CLK CLK 0.12191f
C253 w_n9655_63119# a_n9133_63315# 1.49436f
C254 a_62185_52707# VSSD 0.15428f
C255 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 1.16383f
C256 m3_14060_21578# VCM 0.13579f
C257 m3_45124_83372# c1_45456_82292# 0.01078f
C258 m3_n1472_82252# c1_n1140_82292# 1.74381f
C259 m3_45124_82252# c1_45456_83412# 0.01078f
C260 VDDD sar10b_0.SWN[3] 0.17968f
C261 c1_18628_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 0.02099f
C262 m3_23944_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 0.3358f
C263 VDDD a_64149_64635# 0.29059f
C264 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.95198f
C265 c1_45456_29458# m3_45124_28298# 0.01078f
C266 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[1] 0.05939f
C267 c1_45456_28338# m3_45124_29418# 0.01078f
C268 c1_n1140_28338# m3_n1472_28298# 1.74381f
C269 sar10b_0._10_ a_65021_50292# 0.01778f
C270 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] 0.01377f
C271 VDDD a_66865_52076# 0.38363f
C272 VDDD a_60747_62899# 0.28469f
C273 VDDD a_61358_58354# 0.29057f
C274 sar10b_0.net1 sar10b_0.net31 0.01833f
C275 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C276 a_66109_51982# a_66216_52022# 0.14439f
C277 VDDD a_64188_51135# 0.44289f
C278 a_61153_58263# a_62181_58100# 0.07826f
C279 a_60969_57971# a_61929_57971# 0.03432f
C280 a_n8277_54565# th_dif_sw_0.th_sw_1.CK 0.0999f
C281 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.11339f
C282 VDDD a_66368_49417# 0.10681f
C283 a_61400_63620# sar10b_0.net40 0.02701f
C284 sar10b_0._09_ sar10b_0.net16 0.21215f
C285 c1_45456_82292# VDDR 0.01153f
C286 a_60747_57571# sar10b_0.net6 0.24329f
C287 VDDD a_60747_64605# 0.22504f
C288 m3_19708_21578# m3_21120_21578# 0.23959f
C289 sar10b_0.net3 a_67113_56343# 0.17989f
C290 a_67105_61303# a_67881_61671# 0.3578f
C291 sar10b_0.net3 a_66933_67059# 0.23094f
C292 VSSD a_66254_57356# 0.11996f
C293 VDDD a_65761_58263# 0.22676f
C294 VSSR c1_45456_30578# 0.09348f
C295 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] a_20335_112621# 0.56899f
C296 a_62025_51015# a_62623_50660# 0.06623f
C297 a_61395_63280# sar10b_0.net16 0.20358f
C298 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VCM 2.58383f
C299 VCM CLK 3.07103f
C300 m3_n1472_72172# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C301 a_64338_52411# a_64780_52239# 0.01703f
C302 VSSR m3_29592_97932# 0.49843f
C303 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A VDDR 0.60103f
C304 c1_n1140_67732# c1_n1140_66612# 0.13255f
C305 m3_29592_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.31585f
C306 sar10b_0.CF[6] a_60747_64231# 0.14263f
C307 m3_n1472_47338# VDDR 0.02681f
C308 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26364f
C309 sar10b_0.net16 sar10b_0.net45 0.0717f
C310 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A 0.28117f
C311 m3_n1472_55178# VCM 0.01415f
C312 a_66785_50875# a_67564_50907# 0.015f
C313 a_60945_52617# a_61400_52964# 0.3578f
C314 sar10b_0._08_ a_64188_51135# 0.02387f
C315 a_65061_63428# VSSD 0.2768f
C316 VDDD a_66933_64395# 0.32503f
C317 a_60969_51311# sar10b_0.net16 0.18331f
C318 a_62181_67424# sar10b_0.net16 0.20179f
C319 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A 0.03718f
C320 VSSR c1_7332_97972# 0.05923f
C321 sar10b_0.clk_div_0.COUNT\[0\] sar10b_0.net35 1.10975f
C322 sar10b_0.net34 sar10b_0.net16 0.62928f
C323 sar10b_0.CF[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP 0.20878f
C324 a_60789_51075# VSSD 0.13976f
C325 a_68169_63003# sar10b_0.net3 0.2788f
C326 sar10b_0._07_ sar10b_0._00_ 0.03895f
C327 VDDD VDDA 12.187f
C328 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_n60_21578# 0.03808f
C329 a_64818_49979# VSSD 0.21277f
C330 sar10b_0.CF[5] VCM 3.51414f
C331 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.68971f
C332 tdc_0.OUTP sar10b_0.net16 0.01003f
C333 VDDD a_61395_60616# 0.85583f
C334 a_63457_67583# a_63804_67580# 0.24999f
C335 a_63273_67295# a_63663_67678# 0.06428f
C336 a_60969_57971# sar10b_0.net4 0.2641f
C337 sar10b_0.clknet_0_CLK a_66216_49358# 0.02795f
C338 m3_n1472_87852# VDDR 0.02674f
C339 a_67502_56024# sar10b_0.net35 0.02738f
C340 m3_n1472_95692# VCM 0.01412f
C341 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 2.35116f
C342 sar10b_0.SWN[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 0.31361f
C343 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 0.20887f
C344 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04073f
C345 c1_45456_32818# c1_45456_31698# 0.13255f
C346 VDDR sar10b_0.SWP[2] 3.19104f
C347 sar10b_0.net3 sar10b_0.net26 0.02421f
C348 sar10b_0.SWN[7] sar10b_0.CF[9] 0.16032f
C349 VDDD a_68671_55988# 0.21249f
C350 sar10b_0._03_ a_66961_50219# 0.08313f
C351 c1_27100_97972# VCM 0.01358f
C352 a_64521_60339# sar10b_0.net16 0.26324f
C353 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A 0.03718f
C354 a_61400_63620# sar10b_0.net38 0.01867f
C355 m3_45124_33898# m3_45124_32778# 0.29566f
C356 sar10b_0.net16 a_66197_56924# 0.14914f
C357 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 2.53551f
C358 tdc_0.RDY CLK 0.12383f
C359 VSSR c1_n1140_73332# 0.04956f
C360 th_dif_sw_0.CKB sar10b_0.CF[1] 0.1754f
C361 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP 0.02666f
C362 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A 0.01751f
C363 m3_8412_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.63895f
C364 c1_31336_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C365 a_60693_56643# sar10b_0.net5 0.03106f
C366 a_61153_67587# a_61493_67580# 0.24088f
C367 a_60969_67295# a_62181_67424# 0.07766f
C368 c1_11568_21618# m3_12648_21578# 0.15596f
C369 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y 0.07183f
C370 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP 0.10502f
C371 m3_45124_49578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C372 sar10b_0.net38 a_61358_67678# 0.01594f
C373 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A 0.7488f
C374 VDDD a_63797_56924# 0.19465f
C375 a_65481_59303# a_66079_59638# 0.06623f
C376 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP a_9853_112162# 0.07015f
C377 a_n9133_63315# a_n8277_65767# 0.11069f
C378 tdc_0.OUTP sar10b_0.CF[3] 0.17967f
C379 sar10b_0.net3 sar10b_0._02_ 0.33477f
C380 sar10b_0.CF[5] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] 0.01367f
C381 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A 0.07183f
C382 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A 0.01751f
C383 VCM cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 3.4512f
C384 a_62181_51440# CLK 0.02193f
C385 m3_14060_97932# c1_14392_97972# 1.74381f
C386 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A 0.39559f
C387 VSSR m3_45124_39498# 0.63261f
C388 sar10b_0.SWN[6] sar10b_0.CF[9] 0.1666f
C389 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A 0.10815f
C390 sar10b_0.net47 a_67598_68012# 0.01519f
C391 a_65765_50645# a_66593_50645# 0.27469f
C392 a_66103_50668# a_65996_50650# 0.17275f
C393 a_65586_50645# a_66785_50875# 0.05767f
C394 m3_39476_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C395 VSSD a_67209_66999# 0.55635f
C396 a_63945_63003# a_64197_62956# 0.27388f
C397 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A 0.02842f
C398 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A 0.05472f
C399 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A sar10b_0.CF[4] 0.26294f
C400 VSSR c1_25688_21618# 0.05451f
C401 sar10b_0._16_ VSSD 0.35189f
C402 a_65637_64760# sar10b_0.net16 0.17428f
C403 a_67598_54692# a_67733_54791# 0.35559f
C404 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN 0.41047f
C405 VDDR cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 5.22496f
C406 m3_45124_74412# m3_45124_73292# 0.29566f
C407 VSSR m3_45124_80012# 0.63305f
C408 a_67881_60339# a_68479_59984# 0.06623f
C409 sar10b_0.net3 a_67733_54791# 0.16759f
C410 th_dif_sw_0.VCN a_51603_61205# 0.05296f
C411 m3_45124_23818# VDDR 0.0103f
C412 a_61461_56403# a_61921_55975# 0.26257f
C413 a_61737_56343# a_62126_56024# 0.05462f
C414 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN sar10b_0.SWP[0] 0.24467f
C415 VSSD a_62527_56974# 0.25159f
C416 VDDD a_62017_57307# 0.22272f
C417 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 1.29717f
C418 m3_45124_91212# c1_45456_90132# 0.01078f
C419 m3_45124_90092# c1_45456_91252# 0.01078f
C420 m3_n1472_90092# c1_n1140_90132# 1.74381f
C421 sar10b_0.clknet_1_0__leaf_CLK a_65682_49313# 0.25096f
C422 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A 0.84026f
C423 sar10b_0.net34 sar10b_0._17_ 0.03148f
C424 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 a_20335_112621# 0.36136f
C425 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C426 a_61065_53679# a_62025_53679# 0.03529f
C427 sar10b_0.CF[4] sar10b_0.SWP[0] 0.12511f
C428 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_43712_21578# 0.0162f
C429 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 21.8133f
C430 sar10b_0.net33 a_65928_53032# 0.01942f
C431 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.40046f
C432 VSSR a_43467_106170# 0.05969f
C433 c1_45456_21618# VCM 0.02045f
C434 c1_n1140_36178# m3_n1472_36138# 1.74381f
C435 c1_45456_37298# m3_45124_36138# 0.01078f
C436 c1_45456_36178# m3_45124_37258# 0.01078f
C437 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] a_24259_109594# 1.78742f
C438 a_67297_55975# a_68325_56296# 0.07826f
C439 sar10b_0.CF[9] sar10b_0.CF[7] 0.11758f
C440 m3_45124_64332# VDDR 0.01034f
C441 a_64085_60119# a_64521_60339# 0.16939f
C442 VDDD a_67733_65447# 0.21072f
C443 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.11339f
C444 sar10b_0.net2 a_60693_56643# 0.25896f
C445 a_65673_56639# a_66885_56768# 0.07766f
C446 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] sar10b_0.SWP[7] 0.22609f
C447 sar10b_0.net18 DATA[0] 0.07954f
C448 sar10b_0.net16 a_63285_60399# 0.28321f
C449 VSSD a_60747_57571# 0.34329f
C450 VSSD a_67445_61451# 0.10008f
C451 a_65525_68912# a_65961_68627# 0.16939f
C452 VDDD th_dif_sw_0.CKB 0.2905f
C453 m3_n60_21578# m3_1352_21578# 0.23959f
C454 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C455 VSSR c1_45456_46258# 0.09348f
C456 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.11339f
C457 a_64338_52411# VSSD 0.35318f
C458 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[9] 0.17717f
C459 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN sar10b_0.SWP[6] 0.20876f
C460 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 2.73845f
C461 a_66933_59067# VSSD 0.13832f
C462 m3_n1472_87852# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C463 VDDD sar10b_0._12_ 0.40096f
C464 VDDD a_65188_51977# 0.26737f
C465 c1_n1140_75572# c1_n1140_74452# 0.13255f
C466 m3_36652_21578# c1_35572_21618# 0.15596f
C467 VDDA sar10b_0.CF[2] 0.15777f
C468 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSSR 1.11894f
C469 m3_n1472_24938# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C470 sar10b_0.net35 sar10b_0.net37 0.0285f
C471 sar10b_0.net3 sar10b_0.clk_div_0.COUNT\[2\] 0.21783f
C472 c1_n1140_96852# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C473 a_67423_69308# sar10b_0._06_ 0.01747f
C474 m3_45124_97932# c1_44044_97972# 0.15596f
C475 sar10b_0.net34 a_66789_58100# 0.01301f
C476 VSSR m3_15472_21578# 0.44987f
C477 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] th_dif_sw_0.VCN 17.8827f
C478 a_55282_59893# VDDA 0.19332f
C479 sar10b_0.net3 sar10b_0.net30 0.03037f
C480 c1_45456_30578# VDDR 0.01151f
C481 m3_45124_33898# th_dif_sw_0.VCN 0.17339f
C482 a_64725_68631# sar10b_0.net41 0.01946f
C483 a_61153_67587# VSSD 0.85314f
C484 sar10b_0.SWN[5] sar10b_0.CF[9] 0.17351f
C485 sar10b_0.net3 a_66865_49412# 0.04156f
C486 a_65481_59303# VSSD 0.29342f
C487 sar10b_0.SWP[9] VCM 0.13075f
C488 VSSD DATA[1] 0.61652f
C489 sar10b_0.net19 a_68946_56639# 0.01265f
C490 a_61400_50300# sar10b_0.net1 0.05214f
C491 a_60945_49953# a_61086_49986# 0.27388f
C492 sar10b_0._03_ a_65778_49979# 0.09099f
C493 sar10b_0.SWN[7] sar10b_0.net35 0.08531f
C494 sar10b_0.CF[6] sar10b_0.SWP[2] 0.12254f
C495 sar10b_0.CF[5] sar10b_0.SWP[3] 0.12083f
C496 m3_9824_97932# VCM 0.13573f
C497 sar10b_0.net4 a_62313_61671# 0.02898f
C498 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 a_44345_5779# 0.75105f
C499 sar10b_0.net33 a_65682_49313# 0.02041f
C500 VDDD a_63871_61316# 0.20682f
C501 sar10b_0.SWP[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 0.41985f
C502 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_31336_21618# 0.0106f
C503 a_67598_54692# VSSD 0.1356f
C504 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 0.12068f
C505 c1_45456_40658# c1_45456_39538# 0.13255f
C506 c1_15804_97972# th_dif_sw_0.VCP 0.13255f
C507 sar10b_0.net3 VSSD 11.3917f
C508 sar10b_0.net2 a_61400_62288# 0.01615f
C509 m3_35240_21578# VCM 0.15231f
C510 m3_14060_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C511 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04073f
C512 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A 0.41861f
C513 m3_45124_41738# m3_45124_40618# 0.29566f
C514 VSSR c1_n1140_89012# 0.04956f
C515 a_67733_64115# sar10b_0.net3 0.16788f
C516 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A 0.42509f
C517 VSSR a_29939_111781# 2.46707f
C518 a_64609_64923# a_64949_64916# 0.24088f
C519 a_64425_64631# a_65385_64631# 0.03432f
C520 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 2.58955f
C521 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 0.5837f
C522 a_61400_66284# a_61677_66174# 0.09983f
C523 sar10b_0.SWN[6] sar10b_0.net35 0.07869f
C524 a_67798_52206# sar10b_0.clk_div_0.COUNT\[2\] 0.04351f
C525 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A a_11436_111636# 0.01076f
C526 a_61182_52404# sar10b_0.net16 0.18004f
C527 VDDD a_65765_50645# 0.97264f
C528 sar10b_0.SWP[0] VSSD 1.69971f
C529 VSSR m3_45124_55178# 0.63083f
C530 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A 1.37832f
C531 sar10b_0.net16 a_62793_57675# 0.26553f
C532 c1_n1140_31698# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C533 VDDD a_64356_51029# 0.1056f
C534 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 3.67818f
C535 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] sar10b_0.SWP[3] 0.23248f
C536 m3_n60_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.01492f
C537 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 4.35597f
C538 VSSR c1_n1140_21618# 0.07152f
C539 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A 0.43651f
C540 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.36779f
C541 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSSR 2.48681f
C542 m3_45124_64332# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C543 sar10b_0.net7 a_60693_56643# 0.01085f
C544 a_65577_57971# a_65761_58263# 0.44532f
C545 a_66666_49313# a_66865_49412# 0.29821f
C546 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A 0.42509f
C547 m3_45124_82252# m3_45124_81132# 0.29566f
C548 VSSR m3_45124_95692# 0.63305f
C549 a_68073_56343# sar10b_0.net37 0.02493f
C550 a_64609_64923# VSSD 0.86621f
C551 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 6.32799f
C552 m3_45124_39498# VDDR 0.0103f
C553 a_67798_52206# VSSD 0.28295f
C554 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A 0.60057f
C555 sar10b_0.SWP[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 0.2638f
C556 sar10b_0.CF[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A 0.26294f
C557 sar10b_0.net3 sar10b_0.net31 0.13029f
C558 a_60690_53975# sar10b_0.net5 0.02763f
C559 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP sar10b_0.SWP[9] 0.15994f
C560 sar10b_0.cyclic_flag_0.FINAL a_67598_66680# 0.01208f
C561 a_61395_64612# a_61609_64934# 0.04522f
C562 a_61086_64638# a_61400_64952# 0.07826f
C563 VSSR c1_28512_97972# 0.05685f
C564 sar10b_0._03_ sar10b_0.net35 0.02602f
C565 VDDD a_66825_69663# 0.4077f
C566 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] a_25137_5779# 0.68523f
C567 a_66537_57971# a_67135_58306# 0.06623f
C568 sar10b_0.net8 a_63045_57628# 0.02047f
C569 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_4176_21578# 0.0162f
C570 a_55282_59893# tdc_0.phase_detector_0.pd_out_0.A 0.01858f
C571 sar10b_0.clknet_1_1__leaf_CLK a_65586_50645# 0.23801f
C572 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_21120_21578# 0.45971f
C573 a_66666_49313# VSSD 0.19839f
C574 VSSR sar10b_0.SWN[3] 5.19809f
C575 c1_18628_21618# VCM 0.01358f
C576 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 1.77469f
C577 c1_45456_44018# m3_45124_45098# 0.01078f
C578 c1_45456_45138# m3_45124_43978# 0.01078f
C579 c1_n1140_44018# m3_n1472_43978# 1.74381f
C580 VDDD a_60747_60235# 0.28649f
C581 VSSD a_61086_64638# 0.27173f
C582 m3_45124_80012# VDDR 0.01034f
C583 m3_45124_76652# th_dif_sw_0.VCP 0.17339f
C584 th_dif_sw_0.CKB sar10b_0.CF[2] 0.17064f
C585 VSSD a_66537_57971# 0.2864f
C586 VDDD a_60945_61941# 0.40908f
C587 sar10b_0.net9 a_61609_60938# 0.0392f
C588 sar10b_0.SWP[0] sar10b_0.CF[8] 0.18696f
C589 sar10b_0.net34 a_65682_51977# 0.0218f
C590 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.74879f
C591 a_62933_58787# VSSD 0.09146f
C592 VDDD a_61086_65970# 0.31755f
C593 a_62593_58639# a_63369_59007# 0.3578f
C594 th_dif_sw_0.VCP th_dif_sw_0.th_sw_1.CK 0.85538f
C595 sar10b_0.net4 a_62185_64695# 0.04141f
C596 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSSR 2.51835f
C597 a_65778_49979# a_66464_50363# 0.27693f
C598 a_n8277_54249# th_dif_sw_0.th_sw_1.CKB 0.06685f
C599 sar10b_0._09_ sar10b_0._07_ 0.43136f
C600 m3_45124_66572# c1_45456_66612# 1.74381f
C601 m3_n1472_65452# c1_n1140_66612# 0.01078f
C602 m3_n1472_66572# c1_n1140_65492# 0.01078f
C603 sar10b_0.net33 sar10b_0.clknet_1_0__leaf_CLK 0.4039f
C604 VDDR a_43467_106170# 8.00721f
C605 VSSR c1_45456_65492# 0.0935f
C606 a_67598_64016# VSSD 0.13552f
C607 m3_29592_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.31585f
C608 m3_35240_97932# m3_36652_97932# 0.23959f
C609 a_67209_64335# a_68421_64288# 0.07766f
C610 a_67598_64016# a_67733_64115# 0.35559f
C611 c1_n1140_83412# c1_n1140_82292# 0.13255f
C612 m3_n1472_40618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C613 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C614 sar10b_0.net14 a_65589_69723# 0.04296f
C615 VSSD a_61086_60642# 0.25483f
C616 VDDA tdc_0.OUTN 0.41037f
C617 c1_7332_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26825f
C618 m3_25356_97932# c1_24276_97972# 0.15596f
C619 VSSD a_62949_56296# 0.27524f
C620 sar10b_0.net16 a_64238_67295# 0.25259f
C621 a_65333_66248# a_65769_65963# 0.16939f
C622 VSSR m3_n1472_30538# 0.66371f
C623 sar10b_0.net3 a_68421_65620# 0.17732f
C624 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y 0.07418f
C625 w_n9655_56533# th_dif_sw_0.th_sw_1.CKB 0.23527f
C626 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.01132f
C627 c1_45456_46258# VDDR 0.01151f
C628 m3_45124_49578# th_dif_sw_0.VCN 0.17339f
C629 sar10b_0.net34 sar10b_0._07_ 0.02809f
C630 sar10b_0.net4 a_62185_60699# 0.04013f
C631 a_67209_63003# a_67393_62635# 0.44098f
C632 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 0.01212f
C633 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 2.62306f
C634 VSSA th_dif_sw_0.th_sw_1.CKB 5.70601f
C635 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP sar10b_0.SWN[6] 0.22362f
C636 VSSR VDDA 18.0459f
C637 a_61395_60616# a_61677_60846# 0.05462f
C638 a_61086_60642# a_61400_60956# 0.07826f
C639 a_68767_54656# sar10b_0.net18 0.27376f
C640 a_66049_57307# a_66825_57675# 0.3578f
C641 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VDDR 0.95338f
C642 sar10b_0.CF[4] sar10b_0.SWP[1] 0.12245f
C643 VSSR a_38665_107026# 0.06033f
C644 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_4508_21618# 0.0106f
C645 VSSR m3_n1472_71052# 0.66316f
C646 sar10b_0.net10 a_62497_61303# 0.02354f
C647 c1_45456_48498# c1_45456_47378# 0.13255f
C648 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP a_39543_110941# 0.01676f
C649 a_66593_50645# sar10b_0.net16 0.03713f
C650 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] sar10b_0.SWN[5] 0.07354f
C651 sar10b_0.net32 sar10b_0._10_ 0.16395f
C652 a_62949_56296# a_63295_55988# 0.07649f
C653 sar10b_0.net6 sar10b_0.net5 0.0515f
C654 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A 0.42509f
C655 VSSD a_64831_56974# 0.25627f
C656 m3_n1472_22698# VCM 0.01945f
C657 VDDD a_66049_57307# 0.22783f
C658 c1_n1140_73332# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C659 m3_45124_49578# m3_45124_48458# 0.29566f
C660 sar10b_0.SWP[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 0.31361f
C661 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] a_29939_5779# 0.80139f
C662 a_62313_61671# a_63273_61671# 0.03471f
C663 a_64428_50947# a_64761_51028# 0.14439f
C664 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 0.02632f
C665 sar10b_0.CF[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A 0.03041f
C666 sar10b_0.cyclic_flag_0.FINAL a_67423_57320# 0.02491f
C667 sar10b_0._04_ sar10b_0.clk_div_0.COUNT\[1\] 0.22037f
C668 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.10847f
C669 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] a_5051_113018# 0.58622f
C670 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN 0.08512f
C671 VDDD a_64373_63584# 0.19948f
C672 a_65577_51311# a_66785_50875# 0.02199f
C673 m3_n1472_63212# VCM 0.01412f
C674 EN sar10b_0.CF[9] 4.23948f
C675 VDDD a_61065_51015# 0.81094f
C676 a_64809_63299# a_65407_63634# 0.06623f
C677 sar10b_0.net2 a_61358_57022# 0.06135f
C678 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A sar10b_0.CF[8] 0.02149f
C679 c1_n1140_47378# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C680 a_60843_52216# VSSD 0.26232f
C681 a_60693_51315# sar10b_0.net5 0.05711f
C682 sar10b_0.net32 sar10b_0.net39 0.271f
C683 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP sar10b_0.CF[7] 0.19314f
C684 sar10b_0.net19 sar10b_0.net36 0.09273f
C685 sar10b_0._00_ sar10b_0._02_ 0.08728f
C686 VSSR c1_n1140_37298# 0.04956f
C687 a_60789_51075# a_61454_50696# 0.19065f
C688 a_61065_51015# a_61589_50795# 0.04522f
C689 sar10b_0.CF[4] th_dif_sw_0.CK 0.17698f
C690 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C691 a_65861_51977# VSSD 0.56574f
C692 m3_45124_80012# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C693 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 3.0084f
C694 m3_45124_90092# m3_45124_88972# 0.29566f
C695 VSSR m3_11236_97932# 0.49843f
C696 sar10b_0.net16 a_61677_62178# 0.23618f
C697 m3_11236_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.31716f
C698 m3_45124_55178# VDDR 0.0103f
C699 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A 0.83558f
C700 sar10b_0.net4 a_61395_65944# 0.22054f
C701 a_64831_56974# sar10b_0.net31 0.2982f
C702 a_62497_61303# a_63525_61624# 0.07826f
C703 m3_45124_93452# c1_45456_94612# 0.01078f
C704 VSSR m3_36652_21578# 0.54637f
C705 VSSD a_68169_65667# 0.29048f
C706 tdc_0.phase_detector_0.pd_out_0.A tdc_0.OUTN 0.11718f
C707 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VSSR 2.53903f
C708 sar10b_0.net2 sar10b_0.net6 0.35684f
C709 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] a_43467_106170# 2.98903f
C710 VDDD a_67733_68111# 0.21129f
C711 VSSR cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 20.1986f
C712 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A VDDR 0.38427f
C713 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.59327f
C714 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VDDR 3.04089f
C715 sar10b_0.net14 a_65185_68919# 0.02561f
C716 c1_45456_51858# m3_45124_52938# 0.01078f
C717 c1_45456_52978# m3_45124_51818# 0.01078f
C718 c1_n1140_51858# m3_n1472_51818# 1.74381f
C719 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A 0.10815f
C720 sar10b_0.cyclic_flag_0.FINAL sar10b_0.net41 0.01527f
C721 m3_45124_95692# VDDR 0.01034f
C722 m3_45124_92332# th_dif_sw_0.VCP 0.17339f
C723 VDDD a_66645_60399# 0.33449f
C724 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 8.01368f
C725 m3_31004_97932# VCM 0.13579f
C726 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] c1_20040_21618# 0.02068f
C727 a_60747_58903# sar10b_0.net7 0.29413f
C728 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A 0.42509f
C729 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 0.38262f
C730 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 0.40207f
C731 a_249_113874# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 0.02167f
C732 sar10b_0.CF[1] sar10b_0.CF[3] 0.11644f
C733 a_61153_51603# sar10b_0.net1 0.10989f
C734 sar10b_0.clk_div_0.COUNT\[0\] a_66205_50408# 0.01755f
C735 c1_8744_97972# VCM 0.01358f
C736 m3_35240_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C737 sar10b_0.SWN[4] VSSA 0.24827f
C738 sar10b_0.net7 a_60690_53975# 0.0186f
C739 VSSD sar10b_0.SWP[1] 0.92685f
C740 m3_n1472_74412# c1_n1140_73332# 0.01078f
C741 m3_45124_74412# c1_45456_74452# 1.74381f
C742 m3_n1472_73292# c1_n1140_74452# 0.01078f
C743 VSSR c1_45456_81172# 0.0935f
C744 VDDR sar10b_0.SWN[3] 2.79378f
C745 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A 0.07418f
C746 m3_21120_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.07708f
C747 sar10b_0.net41 a_64491_71265# 0.07567f
C748 VSSR th_dif_sw_0.CKB 11.844f
C749 sar10b_0.cyclic_flag_0.FINAL a_67502_56024# 0.01779f
C750 c1_12980_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C751 m3_15472_97932# m3_16884_97932# 0.23959f
C752 a_61589_53459# sar10b_0.net16 0.14579f
C753 a_34741_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.01247f
C754 c1_3096_21618# m3_2764_21578# 1.74381f
C755 c1_n1140_91252# c1_n1140_90132# 0.13255f
C756 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A 0.02842f
C757 m3_n1472_56298# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C758 VDDD a_61929_56639# 0.31877f
C759 a_64705_59595# sar10b_0.net12 0.02463f
C760 sar10b_0.CF[0] VSSA 0.38778f
C761 m3_5588_97932# c1_4508_97972# 0.15596f
C762 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A 0.05472f
C763 VSSR m3_n1472_46218# 0.66371f
C764 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VDDR 3.46557f
C765 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_12472_111642# 0.01076f
C766 sar10b_0.net16 a_66825_57675# 0.26548f
C767 a_60843_52216# a_61041_52340# 0.06623f
C768 sar10b_0.SWN[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A 0.01417f
C769 sar10b_0.net17 sar10b_0.SWN[3] 0.06244f
C770 c1_45456_62132# th_dif_sw_0.VCP 0.03459f
C771 c1_45456_65492# VDDR 0.01153f
C772 m3_21120_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C773 VSSD a_63804_67580# 0.12497f
C774 a_62709_63063# a_63169_62635# 0.26257f
C775 a_62985_63003# a_63374_62684# 0.05462f
C776 m3_40888_21578# m3_42300_21578# 0.23959f
C777 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A 1.11657f
C778 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN 0.02638f
C779 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C780 VDDD sar10b_0.net16 31.3594f
C781 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR 0.41436f
C782 a_62357_57455# a_62793_57675# 0.16939f
C783 a_63169_62635# sar10b_0.net11 0.02498f
C784 VSSR m3_n1472_86732# 0.66316f
C785 sar10b_0.clknet_0_CLK sar10b_0._16_ 0.04497f
C786 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN sar10b_0.CF[2] 0.12381f
C787 c1_45456_56338# c1_45456_55218# 0.13255f
C788 VSSD sar10b_0.net5 1.5227f
C789 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR 0.36333f
C790 m3_n1472_30538# VDDR 0.02681f
C791 VDDD a_67310_61352# 0.30383f
C792 a_61589_50795# sar10b_0.net16 0.17115f
C793 m3_n1472_38378# VCM 0.01415f
C794 a_65682_51977# sar10b_0._04_ 0.09084f
C795 th_dif_sw_0.CK VSSD 0.69107f
C796 sar10b_0.net19 sar10b_0._04_ 0.04261f
C797 c1_n1140_89012# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C798 a_65996_50650# VSSD 0.01699f
C799 VSSR c1_n1140_95732# 0.04956f
C800 sar10b_0.SWP[1] sar10b_0.CF[8] 0.13856f
C801 sar10b_0.SWP[2] sar10b_0.CF[7] 0.127f
C802 a_64197_62956# VSSD 0.31604f
C803 VDDD a_67209_59007# 0.90273f
C804 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_42300_21578# 0.03017f
C805 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_25356_21578# 0.0162f
C806 VCM cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 4.06768f
C807 CLK a_51603_61205# 0.02753f
C808 VDDA VDDR 13.1273f
C809 sar10b_0._00_ VSSD 0.25341f
C810 sar10b_0.net13 a_60747_65937# 0.28423f
C811 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A 0.07418f
C812 a_52504_59293# VSSA 0.01123f
C813 w_n9655_56533# a_n8277_54249# 68.4698f
C814 c1_27100_21618# VCM 0.01358f
C815 sar10b_0._08_ sar10b_0.net16 0.17462f
C816 VDDR a_38665_107026# 7.21057f
C817 a_67113_56343# a_66837_56403# 0.1263f
C818 th_dif_sw_0.VCN th_dif_sw_0.th_sw_1.CKB 0.25346f
C819 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 2.74303f
C820 m3_n1472_71052# VDDR 0.02674f
C821 sar10b_0.net34 a_66389_57455# 0.02284f
C822 m3_n1472_78892# VCM 0.01412f
C823 m3_29592_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.53894f
C824 a_65301_57975# sar10b_0.net1 0.18555f
C825 a_n8277_54249# VSSA 22.1094f
C826 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP sar10b_0.CF[0] 0.10544f
C827 VDDD sar10b_0.CF[3] 0.46346f
C828 c1_n1140_23858# c1_n1140_22738# 0.13255f
C829 sar10b_0.net7 sar10b_0.net6 0.50633f
C830 VDDD a_60969_67295# 0.89734f
C831 sar10b_0.net13 a_65185_68919# 0.06103f
C832 VDDD a_65733_59432# 0.26904f
C833 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN sar10b_0.CF[8] 0.12367f
C834 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN 0.90176f
C835 a_68169_65667# a_68421_65620# 0.27388f
C836 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[9] 0.01887f
C837 m3_n1472_24938# m3_n1472_23818# 0.29566f
C838 VSSR c1_n1140_52978# 0.04956f
C839 a_61153_58263# sar10b_0.net38 0.02023f
C840 sar10b_0._04_ sar10b_0._07_ 0.16456f
C841 sar10b_0.net14 a_65966_58354# 0.01108f
C842 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VCM 0.12732f
C843 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR 0.95198f
C844 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A sar10b_0.CF[9] 0.06369f
C845 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN sar10b_0.SWP[1] 0.23892f
C846 sar10b_0._06_ VSSD 0.65922f
C847 sar10b_0.clk_div_0.COUNT\[3\] sar10b_0.clk_div_0.COUNT\[2\] 0.10964f
C848 VDDD a_67393_54643# 0.25362f
C849 m3_45124_95692# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C850 m3_26768_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.30253f
C851 m3_45124_97932# m3_45124_96812# 0.29566f
C852 a_68767_63980# sar10b_0.net23 0.27341f
C853 VDDA sar10b_0.SWP[7] 0.24924f
C854 m3_26768_21578# c1_27100_21618# 1.74381f
C855 sar10b_0.net33 a_65865_57675# 0.01688f
C856 w_n9655_56533# VSSA 4.24662f
C857 m3_45124_32778# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C858 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 sar10b_0.SWN[0] 0.35053f
C859 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A 0.4383f
C860 VDDD a_60747_68227# 0.28769f
C861 a_61086_49986# VSSD 0.2702f
C862 sar10b_0.net12 a_60747_64605# 0.27587f
C863 a_62025_51015# CLK 0.01329f
C864 a_66049_69295# a_66389_69443# 0.24088f
C865 sar10b_0.clknet_1_1__leaf_CLK a_65577_51311# 0.03796f
C866 a_65865_69663# a_66825_69663# 0.03529f
C867 th_dif_sw_0.CK sar10b_0.CF[8] 0.18102f
C868 m3_35240_97932# c1_35572_97972# 1.74381f
C869 VSSR m3_45124_22698# 0.63261f
C870 sar10b_0.net2 VSSD 4.06981f
C871 VCM cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 3.45121f
C872 sar10b_0.net47 a_67077_69616# 0.01042f
C873 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05939f
C874 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 0.26289f
C875 VDDD a_64085_60119# 0.20337f
C876 sar10b_0.net7 a_60693_51315# 0.02263f
C877 a_61395_49960# a_62185_50043# 0.1263f
C878 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A 0.42509f
C879 c1_42632_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26825f
C880 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 2.44658f
C881 VSSD a_61609_66266# 0.10006f
C882 a_68169_63003# a_68421_62956# 0.27388f
C883 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[3] 0.17717f
C884 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C885 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C886 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] 17.511f
C887 m3_19708_97932# th_dif_sw_0.VCP 0.01078f
C888 sar10b_0.cyclic_flag_0.FINAL sar10b_0.net37 0.04609f
C889 VDDD sar10b_0._17_ 0.60281f
C890 sar10b_0.clk_div_0.COUNT\[3\] VSSD 1.19324f
C891 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A 0.26364f
C892 m3_n1472_65452# m3_n1472_64332# 0.29566f
C893 VSSR m3_45124_63212# 0.63305f
C894 sar10b_0.CF[6] sar10b_0.SWN[3] 0.12145f
C895 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VDDR 2.60252f
C896 m3_16884_21578# VCM 0.13579f
C897 m3_n1472_81132# c1_n1140_82292# 0.01078f
C898 m3_45124_82252# c1_45456_82292# 1.74381f
C899 m3_n1472_82252# c1_n1140_81172# 0.01078f
C900 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A 1.11457f
C901 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VDDR 3.78834f
C902 a_68562_71291# sar10b_0.net46 0.06663f
C903 sar10b_0.net3 sar10b_0.clknet_0_CLK 0.03132f
C904 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.11339f
C905 sar10b_0.net39 sar10b_0.net40 0.86362f
C906 sar10b_0.net45 a_66933_67059# 0.02615f
C907 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 sar10b_0.CF[3] 0.40665f
C908 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] a_14655_5788# 1.18623f
C909 sar10b_0.net3 a_68421_68284# 0.17518f
C910 VDDD a_67696_52265# 0.40621f
C911 c1_n1140_27218# m3_n1472_28298# 0.01078f
C912 c1_45456_28338# m3_45124_28298# 1.74381f
C913 c1_n1140_28338# m3_n1472_27178# 0.01078f
C914 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 sar10b_0.CF[5] 0.26311f
C915 VDDD sar10b_0.clk_div_0.COUNT\[1\] 1.07817f
C916 a_63745_59971# sar10b_0.net41 0.06853f
C917 a_61249_53311# VSSD 0.85322f
C918 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45324f
C919 a_67310_60020# sar10b_0.net3 0.22845f
C920 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[0] 0.01902f
C921 a_61493_58256# a_61929_57971# 0.16939f
C922 a_60969_57971# a_61358_58354# 0.06034f
C923 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 sar10b_0.SWP[9] 0.2346f
C924 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C925 c1_45456_81172# VDDR 0.01153f
C926 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[0] 0.17732f
C927 VDDA a_51345_60437# 0.65552f
C928 a_67445_61451# a_67881_61671# 0.16939f
C929 VDDR th_dif_sw_0.CKB 0.22815f
C930 m3_21120_21578# m3_22532_21578# 0.23959f
C931 VDDD a_60945_64605# 0.4075f
C932 sar10b_0.net38 a_62997_56643# 0.0667f
C933 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] a_15533_113041# 0.45291f
C934 VSSR c1_45456_29458# 0.09348f
C935 VDDD a_66789_58100# 0.28277f
C936 sar10b_0._10_ CLK 0.04062f
C937 a_61086_63306# sar10b_0.net16 0.17802f
C938 m3_n1472_71052# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C939 a_61035_48621# VSSD 0.30423f
C940 a_66933_63063# sar10b_0.net44 0.1743f
C941 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.41861f
C942 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A 0.02842f
C943 sar10b_0.clknet_1_0__leaf_CLK a_65778_49979# 0.24476f
C944 a_64780_52239# sar10b_0._09_ 0.11155f
C945 VSSR m3_32416_97932# 0.49843f
C946 c1_45456_67732# c1_45456_66612# 0.13255f
C947 sar10b_0.clk_div_0.COUNT\[1\] sar10b_0._08_ 0.37323f
C948 VDDD a_62798_58688# 0.26812f
C949 m3_32416_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.3309f
C950 m3_n1472_46218# VDDR 0.02681f
C951 a_61491_52222# sar10b_0.net1 0.0109f
C952 VSSA a_53652_61050# 0.20064f
C953 m3_n1472_54058# VCM 0.01415f
C954 a_60945_52617# a_61609_52946# 0.16939f
C955 a_61395_52624# a_61677_52854# 0.05462f
C956 a_65407_63634# VSSD 0.27276f
C957 a_61493_51596# sar10b_0.net16 0.15576f
C958 a_67209_59007# a_67598_58688# 0.05462f
C959 VDDD a_67393_63967# 0.24943f
C960 a_66933_59067# a_67393_58639# 0.26257f
C961 a_62527_67630# sar10b_0.net16 0.02498f
C962 sar10b_0.CF[0] th_dif_sw_0.VCN 0.28582f
C963 sar10b_0.CF[6] VDDA 0.39306f
C964 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A 0.05105f
C965 VSSR c1_10156_97972# 0.06746f
C966 a_64149_64635# sar10b_0.net41 0.01534f
C967 a_61249_50647# VSSD 0.85194f
C968 sar10b_0.net16 a_64809_65963# 0.17341f
C969 a_43467_5788# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 0.23957f
C970 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A 0.95262f
C971 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_2764_21578# 0.03017f
C972 sar10b_0.CF[3] sar10b_0.CF[2] 48.4706f
C973 sar10b_0.SWN[9] DATA[1] 0.08532f
C974 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM 4.85257f
C975 sar10b_0.net23 sar10b_0.net25 0.24631f
C976 c1_272_21618# VCM 0.01358f
C977 sar10b_0.net38 sar10b_0.net39 2.68565f
C978 a_63797_56924# a_63662_57022# 0.35559f
C979 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR 0.38833f
C980 VDDD a_60945_60609# 0.40714f
C981 a_63457_67583# a_64238_67295# 0.35777f
C982 a_61493_58256# sar10b_0.net4 0.05296f
C983 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 7.2266f
C984 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 1.88521f
C985 m3_n1472_86732# VDDR 0.02674f
C986 VDDD a_62697_56343# 0.35983f
C987 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR 0.59833f
C988 m3_n1472_94572# VCM 0.01412f
C989 a_60747_65937# a_60945_65937# 0.06623f
C990 th_dif_sw_0.th_sw_1.CKB a_n9133_63315# 0.42326f
C991 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A sar10b_0.CF[8] 0.03041f
C992 a_66865_52076# sar10b_0.clk_div_0.COUNT\[0\] 0.08529f
C993 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 sar10b_0.CF[7] 0.40665f
C994 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] th_dif_sw_0.VCN 1.10485p
C995 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.38218f
C996 sar10b_0.net7 VSSD 2.51539f
C997 c1_n1140_31698# c1_n1140_30578# 0.13255f
C998 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 0.53683f
C999 sar10b_0._03_ a_66205_50408# 0.13181f
C1000 c1_29924_97972# VCM 0.01358f
C1001 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VSSR 20.1987f
C1002 a_61609_63602# sar10b_0.net38 0.02174f
C1003 m3_n1472_32778# m3_n1472_31658# 0.29566f
C1004 sar10b_0.net3 a_67881_61671# 0.293f
C1005 sar10b_0.net16 a_66633_56639# 0.26652f
C1006 VSSR c1_n1140_72212# 0.04956f
C1007 a_68235_71265# sar10b_0.net45 0.27814f
C1008 a_65355_53949# VSSD 2.2902f
C1009 VDDD a_65390_69010# 0.26034f
C1010 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.39384f
C1011 a_67744_51002# VSSD 0.01142f
C1012 sar10b_0.net33 sar10b_0._01_ 0.25417f
C1013 m3_11236_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.31716f
C1014 c1_34160_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C1015 a_68169_68331# VSSD 0.29131f
C1016 a_67393_58639# sar10b_0.net3 0.11379f
C1017 a_60693_51315# a_60969_51311# 0.1263f
C1018 a_61153_67587# a_61929_67295# 0.3578f
C1019 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A 0.11547f
C1020 c1_12980_21618# m3_14060_21578# 0.15596f
C1021 m3_45124_48458# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C1022 VDDD a_64233_56639# 0.32963f
C1023 a_66079_59638# sar10b_0.net34 0.27457f
C1024 a_n8277_66083# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 1.13669f
C1025 a_67105_59971# VSSD 0.85295f
C1026 m3_15472_97932# c1_15804_97972# 1.74381f
C1027 a_62527_51646# CLK 0.01981f
C1028 VSSD a_68946_56639# 0.33159f
C1029 VSSR m3_45124_38378# 0.63261f
C1030 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A 0.10815f
C1031 sar10b_0.CF[4] tdc_0.OUTP 0.27745f
C1032 sar10b_0.clknet_1_0__leaf_CLK sar10b_0.net35 0.33439f
C1033 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.43131f
C1034 VSSA a_52417_60961# 0.14575f
C1035 sar10b_0.net33 a_65778_49979# 0.02339f
C1036 m3_42300_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C1037 a_66837_56403# VSSD 0.13927f
C1038 a_68331_52243# a_68946_52411# 0.02515f
C1039 a_64197_62956# a_64543_62648# 0.07649f
C1040 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C1041 a_62187_48621# sar10b_0.SWN[2] 0.15514f
C1042 VSSR c1_28512_21618# 0.05685f
C1043 a_67393_54643# a_68169_55011# 0.3578f
C1044 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] a_34741_111361# 0.91754f
C1045 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A 0.38427f
C1046 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 a_10731_5779# 0.20413f
C1047 m3_n1472_73292# m3_n1472_72172# 0.29566f
C1048 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 0.40665f
C1049 VSSR m3_45124_78892# 0.63305f
C1050 a_65577_57971# sar10b_0.net16 0.19011f
C1051 sar10b_0.net34 a_65857_56931# 0.0251f
C1052 sar10b_0.net40 sar10b_0.net11 0.02673f
C1053 m3_45124_22698# VDDR 0.0103f
C1054 sar10b_0.net8 a_62497_61303# 0.06724f
C1055 VDDD a_62357_57455# 0.2051f
C1056 sar10b_0.net32 sar10b_0.SWN[4] 0.01678f
C1057 m3_n1472_90092# c1_n1140_89012# 0.01078f
C1058 m3_n1472_88972# c1_n1140_90132# 0.01078f
C1059 m3_45124_90092# c1_45456_90132# 1.74381f
C1060 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR 2.40416f
C1061 a_68421_62956# VSSD 0.27186f
C1062 VSSA th_dif_sw_0.VCN 9.49539f
C1063 VDDD a_65682_51977# 0.40622f
C1064 VDDD sar10b_0.net19 1.1114f
C1065 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 a_15533_113041# 0.28343f
C1066 sar10b_0.SWP[4] VDDD 0.35153f
C1067 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C1068 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A 0.39559f
C1069 sar10b_0.net16 a_61677_64842# 0.22675f
C1070 sar10b_0.net2 a_64492_67433# 0.0229f
C1071 sar10b_0.SWN[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP 0.30835f
C1072 VSSD DATA[2] 0.59996f
C1073 c1_n1140_93492# c1_n1140_94612# 0.13255f
C1074 c1_45456_36178# m3_45124_36138# 1.74381f
C1075 c1_n1140_36178# m3_n1472_35018# 0.01078f
C1076 c1_n1140_35058# m3_n1472_36138# 0.01078f
C1077 m3_45124_63212# VDDR 0.01034f
C1078 sar10b_0.clk_div_0.COUNT\[1\] sar10b_0._15_ 0.06704f
C1079 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.12357f
C1080 a_63621_58960# sar10b_0.net16 0.17344f
C1081 sar10b_0.net7 a_61041_52340# 0.01908f
C1082 a_65857_56931# a_66197_56924# 0.24088f
C1083 a_n9133_57045# th_dif_sw_0.th_sw_1.CKB 0.42326f
C1084 sar10b_0.CF[6] th_dif_sw_0.CKB 0.08605f
C1085 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A 0.95194f
C1086 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] 2.78254f
C1087 a_62133_59067# sar10b_0.net39 0.06074f
C1088 th_dif_sw_0.CKB sar10b_0.SWN[1] 0.09905f
C1089 c1_28512_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.26825f
C1090 a_65865_69663# sar10b_0.net16 0.18948f
C1091 a_66213_68756# a_66559_68962# 0.07649f
C1092 m3_1352_21578# m3_2764_21578# 0.23959f
C1093 sar10b_0._05_ a_65394_52643# 0.08239f
C1094 sar10b_0.net19 sar10b_0._08_ 0.03079f
C1095 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM 1.75389f
C1096 VSSR c1_45456_45138# 0.09348f
C1097 sar10b_0.net14 sar10b_0.net39 0.05682f
C1098 sar10b_0._09_ VSSD 0.71276f
C1099 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP sar10b_0.CF[8] 0.10502f
C1100 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A 0.41861f
C1101 sar10b_0.net16 a_61677_60846# 0.23706f
C1102 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 0.21775f
C1103 m3_n1472_86732# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C1104 VDDD sar10b_0._07_ 0.97274f
C1105 c1_45456_75572# c1_45456_74452# 0.13255f
C1106 sar10b_0.net34 a_66865_49412# 0.081f
C1107 VDDD DATA[5] 0.35476f
C1108 m3_38064_21578# c1_36984_21618# 0.15596f
C1109 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A sar10b_0.CF[9] 0.26294f
C1110 sar10b_0.clknet_0_CLK a_65861_51977# 0.01386f
C1111 m3_n1472_23818# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C1112 sar10b_0.SWP[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A 0.01506f
C1113 a_61395_63280# VSSD 0.51666f
C1114 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A 0.28117f
C1115 sar10b_0.net38 sar10b_0.net11 0.02621f
C1116 a_62997_56643# a_63457_56931# 0.26257f
C1117 c1_n1140_95732# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C1118 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A 1.29796f
C1119 VSSR m3_18296_21578# 0.39907f
C1120 c1_22864_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 0.01334f
C1121 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A 0.10815f
C1122 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C1123 sar10b_0.net45 VSSD 1.16053f
C1124 c1_45456_29458# VDDR 0.01151f
C1125 m3_45124_32778# th_dif_sw_0.VCN 0.17339f
C1126 a_60969_51311# VSSD 0.48409f
C1127 a_62181_67424# VSSD 0.27002f
C1128 sar10b_0.net34 VSSD 1.56686f
C1129 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17717f
C1130 sar10b_0.CF[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP 0.16021f
C1131 tdc_0.OUTN sar10b_0.CF[3] 0.56605f
C1132 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A sar10b_0.CF[8] 0.06369f
C1133 a_61086_49986# a_61400_50300# 0.07826f
C1134 sar10b_0._07_ sar10b_0._08_ 0.84246f
C1135 m3_12648_97932# VCM 0.13579f
C1136 sar10b_0.SWP[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 0.39898f
C1137 tdc_0.OUTP VSSD 1.33537f
C1138 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A 0.05472f
C1139 sar10b_0.SWN[2] VCM 0.13074f
C1140 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_34160_21618# 0.0106f
C1141 c1_n1140_39538# c1_n1140_38418# 0.13255f
C1142 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.02638f
C1143 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A a_1832_111636# 0.01076f
C1144 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[1] 0.01887f
C1145 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 sar10b_0.SWN[6] 0.39899f
C1146 c1_18628_97972# th_dif_sw_0.VCP 0.13255f
C1147 VDDD a_63457_67583# 0.24365f
C1148 a_61400_62288# a_61677_62178# 0.09983f
C1149 sar10b_0.net39 a_63457_56931# 0.02517f
C1150 m3_38064_21578# VCM 0.15231f
C1151 VSSR sar10b_0.CF[3] 19.7771f
C1152 m3_16884_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C1153 a_68946_59303# sar10b_0.net22 0.02944f
C1154 m3_n1472_40618# m3_n1472_39498# 0.29566f
C1155 sar10b_0._12_ a_67611_50645# 0.07728f
C1156 VSSR c1_n1140_87892# 0.04956f
C1157 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26364f
C1158 sar10b_0.SWN[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 0.29562f
C1159 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.02632f
C1160 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 4.3082f
C1161 a_64521_60339# VSSD 0.28722f
C1162 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A 0.43728f
C1163 VSSD a_66197_56924# 0.1003f
C1164 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 a_34741_111361# 0.59518f
C1165 a_64425_64631# a_64814_65014# 0.06034f
C1166 VDDD a_60693_56643# 0.31734f
C1167 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C1168 a_64609_64923# a_65385_64631# 0.3578f
C1169 sar10b_0.net47 sar10b_0.net3 0.23747f
C1170 a_61609_66266# a_61677_66174# 0.35559f
C1171 sar10b_0.clk_div_0.COUNT\[0\] sar10b_0._12_ 0.10327f
C1172 a_61400_66284# a_62185_66027# 0.26257f
C1173 sar10b_0.net21 a_68421_54964# 0.022f
C1174 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C1175 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.59283f
C1176 a_64521_60339# a_63561_60339# 0.03471f
C1177 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] a_38665_107026# 2.68762f
C1178 a_61035_48621# sar10b_0.SWN[0] 0.04462f
C1179 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSSR 6.0472f
C1180 a_61496_52091# sar10b_0.net16 0.11837f
C1181 VDDD a_66103_50668# 0.15622f
C1182 VDDD a_63945_63003# 0.35368f
C1183 VSSR m3_45124_54058# 0.63261f
C1184 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A 0.28117f
C1185 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VDDR 3.78835f
C1186 c1_n1140_30578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C1187 m3_2764_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C1188 a_66933_63063# sar10b_0.cyclic_flag_0.FINAL 0.06686f
C1189 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP 0.02666f
C1190 sar10b_0.net41 a_63871_61316# 0.27484f
C1191 VSSR c1_1684_21618# 0.05923f
C1192 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.11339f
C1193 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VCM 2.33869f
C1194 m3_45124_63212# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C1195 a_66865_49412# a_67371_49579# 0.0192f
C1196 a_65577_57971# a_66789_58100# 0.07766f
C1197 tdc_0.OUTP sar10b_0.CF[8] 0.17891f
C1198 m3_n1472_81132# m3_n1472_80012# 0.29566f
C1199 VSSR m3_45124_94572# 0.63305f
C1200 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A 0.11547f
C1201 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.36435f
C1202 a_65637_64760# VSSD 0.27401f
C1203 sar10b_0.net10 sar10b_0.net39 0.02514f
C1204 m3_45124_38378# VDDR 0.0103f
C1205 a_65001_68627# sar10b_0.net16 0.21148f
C1206 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.02632f
C1207 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.11339f
C1208 sar10b_0.net13 sar10b_0.net39 0.05733f
C1209 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 0.20006f
C1210 a_68169_59007# a_68767_58652# 0.06623f
C1211 VSSR c1_31336_97972# 0.05685f
C1212 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] sar10b_0.SWN[9] 0.22371f
C1213 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] m3_19708_97932# 0.13306f
C1214 VDDD a_67423_69308# 0.22511f
C1215 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP 0.02666f
C1216 sar10b_0.net19 sar10b_0._15_ 0.21126f
C1217 a_67135_58306# sar10b_0.net36 0.275f
C1218 m3_32416_21578# th_dif_sw_0.VCN 0.01078f
C1219 a_67371_49579# VSSD 0.30708f
C1220 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_23944_21578# 0.03017f
C1221 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_7000_21578# 0.0162f
C1222 VSSA a_n9133_63315# 0.87222f
C1223 a_61041_52340# a_60969_51311# 0.01304f
C1224 sar10b_0.SWN[3] sar10b_0.CF[7] 0.12514f
C1225 sar10b_0.net26 a_68946_65963# 0.26142f
C1226 c1_45456_44018# m3_45124_43978# 1.74381f
C1227 c1_n1140_42898# m3_n1472_43978# 0.01078f
C1228 c1_n1140_44018# m3_n1472_42858# 0.01078f
C1229 VDDD a_60945_49953# 0.40485f
C1230 a_61677_63510# a_62185_63363# 0.19065f
C1231 m3_45124_78892# VDDR 0.01034f
C1232 sar10b_0.net12 a_66049_57307# 0.0155f
C1233 m3_45124_75532# th_dif_sw_0.VCP 0.17339f
C1234 VSSD sar10b_0.net36 3.49298f
C1235 VDDD a_61400_62288# 0.25246f
C1236 m3_11236_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.53633f
C1237 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VSSR 3.55942f
C1238 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A 1.3401f
C1239 sar10b_0.SWP[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.45618f
C1240 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN 0.01165f
C1241 a_62933_58787# a_63369_59007# 0.16939f
C1242 CLK th_dif_sw_0.th_sw_1.CKB 0.24353f
C1243 a_65778_49979# a_66961_50219# 0.0649f
C1244 a_67209_65667# a_67598_65348# 0.05462f
C1245 a_66933_65727# a_67393_65299# 0.26257f
C1246 a_68562_71291# CKO 0.1431f
C1247 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A 0.60057f
C1248 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04073f
C1249 m3_45124_65452# c1_45456_66612# 0.01078f
C1250 m3_45124_66572# c1_45456_65492# 0.01078f
C1251 m3_n1472_65452# c1_n1140_65492# 1.74381f
C1252 VSSR c1_45456_64372# 0.0935f
C1253 VSSD a_63285_60399# 0.142f
C1254 sar10b_0.net4 a_62281_52347# 0.05536f
C1255 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.39835f
C1256 sar10b_0.net13 a_65333_66248# 0.02093f
C1257 m3_32416_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.3309f
C1258 m3_36652_97932# m3_38064_97932# 0.23959f
C1259 a_67393_63967# a_68169_64335# 0.3578f
C1260 c1_45456_83412# c1_45456_82292# 0.13255f
C1261 a_63561_60339# a_63285_60399# 0.1263f
C1262 th_dif_sw_0.VCP VCM 2.8337f
C1263 a_61249_53311# a_61454_53360# 0.09983f
C1264 VDDD a_65394_52643# 0.43391f
C1265 m3_n1472_39498# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C1266 m3_18296_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.80922f
C1267 sar10b_0.net14 a_66049_69295# 0.02005f
C1268 c1_10156_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.01541f
C1269 sar10b_0.net20 sar10b_0.net36 0.16164f
C1270 m3_26768_97932# c1_25688_97972# 0.15596f
C1271 VSSR m3_n1472_29418# 0.66371f
C1272 a_65333_66248# a_65198_66346# 0.35559f
C1273 a_66021_66092# a_66367_66298# 0.07649f
C1274 sar10b_0.net16 a_63663_67678# 0.22385f
C1275 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A 1.37879f
C1276 c1_45456_45138# VDDR 0.01151f
C1277 a_67209_66999# a_67393_66631# 0.44098f
C1278 m3_45124_48458# th_dif_sw_0.VCN 0.17339f
C1279 a_65045_59588# a_64910_59686# 0.35559f
C1280 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VCM 0.12074f
C1281 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN 0.01152f
C1282 sar10b_0.net18 a_68946_53975# 0.03194f
C1283 a_n8277_54249# a_n9133_57045# 0.97211f
C1284 a_66933_63063# a_67598_62684# 0.19065f
C1285 a_67209_63003# a_67733_62783# 0.04522f
C1286 a_35446_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.01076f
C1287 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VSSR 1.37544f
C1288 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A 0.05472f
C1289 a_61395_60616# a_62185_60699# 0.1263f
C1290 VDDA sar10b_0.CF[7] 0.39307f
C1291 a_66389_57455# a_66825_57675# 0.16939f
C1292 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_7332_21618# 0.0106f
C1293 c1_15804_21618# th_dif_sw_0.VCN 0.13255f
C1294 VSSR m3_n1472_69932# 0.66316f
C1295 sar10b_0.net3 sar10b_0.net43 0.13233f
C1296 c1_n1140_47378# c1_n1140_46258# 0.13255f
C1297 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A a_25842_111636# 0.01076f
C1298 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A 0.74881f
C1299 VSSR a_5929_113881# 0.77753f
C1300 sar10b_0.clknet_0_CLK sar10b_0.clk_div_0.COUNT\[3\] 0.02709f
C1301 m3_n1472_21578# VCM 0.16646f
C1302 VDDD a_66389_57455# 0.20777f
C1303 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR 1.10847f
C1304 c1_n1140_72212# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C1305 m3_n1472_48458# m3_n1472_47338# 0.29566f
C1306 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] th_dif_sw_0.VCP 70.5858f
C1307 w_n9655_56533# a_n9133_57045# 1.49436f
C1308 sar10b_0._04_ sar10b_0.clk_div_0.COUNT\[2\] 0.28942f
C1309 sar10b_0.net4 a_61400_52964# 0.05656f
C1310 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A 0.39629f
C1311 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 sar10b_0.SWN[6] 0.27668f
C1312 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A VSSR 0.39674f
C1313 VSSA a_n9133_57045# 0.87222f
C1314 a_66961_50219# sar10b_0.net35 0.02586f
C1315 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] a_5929_5779# 0.22044f
C1316 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 21.6018f
C1317 VDDD a_64809_63299# 0.36072f
C1318 m3_n1472_62092# VCM 0.01412f
C1319 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A 0.05472f
C1320 sar10b_0.net19 a_68946_49747# 0.25539f
C1321 sar10b_0.net10 a_62709_63063# 0.06345f
C1322 VDDR sar10b_0.CF[3] 1.70274f
C1323 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 0.30288f
C1324 VDDD a_66762_50329# 0.10132f
C1325 c1_n1140_46258# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C1326 a_61153_51603# sar10b_0.net5 0.01585f
C1327 a_61182_52404# VSSD 0.26904f
C1328 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A VDDR 0.38397f
C1329 VSSD a_62793_57675# 0.27102f
C1330 VSSR c1_n1140_36178# 0.04956f
C1331 sar10b_0.net10 sar10b_0.net11 1.39736f
C1332 a_61249_50647# a_61454_50696# 0.09983f
C1333 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS th_dif_sw_0.th_sw_1.CKB 0.35456f
C1334 a_64609_64923# sar10b_0.net43 0.02568f
C1335 sar10b_0._04_ VSSD 0.39873f
C1336 sar10b_0.net16 a_61677_50190# 0.23982f
C1337 m3_45124_78892# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C1338 sar10b_0.CF[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP 0.1053f
C1339 VDDD a_60747_58903# 0.28292f
C1340 m3_n1472_88972# m3_n1472_87852# 0.29566f
C1341 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VDDR 3.50612f
C1342 VSSR m3_14060_97932# 0.49683f
C1343 sar10b_0.net16 a_62185_62031# 0.22212f
C1344 m3_14060_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.31585f
C1345 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A 0.05472f
C1346 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP sar10b_0.SWP[3] 0.28713f
C1347 m3_45124_54058# VDDR 0.0103f
C1348 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A sar10b_0.CF[3] 0.02149f
C1349 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A sar10b_0.CF[5] 0.03041f
C1350 VDDD a_60690_53975# 0.54105f
C1351 VSSR m3_39476_21578# 0.54637f
C1352 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP 1.16923f
C1353 sar10b_0.net16 sar10b_0.net12 1.08622f
C1354 VSSD a_68767_65312# 0.26804f
C1355 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN sar10b_0.CF[9] 0.12367f
C1356 c1_n1140_51858# m3_n1472_50698# 0.01078f
C1357 c1_n1140_50738# m3_n1472_51818# 0.01078f
C1358 sar10b_0.SWP[4] VSSR 4.79472f
C1359 c1_45456_51858# m3_45124_51818# 1.74381f
C1360 VSSD a_68946_65963# 0.33161f
C1361 sar10b_0.CF[5] sar10b_0.SWN[4] 0.11875f
C1362 sar10b_0.CF[0] CLK 0.18538f
C1363 m3_45124_91212# th_dif_sw_0.VCP 0.17339f
C1364 m3_45124_94572# VDDR 0.01034f
C1365 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.59739f
C1366 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A 0.45324f
C1367 m3_33828_97932# VCM 0.15071f
C1368 a_65643_71265# VSSD 0.33898f
C1369 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 0.90172f
C1370 sar10b_0.CF[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN 0.10438f
C1371 sar10b_0.net3 a_67393_66631# 0.1112f
C1372 VDDD a_67113_56343# 0.89606f
C1373 VDDD a_66933_67059# 0.32565f
C1374 a_62181_51440# sar10b_0.net1 0.0155f
C1375 VDDA th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 0.12838f
C1376 c1_11568_97972# VCM 0.01358f
C1377 m3_38064_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C1378 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP a_39543_5779# 0.01676f
C1379 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y sar10b_0.CF[3] 0.12541f
C1380 sar10b_0.net16 a_63662_57022# 0.22534f
C1381 m3_45124_74412# c1_45456_73332# 0.01078f
C1382 m3_45124_73292# c1_45456_74452# 0.01078f
C1383 m3_n1472_73292# c1_n1140_73332# 1.74381f
C1384 VSSR c1_45456_80052# 0.0935f
C1385 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.38722f
C1386 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.5837f
C1387 sar10b_0.CF[5] sar10b_0.CF[0] 0.11689f
C1388 m3_23944_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.09358f
C1389 sar10b_0.CF[4] sar10b_0.CF[1] 0.11415f
C1390 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 1.79797f
C1391 sar10b_0.net46 a_66049_69295# 0.01942f
C1392 th_dif_sw_0.CKB sar10b_0.CF[7] 0.08666f
C1393 c1_15804_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C1394 a_64491_48621# sar10b_0.SWN[4] 0.17846f
C1395 a_65355_53949# sar10b_0.clknet_0_CLK 0.50561f
C1396 m3_16884_97932# m3_18296_97932# 0.23959f
C1397 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A 0.02842f
C1398 sar10b_0.net2 a_64533_65967# 0.2264f
C1399 c1_45456_91252# c1_45456_90132# 0.13255f
C1400 c1_4508_21618# m3_4176_21578# 1.74381f
C1401 m3_n1472_55178# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C1402 a_65001_68627# a_65390_69010# 0.06034f
C1403 sar10b_0._03_ sar10b_0._12_ 0.2457f
C1404 VDDD a_61358_57022# 0.27761f
C1405 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VDDR 3.71081f
C1406 a_64521_59303# a_64705_59595# 0.44532f
C1407 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A 0.76105f
C1408 VDDD a_68169_63003# 0.36697f
C1409 m3_7000_97932# c1_5920_97972# 0.15596f
C1410 VSSR m3_n1472_45098# 0.66371f
C1411 a_68169_68331# a_68421_68284# 0.27388f
C1412 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A 0.07183f
C1413 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A 0.01751f
C1414 sar10b_0.SWP[8] sar10b_0.SWP[9] 21.3566f
C1415 a_61041_52340# a_61182_52404# 0.27388f
C1416 c1_45456_64372# VDDR 0.01153f
C1417 sar10b_0.net21 sar10b_0.net22 0.13043f
C1418 m3_23944_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C1419 a_66645_60399# sar10b_0.net41 0.17955f
C1420 sar10b_0.CF[6] sar10b_0.net16 0.01525f
C1421 VSSD a_64238_67295# 0.30902f
C1422 a_62181_58100# sar10b_0.net40 0.02272f
C1423 sar10b_0._05_ VSSD 0.26664f
C1424 m3_42300_21578# m3_43712_21578# 0.23959f
C1425 a_n8277_54249# CLK 0.17329f
C1426 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A sar10b_0.CF[7] 0.02149f
C1427 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 2.74732f
C1428 VDDD sar10b_0.net26 0.52164f
C1429 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A 0.45324f
C1430 VSSR m3_n1472_85612# 0.66316f
C1431 a_60969_57971# sar10b_0.net16 0.16385f
C1432 a_66921_60339# a_67881_60339# 0.03471f
C1433 a_67105_59971# a_67310_60020# 0.09983f
C1434 c1_n1140_55218# c1_n1140_54098# 0.13255f
C1435 VDDD sar10b_0.net6 2.01297f
C1436 m3_n1472_29418# VDDR 0.02681f
C1437 a_60747_69559# sar10b_0.CF[9] 0.14208f
C1438 m3_n1472_37258# VCM 0.01415f
C1439 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A sar10b_0.CF[0] 0.03041f
C1440 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A 0.83578f
C1441 c1_n1140_87892# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C1442 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 5.16397f
C1443 m3_n1472_56298# m3_n1472_55178# 0.29566f
C1444 VDDD a_64780_52239# 0.2043f
C1445 a_66593_50645# VSSD 0.19194f
C1446 VSSR c1_n1140_94612# 0.04956f
C1447 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A 0.05472f
C1448 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VDDR 0.84106f
C1449 a_9853_112162# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 0.28709f
C1450 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_28180_21578# 0.0162f
C1451 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_45124_21578# 0.03017f
C1452 a_53652_59132# VSSA 0.20064f
C1453 c1_29924_21618# VCM 0.01358f
C1454 sar10b_0.net4 a_60969_56639# 0.02979f
C1455 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C1456 VDDD a_60747_63273# 0.22504f
C1457 VDDD sar10b_0._02_ 0.37717f
C1458 m3_n1472_69932# VDDR 0.02674f
C1459 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.10815f
C1460 sar10b_0.CF[6] sar10b_0.CF[3] 0.10965f
C1461 sar10b_0.SWN[3] EN 0.15924f
C1462 VSSA CLK 5.40882f
C1463 sar10b_0.SWN[1] sar10b_0.CF[3] 0.12225f
C1464 a_66101_58256# a_65966_58354# 0.35559f
C1465 m3_32416_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.33071f
C1466 m3_n1472_77772# VCM 0.01412f
C1467 VDDD a_68235_71265# 0.23014f
C1468 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR 0.95198f
C1469 c1_45456_23858# c1_45456_22738# 0.13255f
C1470 VDDD a_60693_51315# 0.33295f
C1471 a_60747_58903# sar10b_0.CF[2] 0.15195f
C1472 VDDD a_61493_67580# 0.20576f
C1473 sar10b_0.net16 sar10b_0.net41 1.45941f
C1474 VDDD a_66079_59638# 0.2054f
C1475 a_68421_65620# a_68767_65312# 0.07649f
C1476 sar10b_0.cyclic_flag_0.FINAL a_66933_65727# 0.0786f
C1477 sar10b_0.CF[4] VDDD 0.38234f
C1478 m3_45124_24938# m3_45124_23818# 0.29566f
C1479 sar10b_0._10_ a_67084_53565# 0.09174f
C1480 VSSR c1_n1140_51858# 0.04956f
C1481 a_67372_52833# sar10b_0.net35 0.03051f
C1482 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP sar10b_0.SWN[8] 0.18139f
C1483 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.07723f
C1484 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A VDDR 0.60027f
C1485 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 2.77549f
C1486 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A VDDR 0.60103f
C1487 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C1488 VDDD a_67733_54791# 0.21294f
C1489 sar10b_0.CF[5] VSSA 0.11644f
C1490 sar10b_0.clk_div_0.COUNT\[0\] sar10b_0.net16 0.13624f
C1491 m3_45124_94572# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C1492 sar10b_0.SWP[8] sar10b_0.net46 0.0472f
C1493 m3_29592_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.53894f
C1494 sar10b_0._08_ sar10b_0._02_ 0.13649f
C1495 m3_n1472_96812# m3_n1472_95692# 0.29566f
C1496 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y 0.32492f
C1497 a_61705_51992# sar10b_0.net1 0.01198f
C1498 m3_28180_21578# c1_28512_21618# 1.74381f
C1499 sar10b_0.net16 a_61737_56343# 0.1909f
C1500 m3_45124_31658# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C1501 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 0.21044f
C1502 sar10b_0.CF[1] VSSD 0.55164f
C1503 VSSD a_61677_62178# 0.13536f
C1504 m3_36652_97932# c1_36984_97972# 1.74381f
C1505 VSSR m3_n60_21578# 0.54178f
C1506 sar10b_0.net47 sar10b_0._06_ 0.18577f
C1507 sar10b_0.net46 a_66213_68756# 0.01005f
C1508 sar10b_0.net7 a_61153_51603# 0.01491f
C1509 sar10b_0.SWN[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 0.15996f
C1510 VDDD a_65857_56931# 0.22504f
C1511 c1_17216_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.28565f
C1512 a_68421_62956# a_68767_62648# 0.07649f
C1513 m3_22532_97932# th_dif_sw_0.VCP 0.01078f
C1514 sar10b_0.net34 sar10b_0.clknet_0_CLK 1.09676f
C1515 VSSD DATA[9] 0.7936f
C1516 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A sar10b_0.CF[3] 0.26294f
C1517 c1_24276_21618# th_dif_sw_0.VCN 0.13255f
C1518 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] a_15533_5779# 0.45291f
C1519 m3_45124_65452# m3_45124_64332# 0.29566f
C1520 a_n8277_54249# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 1.13669f
C1521 VSSR m3_45124_62092# 0.69778f
C1522 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.41774f
C1523 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 2.51837f
C1524 m3_19708_21578# VCM 0.13579f
C1525 m3_n1472_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C1526 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A 0.68875f
C1527 m3_n1472_81132# c1_n1140_81172# 1.74381f
C1528 m3_45124_82252# c1_45456_81172# 0.01078f
C1529 m3_45124_81132# c1_45456_82292# 0.01078f
C1530 c1_24276_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 0.01078f
C1531 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[2] 0.01887f
C1532 VDDA a_n4470_53722# 1.54446f
C1533 sar10b_0.SWP[4] VDDR 2.53551f
C1534 sar10b_0.SWN[2] a_33863_5788# 0.86021f
C1535 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_2868_8700# 0.01076f
C1536 VDDD a_64949_64916# 0.20573f
C1537 VDDD sar10b_0.clk_div_0.COUNT\[2\] 0.6004f
C1538 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[2] 0.17717f
C1539 a_29061_108738# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 0.70991f
C1540 c1_n1140_27218# m3_n1472_27178# 1.74381f
C1541 c1_45456_27218# m3_45124_28298# 0.01078f
C1542 c1_45456_28338# m3_45124_27178# 0.01078f
C1543 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C1544 w_n9655_56533# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 0.99238f
C1545 a_61395_52624# sar10b_0.net1 0.01311f
C1546 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 0.20503f
C1547 a_64085_60119# sar10b_0.net41 0.01157f
C1548 sar10b_0.net39 a_61419_71265# 0.09809f
C1549 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP sar10b_0.CF[2] 0.16026f
C1550 a_61589_53459# VSSD 0.09896f
C1551 sar10b_0.CF[1] sar10b_0.CF[8] 0.11291f
C1552 VSSA a_52417_59293# 0.14573f
C1553 c1_12980_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.26825f
C1554 VDDD sar10b_0.net30 0.81665f
C1555 sar10b_0.net8 a_62997_56643# 0.03741f
C1556 a_62181_58100# a_62527_58306# 0.07649f
C1557 a_61493_58256# a_61358_58354# 0.35559f
C1558 VDDD a_66865_49412# 0.39237f
C1559 VSSA th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 2.12202f
C1560 c1_45456_80052# VDDR 0.01153f
C1561 VDDA tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A 0.44525f
C1562 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.09687f
C1563 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR 4.47988f
C1564 VDDD a_61400_64952# 0.2536f
C1565 m3_22532_21578# m3_23944_21578# 0.23959f
C1566 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VCM 10.6522f
C1567 sar10b_0.net3 a_67297_55975# 0.10946f
C1568 VSSD a_66825_57675# 0.27918f
C1569 VSSR c1_45456_28338# 0.09348f
C1570 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSSR 6.45046f
C1571 VDDD a_67135_58306# 0.25389f
C1572 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 0.02632f
C1573 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[2] 0.01887f
C1574 a_66795_71265# sar10b_0.SWP[6] 0.1431f
C1575 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A a_45050_111636# 0.01076f
C1576 a_61803_48621# VSSD 0.29049f
C1577 m3_n1472_69932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C1578 sar10b_0.SWP[5] sar10b_0.SWP[6] 16.0927f
C1579 sar10b_0.clk_div_0.COUNT\[2\] sar10b_0._08_ 0.08449f
C1580 a_65682_49313# a_66368_49417# 0.27693f
C1581 a_65861_49313# a_66109_49318# 0.05308f
C1582 VSSR m3_35240_97932# 0.54637f
C1583 c1_n1140_66612# c1_n1140_65492# 0.13255f
C1584 VDDD VSSD 0.83276p
C1585 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26364f
C1586 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 0.24766f
C1587 m3_35240_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.53847f
C1588 a_61773_52237# sar10b_0.net1 0.02075f
C1589 m3_n1472_45098# VDDR 0.02681f
C1590 sar10b_0.net16 a_62313_61671# 0.19132f
C1591 a_61400_52964# a_61609_52946# 0.24088f
C1592 a_61395_52624# a_62185_52707# 0.1263f
C1593 m3_n1472_52938# VCM 0.01415f
C1594 sar10b_0.SWN[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A 0.01417f
C1595 a_61929_51311# sar10b_0.net16 0.27693f
C1596 VDDD a_67733_64115# 0.20863f
C1597 sar10b_0.net39 sar10b_0.net8 0.60018f
C1598 VDDD a_63561_60339# 0.83314f
C1599 VSSR c1_12980_97972# 0.05685f
C1600 a_55121_59650# a_55085_59917# 0.01114f
C1601 a_61589_50795# VSSD 0.09962f
C1602 sar10b_0.CF[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 0.12389f
C1603 sar10b_0.net16 a_64993_66255# 0.12529f
C1604 sar10b_0.clk_div_0.COUNT\[1\] a_67611_50645# 0.01819f
C1605 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_5588_21578# 0.03017f
C1606 c1_3096_21618# VCM 0.01358f
C1607 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VSSR 1.31843f
C1608 VDDD a_61400_60956# 0.2526f
C1609 a_63457_67583# a_63663_67678# 0.11249f
C1610 a_64492_67433# a_64238_67295# 0.28698f
C1611 a_61929_57971# sar10b_0.net4 0.08043f
C1612 a_61395_63280# a_60945_63273# 0.03471f
C1613 a_60747_63273# a_61086_63306# 0.07649f
C1614 sar10b_0.net42 sar10b_0.net11 0.0129f
C1615 sar10b_0.clk_div_0.COUNT\[0\] a_67696_52265# 0.18186f
C1616 m3_n1472_85612# VDDR 0.02674f
C1617 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[5] 0.05939f
C1618 sar10b_0.CF[4] sar10b_0.CF[2] 0.10792f
C1619 a_66027_53575# sar10b_0._10_ 0.0475f
C1620 sar10b_0.net38 a_61833_57675# 0.01363f
C1621 VDDD a_63295_55988# 0.2087f
C1622 m3_n1472_93452# VCM 0.01412f
C1623 a_61395_65944# a_61086_65970# 0.07766f
C1624 sar10b_0.clk_div_0.COUNT\[1\] sar10b_0.clk_div_0.COUNT\[0\] 1.31612f
C1625 sar10b_0._08_ VSSD 1.78237f
C1626 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] 21.6018f
C1627 sar10b_0.SWP[0] VCM 0.13076f
C1628 CLK a_52417_60961# 0.19115f
C1629 sar10b_0.SWP[2] sar10b_0.CF[9] 0.23628f
C1630 c1_45456_31698# c1_45456_30578# 0.13255f
C1631 VDDD sar10b_0.net20 0.73659f
C1632 a_67372_52833# a_67419_52937# 0.19021f
C1633 c1_32748_97972# VCM 0.01358f
C1634 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A 1.40448f
C1635 sar10b_0.net8 a_62037_61731# 0.05668f
C1636 m3_45124_32778# m3_45124_31658# 0.29566f
C1637 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A 0.03041f
C1638 VSSR c1_n1140_71092# 0.04956f
C1639 a_62187_71265# sar10b_0.SWP[2] 0.1431f
C1640 a_65573_52937# a_65682_51977# 0.01486f
C1641 m3_14060_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.31585f
C1642 c1_36984_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C1643 a_68767_67976# VSSD 0.26795f
C1644 a_62409_59007# sar10b_0.net4 0.02224f
C1645 a_67733_58787# sar10b_0.net3 0.16759f
C1646 a_60969_51311# a_61153_51603# 0.44532f
C1647 a_60690_53975# tdc_0.OUTN 0.02782f
C1648 VSSD DATA[6] 0.61076f
C1649 a_61153_67587# a_61358_67678# 0.09983f
C1650 a_62181_67424# a_61929_67295# 0.27388f
C1651 a_64910_59686# sar10b_0.net1 0.0683f
C1652 c1_14392_21618# m3_15472_21578# 0.15596f
C1653 a_60747_49953# sar10b_0.net29 0.2715f
C1654 m3_45124_47338# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C1655 VDDD sar10b_0.net31 1.4942f
C1656 VDDD sar10b_0.CF[8] 0.59652f
C1657 th_dif_sw_0.CKB EN 0.88994f
C1658 sar10b_0.net16 a_62702_61352# 0.2188f
C1659 sar10b_0.net2 sar10b_0.net43 0.03932f
C1660 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] th_dif_sw_0.VCN 8.84761f
C1661 CLK th_dif_sw_0.VCN 3.67999f
C1662 a_67445_60119# VSSD 0.09927f
C1663 m3_16884_97932# c1_17216_97972# 1.74381f
C1664 VSSR m3_45124_37258# 0.63261f
C1665 VSSA a_51861_60437# 0.01076f
C1666 m3_45124_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C1667 a_n4470_53722# th_dif_sw_0.CKB 0.77401f
C1668 sar10b_0._13_ sar10b_0._12_ 0.0113f
C1669 a_67419_52937# sar10b_0.net35 0.01512f
C1670 VSSR c1_31336_21618# 0.05685f
C1671 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y 0.31983f
C1672 a_67733_54791# a_68169_55011# 0.16939f
C1673 c1_22864_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.02548f
C1674 sar10b_0.CF[5] th_dif_sw_0.VCN 0.28582f
C1675 m3_45124_73292# m3_45124_72172# 0.29566f
C1676 VSSR m3_45124_77772# 0.63305f
C1677 VDDD a_61041_52340# 0.40229f
C1678 sar10b_0.net3 a_68421_54964# 0.17726f
C1679 a_62985_63003# sar10b_0.net16 0.16799f
C1680 a_61921_55975# a_62261_56123# 0.24088f
C1681 a_61737_56343# a_62697_56343# 0.03529f
C1682 sar10b_0.net8 a_62837_61451# 0.01222f
C1683 a_64188_51135# sar10b_0.clknet_1_0__leaf_CLK 0.2427f
C1684 sar10b_0.net9 sar10b_0.net39 0.09942f
C1685 sar10b_0.CF[6] sar10b_0.SWP[4] 0.12054f
C1686 sar10b_0.SWP[5] sar10b_0.CF[5] 2.41011f
C1687 m3_45124_90092# c1_45456_89012# 0.01078f
C1688 m3_45124_88972# c1_45456_90132# 0.01078f
C1689 m3_n1472_88972# c1_n1140_89012# 1.74381f
C1690 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A 0.03718f
C1691 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP a_19457_5788# 0.11862f
C1692 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VCM 0.12068f
C1693 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A 0.43728f
C1694 a_67393_54643# sar10b_0.net37 0.01277f
C1695 sar10b_0.net16 a_62185_64695# 0.22594f
C1696 sar10b_0.net32 sar10b_0.net40 0.02972f
C1697 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A 0.07183f
C1698 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A 0.01751f
C1699 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR 0.36439f
C1700 c1_n1140_35058# m3_n1472_35018# 1.74381f
C1701 c1_45456_36178# m3_45124_35018# 0.01078f
C1702 c1_45456_93492# c1_45456_94612# 0.13255f
C1703 c1_45456_35058# m3_45124_36138# 0.01078f
C1704 sar10b_0.clk_div_0.COUNT\[2\] sar10b_0._15_ 0.23043f
C1705 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A 0.39629f
C1706 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_26878_8700# 0.01076f
C1707 sar10b_0.SWN[9] sar10b_0.net36 0.05936f
C1708 m3_45124_62092# VDDR 0.01034f
C1709 sar10b_0.SWP[9] a_68946_71059# 0.14171f
C1710 VDDD a_68421_65620# 0.27523f
C1711 a_64521_60339# a_64773_60292# 0.27388f
C1712 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38377f
C1713 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.4143f
C1714 sar10b_0.net33 a_65397_56643# 0.01183f
C1715 sar10b_0._11_ sar10b_0._01_ 0.25543f
C1716 a_20335_112621# VSSR 1.79211f
C1717 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 3.46562f
C1718 a_65857_56931# a_66633_56639# 0.3578f
C1719 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 0.02632f
C1720 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.41774f
C1721 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 2.32591f
C1722 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSSR 2.47129f
C1723 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_12472_8700# 0.01076f
C1724 a_62593_58639# sar10b_0.net39 0.15044f
C1725 sar10b_0.CF[1] sar10b_0.SWN[0] 0.1215f
C1726 sar10b_0.net18 sar10b_0.net35 0.07915f
C1727 sar10b_0.net9 a_62037_61731# 0.03234f
C1728 VSSD a_68133_61624# 0.27171f
C1729 VSSD sar10b_0.CF[2] 0.78861f
C1730 c1_31336_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.26825f
C1731 m3_2764_21578# m3_4176_21578# 0.23959f
C1732 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.36778f
C1733 VSSR c1_45456_44018# 0.09348f
C1734 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A 0.45324f
C1735 sar10b_0.SWN[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.32591f
C1736 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VCM 0.12565f
C1737 sar10b_0.net16 a_62185_60699# 0.22647f
C1738 a_67598_58688# VSSD 0.13557f
C1739 m3_n1472_85612# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C1740 sar10b_0.net8 sar10b_0.net11 0.20344f
C1741 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP 5.97252f
C1742 c1_n1140_74452# c1_n1140_73332# 0.13255f
C1743 a_65407_63634# sar10b_0.net43 0.26926f
C1744 sar10b_0._15_ VSSD 0.56321f
C1745 sar10b_0.net16 sar10b_0.CF[7] 0.02393f
C1746 m3_39476_21578# c1_38396_21618# 0.15596f
C1747 sar10b_0.net32 a_64339_51661# 0.01289f
C1748 m3_n1472_22698# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C1749 sar10b_0.clknet_0_CLK sar10b_0._04_ 0.03387f
C1750 sar10b_0.clknet_1_1__leaf_CLK a_65861_51977# 0.01091f
C1751 a_61086_63306# VSSD 0.27173f
C1752 sar10b_0.SWP[4] sar10b_0.net41 0.04979f
C1753 c1_n1140_94612# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C1754 a_63273_56639# a_63797_56924# 0.05022f
C1755 VSSR m3_21120_21578# 0.34859f
C1756 VSSR a_44345_5779# 3.47951f
C1757 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR 0.96907f
C1758 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VDDR 2.42754f
C1759 th_dif_sw_0.VCN th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 0.09766f
C1760 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.41774f
C1761 c1_45456_28338# VDDR 0.01151f
C1762 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VDDR 3.77691f
C1763 m3_45124_31658# th_dif_sw_0.VCN 0.17339f
C1764 a_61493_51596# VSSD 0.0965f
C1765 a_62185_63363# sar10b_0.net4 0.03606f
C1766 a_62527_67630# VSSD 0.25983f
C1767 sar10b_0.net32 sar10b_0.net38 0.02875f
C1768 sar10b_0.net13 a_60693_67299# 0.21731f
C1769 VSSD a_64809_65963# 0.51846f
C1770 sar10b_0.SWP[4] a_25137_112201# 0.48461f
C1771 m3_43712_97932# th_dif_sw_0.VCP 0.01078f
C1772 sar10b_0.cyclic_flag_0.FINAL a_66933_68391# 0.05009f
C1773 m3_15472_97932# VCM 0.13579f
C1774 sar10b_0.net32 CLK 0.04119f
C1775 a_60945_52617# sar10b_0.net16 0.28151f
C1776 sar10b_0.net47 sar10b_0.net45 0.19839f
C1777 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_36984_21618# 0.0106f
C1778 a_68169_55011# VSSD 0.29076f
C1779 sar10b_0.net14 a_65769_65963# 0.03601f
C1780 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 1.76305f
C1781 c1_45456_39538# c1_45456_38418# 0.13255f
C1782 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN 8.05651f
C1783 VDDD a_64492_67433# 0.24883f
C1784 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[8] 0.05939f
C1785 a_61400_62288# a_62185_62031# 0.26257f
C1786 a_61609_62270# a_61677_62178# 0.35559f
C1787 sar10b_0.net4 a_60789_53739# 0.07102f
C1788 sar10b_0.net33 a_65761_58263# 0.01271f
C1789 m3_40888_21578# VCM 0.15231f
C1790 m3_19708_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C1791 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 sar10b_0.CF[2] 0.40679f
C1792 m3_45124_40618# m3_45124_39498# 0.29566f
C1793 a_64245_59307# sar10b_0.net1 0.21451f
C1794 sar10b_0.CF[3] sar10b_0.CF[7] 0.10897f
C1795 sar10b_0.CF[2] sar10b_0.CF[8] 0.10488f
C1796 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP 3.3819f
C1797 VSSR c1_n1140_86772# 0.04956f
C1798 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP sar10b_0.SWN[7] 0.2025f
C1799 sar10b_0._10_ a_64924_52385# 0.04086f
C1800 a_68421_64288# sar10b_0.net3 0.17732f
C1801 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VDDR 0.74911f
C1802 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP 5.18041f
C1803 sar10b_0.CF[4] VSSR 20.8404f
C1804 a_65119_59984# VSSD 0.2614f
C1805 VSSD a_66633_56639# 0.28526f
C1806 a_64609_64923# a_64814_65014# 0.09983f
C1807 a_60690_54641# sar10b_0.net1 0.24179f
C1808 a_65637_64760# a_65385_64631# 0.27388f
C1809 sar10b_0.net40 a_65589_57735# 0.0448f
C1810 sar10b_0.clk_div_0.COUNT\[0\] sar10b_0._07_ 0.16703f
C1811 a_61803_48621# sar10b_0.SWN[0] 0.14362f
C1812 VDDD a_64543_62648# 0.2037f
C1813 VDDD sar10b_0.SWN[0] 0.63674f
C1814 VSSR m3_45124_52938# 0.63261f
C1815 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A 0.28117f
C1816 a_66933_68391# a_67393_67963# 0.26257f
C1817 a_67209_68331# a_67598_68012# 0.05462f
C1818 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A 0.83476f
C1819 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] VCM 16.1243f
C1820 c1_n1140_29458# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C1821 sar10b_0.net9 a_62709_63063# 0.03378f
C1822 sar10b_0.net16 a_61395_65944# 0.19058f
C1823 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.24766f
C1824 m3_5588_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C1825 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45324f
C1826 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 4.15629f
C1827 a_68562_48647# VSSD 0.29268f
C1828 a_64425_64631# sar10b_0.net11 0.22485f
C1829 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.09687f
C1830 VSSR c1_4508_21618# 0.05923f
C1831 sar10b_0.SWP[8] CKO 0.8498f
C1832 sar10b_0.net32 a_64491_48621# 0.26661f
C1833 sar10b_0.CF[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 0.10431f
C1834 sar10b_0.net9 sar10b_0.net11 0.18612f
C1835 a_63810_50901# a_64199_50761# 0.06302f
C1836 m3_45124_62092# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C1837 a_62025_53679# sar10b_0.net1 0.03515f
C1838 a_67371_49579# a_68562_49747# 0.01073f
C1839 m3_45124_81132# m3_45124_80012# 0.29566f
C1840 VSSR m3_45124_93452# 0.63305f
C1841 sar10b_0.net4 a_63273_67295# 0.22606f
C1842 a_65983_64966# VSSD 0.26586f
C1843 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_46086_111642# 0.01076f
C1844 m3_45124_37258# VDDR 0.0103f
C1845 a_65525_68912# sar10b_0.net16 0.17488f
C1846 VSSR cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 94.3862f
C1847 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 0.19757f
C1848 a_65394_52643# a_65573_52937# 0.54361f
C1849 a_65577_57971# VSSD 0.5498f
C1850 VCM sar10b_0.SWP[1] 0.13076f
C1851 a_61400_64952# a_61677_64842# 0.09983f
C1852 VSSR c1_34160_97972# 0.05923f
C1853 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A 1.31843f
C1854 sar10b_0._04_ a_68178_51635# 0.09393f
C1855 sar10b_0.cyclic_flag_0.FINAL a_66645_61731# 0.04985f
C1856 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C1857 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A 0.11547f
C1858 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_26768_21578# 0.03017f
C1859 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_9824_21578# 0.0162f
C1860 a_68946_49747# VSSD 0.29465f
C1861 a_61491_52222# a_60969_51311# 0.12076f
C1862 sar10b_0.clknet_0_CLK a_66593_50645# 0.01318f
C1863 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VSSR 1.3401f
C1864 c1_n1140_42898# m3_n1472_42858# 1.74381f
C1865 c1_45456_42898# m3_45124_43978# 0.01078f
C1866 c1_45456_44018# m3_45124_42858# 0.01078f
C1867 VDDD a_61400_50300# 0.24576f
C1868 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN sar10b_0.SWN[5] 0.2156f
C1869 VSSD a_61677_64842# 0.13539f
C1870 a_67696_52265# sar10b_0._03_ 0.22746f
C1871 m3_45124_77772# VDDR 0.01034f
C1872 m3_45124_74412# th_dif_sw_0.VCP 0.17339f
C1873 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 0.02632f
C1874 VDDD a_61609_62270# 0.2082f
C1875 m3_14060_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.54821f
C1876 sar10b_0.net5 a_60747_56239# 0.26268f
C1877 sar10b_0.clk_div_0.COUNT\[1\] sar10b_0._03_ 0.55713f
C1878 a_61153_58263# sar10b_0.net1 0.02102f
C1879 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP sar10b_0.CF[7] 0.10502f
C1880 a_62025_51015# sar10b_0.net1 0.03088f
C1881 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A sar10b_0.CF[7] 0.06369f
C1882 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A 0.28117f
C1883 a_63621_58960# VSSD 0.26751f
C1884 VDDD a_61677_66174# 0.2729f
C1885 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VCM 3.00607f
C1886 a_65778_49979# a_66205_50408# 0.04602f
C1887 sar10b_0._02_ a_65485_50273# 0.01649f
C1888 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A 0.38397f
C1889 a_n8277_54565# th_dif_sw_0.th_sw_1.CKB 0.03405f
C1890 m3_45124_65452# c1_45456_65492# 1.74381f
C1891 m3_n1472_64332# c1_n1140_65492# 0.01078f
C1892 m3_n1472_65452# c1_n1140_64372# 0.01078f
C1893 a_64809_63299# sar10b_0.net12 0.03114f
C1894 VSSR c1_45456_63252# 0.0935f
C1895 sar10b_0.net19 a_68767_54656# 0.02268f
C1896 a_68169_64335# VSSD 0.29048f
C1897 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR 0.59908f
C1898 VSSD tdc_0.OUTN 0.89784f
C1899 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A 0.60027f
C1900 sar10b_0.net13 a_65769_65963# 0.013f
C1901 a_65865_69663# VSSD 0.50051f
C1902 a_38665_5788# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.92132f
C1903 m3_35240_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.53847f
C1904 m3_11236_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.53633f
C1905 m3_38064_97932# m3_39476_97932# 0.23959f
C1906 a_67733_64115# a_68169_64335# 0.16939f
C1907 c1_n1140_82292# c1_n1140_81172# 0.13255f
C1908 a_61454_53360# a_61589_53459# 0.35559f
C1909 m3_n1472_38378# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C1910 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38781f
C1911 m3_21120_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.07708f
C1912 VSSD a_61677_60846# 0.12188f
C1913 VCM cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 2.92973f
C1914 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A 0.43773f
C1915 sar10b_0.cyclic_flag_0.FINAL a_67209_55011# 0.23275f
C1916 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38377f
C1917 th_dif_sw_0.CK VCM 0.25227f
C1918 a_60969_56639# a_61493_56924# 0.05022f
C1919 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VDDR 2.82798f
C1920 VSSR VSSD 0.14702f
C1921 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VSSR 2.35116f
C1922 a_51603_58977# a_51345_58977# 0.06738f
C1923 m3_28180_97932# c1_27100_97972# 0.15596f
C1924 VSSR m3_n1472_28298# 0.66371f
C1925 sar10b_0.net19 sar10b_0.net37 0.45667f
C1926 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 32.8146f
C1927 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.59327f
C1928 a_66933_67059# a_67598_66680# 0.19065f
C1929 a_67209_66999# a_67733_66779# 0.04522f
C1930 c1_45456_44018# VDDR 0.01151f
C1931 m3_45124_47338# th_dif_sw_0.VCN 0.17339f
C1932 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 sar10b_0.CF[0] 0.26334f
C1933 sar10b_0.net46 a_66795_71265# 0.07022f
C1934 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A sar10b_0.CF[7] 0.26294f
C1935 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP 7.39379f
C1936 a_61400_60956# a_61677_60846# 0.09983f
C1937 VDDD a_61454_53360# 0.27686f
C1938 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VSSR 4.77312f
C1939 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_10156_21618# 0.0106f
C1940 c1_18628_21618# th_dif_sw_0.VCN 0.13255f
C1941 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 4.15627f
C1942 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 0.21775f
C1943 sar10b_0.net1 a_61461_56403# 0.01427f
C1944 VSSR m3_n1472_68812# 0.66316f
C1945 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A 1.37552f
C1946 c1_45456_47378# c1_45456_46258# 0.13255f
C1947 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y VSSR 0.32296f
C1948 sar10b_0.clknet_1_0__leaf_CLK a_65765_50645# 0.02212f
C1949 a_60747_52617# VSSD 0.26212f
C1950 sar10b_0.net32 a_63457_56931# 0.01355f
C1951 m3_1352_21578# VCM 0.15231f
C1952 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38377f
C1953 c1_n1140_71092# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C1954 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A sar10b_0.CF[5] 0.06369f
C1955 m3_45124_48458# m3_45124_47338# 0.29566f
C1956 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A 1.40448f
C1957 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.20752f
C1958 sar10b_0._00_ a_64761_51028# 0.12121f
C1959 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 4.02253f
C1960 sar10b_0.net38 a_66062_57022# 0.0468f
C1961 VDDD a_61419_48621# 0.23485f
C1962 sar10b_0.SWN[0] sar10b_0.CF[2] 0.12301f
C1963 tdc_0.RDY sar10b_0.net5 0.50539f
C1964 sar10b_0.cyclic_flag_0.FINAL sar10b_0.net35 1.07687f
C1965 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A 0.68875f
C1966 sar10b_0.net4 a_61609_52946# 0.02747f
C1967 VSSA a_51861_59345# 0.01076f
C1968 VDDD a_64238_63682# 0.25631f
C1969 a_65643_48621# VSSD 0.33428f
C1970 sar10b_0.net1 a_62997_56643# 0.17079f
C1971 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.41934f
C1972 m3_n1472_57418# VCM 0.01415f
C1973 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN 4.85899f
C1974 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 3.28979f
C1975 a_68169_66999# a_68767_66644# 0.06623f
C1976 VSSR sar10b_0.CF[8] 25.1643f
C1977 VDDD a_61454_50696# 0.27534f
C1978 sar10b_0.net10 a_63169_62635# 0.05797f
C1979 c1_n1140_45138# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C1980 a_61496_52091# VSSD 0.84834f
C1981 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP 6.18181f
C1982 sar10b_0.CF[4] VDDR 1.72081f
C1983 a_66921_61671# a_67105_61303# 0.44098f
C1984 VSSD a_63391_57320# 0.25378f
C1985 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR 0.41429f
C1986 VSSR c1_n1140_35058# 0.04956f
C1987 a_61454_50696# a_61589_50795# 0.35559f
C1988 a_61065_51015# a_62277_50968# 0.07766f
C1989 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C1990 sar10b_0.net16 a_62185_50043# 0.22144f
C1991 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A 0.28117f
C1992 m3_45124_77772# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C1993 sar10b_0.net14 a_65589_57735# 0.0183f
C1994 m3_45124_88972# m3_45124_87852# 0.29566f
C1995 sar10b_0.net38 sar10b_0.net40 0.38378f
C1996 VSSR m3_16884_97932# 0.43913f
C1997 m3_16884_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26806f
C1998 m3_45124_52938# VDDR 0.0103f
C1999 sar10b_0.net39 sar10b_0.net1 0.11968f
C2000 sar10b_0.net7 a_60693_57975# 0.18483f
C2001 VDDD sar10b_0.clknet_0_CLK 3.01735f
C2002 VSSR m3_42300_21578# 0.54637f
C2003 a_64521_59303# sar10b_0.net16 0.18721f
C2004 a_65001_68627# VSSD 0.50973f
C2005 VCM cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 3.63692f
C2006 a_68235_71265# sar10b_0.SWP[7] 0.14231f
C2007 a_67209_63003# sar10b_0.net3 0.19165f
C2008 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.96901f
C2009 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 7.63331f
C2010 VDDD a_68421_68284# 0.27537f
C2011 a_64809_63299# sar10b_0.net41 0.0257f
C2012 sar10b_0.net39 a_61400_66284# 0.01673f
C2013 sar10b_0._06_ a_67890_69727# 0.2612f
C2014 c1_n1140_50738# m3_n1472_50698# 1.74381f
C2015 c1_45456_51858# m3_45124_50698# 0.01078f
C2016 c1_45456_50738# m3_45124_51818# 0.01078f
C2017 c1_45456_97972# c1_45456_96852# 0.13255f
C2018 sar10b_0.net33 a_65765_50645# 0.02734f
C2019 sar10b_0.SWP[4] sar10b_0.CF[7] 0.12409f
C2020 VSSR a_9853_112162# 0.06033f
C2021 m3_45124_90092# th_dif_sw_0.VCP 0.17339f
C2022 m3_45124_93452# VDDR 0.01034f
C2023 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS a_n9133_57045# 1.06244f
C2024 VDDD a_67310_60020# 0.30248f
C2025 sar10b_0.CF[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.40692f
C2026 m3_36652_97932# VCM 0.15231f
C2027 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 0.12068f
C2028 VDDR cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 12.9105f
C2029 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 0.19259f
C2030 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.36333f
C2031 sar10b_0.net3 a_67733_66779# 0.16771f
C2032 sar10b_0.clknet_0_CLK sar10b_0._08_ 0.85465f
C2033 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A 0.74911f
C2034 sar10b_0.clk_div_0.COUNT\[0\] a_66762_50329# 0.06634f
C2035 sar10b_0.SWN[3] sar10b_0.CF[9] 0.20114f
C2036 c1_14392_97972# VCM 0.01358f
C2037 m3_40888_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C2038 m3_45124_73292# c1_45456_73332# 1.74381f
C2039 m3_n1472_73292# c1_n1140_72212# 0.01078f
C2040 m3_n1472_72172# c1_n1140_73332# 0.01078f
C2041 VSSR c1_45456_78932# 0.0935f
C2042 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP a_5051_5788# 0.04592f
C2043 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VDDR 0.76083f
C2044 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN sar10b_0.CF[0] 0.12404f
C2045 a_64339_51661# CLK 0.01475f
C2046 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 0.24779f
C2047 m3_26768_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.33071f
C2048 VSSR a_15533_113041# 1.45369f
C2049 sar10b_0.net46 a_66389_69443# 0.02773f
C2050 c1_18628_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C2051 a_65355_53949# sar10b_0.clknet_1_1__leaf_CLK 1.83449f
C2052 m3_18296_97932# m3_19708_97932# 0.23959f
C2053 a_62277_53632# sar10b_0.net16 0.17424f
C2054 c1_n1140_90132# c1_n1140_89012# 0.13255f
C2055 c1_5920_21618# m3_5588_21578# 1.74381f
C2056 a_65525_68912# a_65390_69010# 0.35559f
C2057 VDDD sar10b_0.SWN[8] 0.1348f
C2058 m3_n1472_54058# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C2059 a_64521_59303# a_65733_59432# 0.07766f
C2060 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 0.02632f
C2061 VDDD a_68767_62648# 0.2142f
C2062 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A sar10b_0.CF[4] 0.03041f
C2063 m3_8412_97932# c1_7332_97972# 0.15596f
C2064 VSSR m3_n1472_43978# 0.66371f
C2065 a_68421_68284# a_68767_67976# 0.07649f
C2066 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 2.62172f
C2067 sar10b_0._10_ a_64818_49979# 0.0141f
C2068 c1_272_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26825f
C2069 a_61182_52404# a_61491_52222# 0.07766f
C2070 a_61041_52340# a_61496_52091# 0.3578f
C2071 sar10b_0.net38 a_66933_55071# 0.1762f
C2072 c1_45456_63252# VDDR 0.01153f
C2073 sar10b_0.SWP[0] a_44345_110521# 0.79636f
C2074 m3_26768_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C2075 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 a_39543_5779# 0.67311f
C2076 sar10b_0.SWN[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP 0.32961f
C2077 VSSD a_63663_67678# 0.15049f
C2078 a_63169_62635# a_63509_62783# 0.24088f
C2079 a_62985_63003# a_63945_63003# 0.03529f
C2080 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A sar10b_0.CF[2] 0.03041f
C2081 m3_43712_21578# m3_45124_21578# 0.23959f
C2082 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 1.80961f
C2083 a_n8277_54249# a_n8277_54565# 0.64152f
C2084 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 2.76716f
C2085 a_62793_57675# a_63045_57628# 0.27388f
C2086 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A 0.45324f
C2087 VDDD sar10b_0.SWN[9] 0.67918f
C2088 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A 0.38472f
C2089 VSSR m3_n1472_84492# 0.66316f
C2090 a_61493_58256# sar10b_0.net16 0.147f
C2091 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 0.39671f
C2092 a_67310_60020# a_67445_60119# 0.35559f
C2093 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A sar10b_0.CF[1] 0.06369f
C2094 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 2.62169f
C2095 c1_45456_55218# c1_45456_54098# 0.13255f
C2096 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VDDR 2.58955f
C2097 sar10b_0.net30 sar10b_0.net17 0.08434f
C2098 m3_n1472_28298# VDDR 0.02681f
C2099 VDDD a_67881_61671# 0.36642f
C2100 a_62277_50968# sar10b_0.net16 0.17886f
C2101 m3_n1472_36138# VCM 0.01415f
C2102 c1_n1140_86772# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C2103 m3_45124_56298# m3_45124_55178# 0.29566f
C2104 sar10b_0.CF[5] CLK 0.0933f
C2105 VDDD a_67393_58639# 0.24874f
C2106 VDDA sar10b_0.CF[9] 2.12323f
C2107 a_62133_59067# sar10b_0.net40 0.02291f
C2108 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_31004_21578# 0.0162f
C2109 sar10b_0.net32 a_64428_50947# 0.02444f
C2110 VDDD a_68178_51635# 0.48266f
C2111 w_n9655_56533# a_n8277_54565# 0.05534f
C2112 c1_32748_21618# VCM 0.01358f
C2113 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VDDR 5.56107f
C2114 VDDD a_60945_63273# 0.40821f
C2115 a_67113_56343# a_67502_56024# 0.05462f
C2116 a_66837_56403# a_67297_55975# 0.26257f
C2117 sar10b_0.net14 sar10b_0.net40 0.20589f
C2118 m3_n1472_68812# VDDR 0.02674f
C2119 th_dif_sw_0.CK w_n9655_63119# 0.0364f
C2120 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VDDR 0.83965f
C2121 sar10b_0.net17 VSSD 1.22632f
C2122 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP 0.02666f
C2123 sar10b_0.net10 a_63849_63299# 0.22494f
C2124 m3_n1472_76652# VCM 0.01412f
C2125 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y VDDR 0.31995f
C2126 a_n8277_54565# VSSA 3.41647f
C2127 c1_n1140_22738# c1_n1140_21618# 0.13255f
C2128 VSSD a_67598_66680# 0.13557f
C2129 sar10b_0.CF[6] sar10b_0.CF[4] 0.11629f
C2130 VDDA VINN 0.87608f
C2131 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VDDR 0.83476f
C2132 VDDD a_61153_51603# 0.25172f
C2133 VDDD a_61929_67295# 0.35681f
C2134 sar10b_0.CF[4] sar10b_0.SWN[1] 0.12243f
C2135 VSSD sar10b_0.SWP[7] 0.94977f
C2136 a_64949_64916# sar10b_0.net12 0.02022f
C2137 VSSR sar10b_0.SWN[0] 7.20022f
C2138 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VCM 0.59215f
C2139 c1_12980_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.26825f
C2140 sar10b_0.cyclic_flag_0.FINAL a_67393_65299# 0.07652f
C2141 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y VSSR 0.32296f
C2142 VDDD a_64533_65967# 0.29488f
C2143 m3_n1472_23818# m3_n1472_22698# 0.29566f
C2144 sar10b_0._10_ sar10b_0._16_ 0.12593f
C2145 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 1.14734f
C2146 VSSR c1_n1140_50738# 0.04956f
C2147 sar10b_0.net1 sar10b_0.net11 0.74446f
C2148 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A a_39543_5779# 0.01247f
C2149 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM 0.99611f
C2150 sar10b_0.clk_div_0.COUNT\[1\] sar10b_0._13_ 0.02357f
C2151 tdc_0.RDY sar10b_0.net7 0.42734f
C2152 sar10b_0._08_ a_68178_51635# 0.04009f
C2153 m3_45124_93452# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C2154 sar10b_0.cyclic_flag_0.FINAL sar10b_0.net44 1.08798f
C2155 m3_32416_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.33071f
C2156 m3_45124_96812# m3_45124_95692# 0.29566f
C2157 m3_29592_21578# c1_29924_21618# 1.74381f
C2158 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.43221f
C2159 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 2.6566f
C2160 sar10b_0.net33 a_66049_57307# 0.0259f
C2161 m3_45124_30538# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C2162 th_dif_sw_0.VCN a_51861_59345# 0.06955f
C2163 VDDR sar10b_0.CF[8] 1.75928f
C2164 a_61677_50190# VSSD 0.13649f
C2165 c1_34160_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26825f
C2166 a_66049_69295# a_67077_69616# 0.07826f
C2167 VSSD a_62185_62031# 0.15425f
C2168 m3_38064_97932# c1_38396_97972# 1.74381f
C2169 VSSR m3_2764_21578# 0.54637f
C2170 sar10b_0.net6 a_61737_56343# 0.23202f
C2171 sar10b_0.net46 a_66559_68962# 0.28941f
C2172 VDDD a_64773_60292# 0.26785f
C2173 c1_20040_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.01445f
C2174 VDDD a_66885_56768# 0.29585f
C2175 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR 0.38768f
C2176 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] VCM 16.1243f
C2177 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN 6.85522f
C2178 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C2179 VSSD sar10b_0.net12 3.04889f
C2180 sar10b_0.net3 a_65068_49569# 0.12376f
C2181 a_65643_71265# sar10b_0.net43 0.30172f
C2182 sar10b_0.net2 a_65589_69723# 0.16776f
C2183 CLK a_52417_59293# 0.19115f
C2184 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 0.53683f
C2185 sar10b_0.clk_div_0.COUNT\[0\] sar10b_0._02_ 0.0764f
C2186 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] th_dif_sw_0.VCN 0.55567p
C2187 sar10b_0.net34 sar10b_0.clknet_1_1__leaf_CLK 0.06387f
C2188 sar10b_0.net17 sar10b_0.net31 0.48832f
C2189 m3_22532_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 0.24105f
C2190 sar10b_0.net38 sar10b_0.net14 0.05463f
C2191 sar10b_0.net16 a_63273_56639# 0.17903f
C2192 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A 0.28117f
C2193 c1_27100_21618# th_dif_sw_0.VCN 0.13255f
C2194 m3_n1472_64332# m3_n1472_63212# 0.29566f
C2195 VINP th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 0.36273f
C2196 a_63339_48621# sar10b_0.SWN[3] 0.15514f
C2197 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.45324f
C2198 a_51603_58977# VDDA 0.01057f
C2199 a_65573_52937# VSSD 0.59628f
C2200 VDDD a_68235_48621# 0.22633f
C2201 sar10b_0.CF[8] sar10b_0.SWP[7] 0.12093f
C2202 sar10b_0._06_ sar10b_0.net27 0.01028f
C2203 m3_22532_21578# VCM 0.11203f
C2204 m3_1352_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C2205 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 4.5807f
C2206 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] sar10b_0.CF[9] 0.01482f
C2207 m3_n1472_80012# c1_n1140_81172# 0.01078f
C2208 m3_45124_81132# c1_45456_81172# 1.74381f
C2209 m3_n1472_81132# c1_n1140_80052# 0.01078f
C2210 th_dif_sw_0.VCP th_dif_sw_0.th_sw_1.CKB 0.25482f
C2211 a_66865_52076# sar10b_0.net35 0.03098f
C2212 VDDR a_9853_112162# 2.42521f
C2213 VSSD a_63662_57022# 0.13881f
C2214 m3_n1472_97932# m3_n60_97932# 0.23959f
C2215 VDDD a_65385_64631# 0.36326f
C2216 c1_45456_27218# m3_45124_27178# 1.74381f
C2217 c1_n1140_26098# m3_n1472_27178# 0.01078f
C2218 c1_n1140_27218# m3_n1472_26058# 0.01078f
C2219 sar10b_0.clknet_1_0__leaf_CLK sar10b_0.net16 0.06422f
C2220 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 0.22396f
C2221 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 0.24771f
C2222 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 8.70956f
C2223 VDDD a_65301_57975# 0.30137f
C2224 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.59833f
C2225 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A 0.42509f
C2226 c1_15804_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.01532f
C2227 a_67881_60339# sar10b_0.net3 0.29276f
C2228 sar10b_0.SWP[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 0.25013f
C2229 VDDD a_68562_49747# 0.25277f
C2230 c1_45456_22738# c1_45456_21618# 0.13255f
C2231 sar10b_0.net10 sar10b_0.net40 0.02564f
C2232 c1_45456_78932# VDDR 0.01153f
C2233 th_dif_sw_0.CKB sar10b_0.CF[9] 4.43166f
C2234 VSSD DATA[0] 0.98421f
C2235 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y VSSR 0.32296f
C2236 sar10b_0.net13 sar10b_0.net40 0.03114f
C2237 a_67881_61671# a_68133_61624# 0.27388f
C2238 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 0.19259f
C2239 VDDD a_61609_64934# 0.20839f
C2240 m3_23944_21578# m3_25356_21578# 0.23959f
C2241 sar10b_0.net3 a_67637_56123# 0.16877f
C2242 VSSD a_67423_57320# 0.26819f
C2243 sar10b_0.net38 a_63457_56931# 0.01247f
C2244 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] th_dif_sw_0.VCN 0.13856p
C2245 VSSR c1_45456_27218# 0.09348f
C2246 a_63810_50901# a_64188_51135# 0.0649f
C2247 sar10b_0.CF[6] VSSD 0.77503f
C2248 a_61677_63510# sar10b_0.net16 0.31615f
C2249 a_66933_59067# sar10b_0.net39 0.1793f
C2250 m3_n1472_68812# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C2251 sar10b_0.SWN[1] VSSD 1.02169f
C2252 VSSR a_38665_5788# 0.06033f
C2253 a_65861_49313# a_66216_49358# 0.18752f
C2254 VSSR m3_38064_97932# 0.54637f
C2255 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 0.32628f
C2256 sar10b_0.SWP[7] a_9853_112162# 0.33169f
C2257 c1_45456_66612# c1_45456_65492# 0.13255f
C2258 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A sar10b_0.CF[2] 0.02149f
C2259 VDDD a_63369_59007# 0.37108f
C2260 VSSA a_53564_60302# 0.02937f
C2261 m3_38064_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.53746f
C2262 sar10b_0.net3 sar10b_0._10_ 0.08617f
C2263 m3_n1472_43978# VDDR 0.02681f
C2264 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.95009f
C2265 m3_n1472_51818# VCM 0.01415f
C2266 sar10b_0.net46 sar10b_0.SWP[6] 0.04776f
C2267 a_67393_58639# a_67598_58688# 0.09983f
C2268 a_67209_59007# a_68169_59007# 0.03529f
C2269 a_60969_57971# VSSD 0.51115f
C2270 sar10b_0.net28 sar10b_0.net16 0.3364f
C2271 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.39559f
C2272 VSSR c1_15804_97972# 0.06681f
C2273 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] a_249_5788# 0.28719f
C2274 a_55121_59650# tdc_0.RDY 0.14294f
C2275 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 0.21212f
C2276 sar10b_0.net16 a_66021_66092# 0.17391f
C2277 a_60690_49683# VSSD 0.95563f
C2278 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_8412_21578# 0.03017f
C2279 VDDD sar10b_0.net47 1.39471f
C2280 sar10b_0.SWP[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.02059f
C2281 a_61153_67587# sar10b_0.net39 0.01979f
C2282 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.11339f
C2283 c1_5920_21618# VCM 0.01358f
C2284 a_68178_51635# sar10b_0._15_ 0.0207f
C2285 sar10b_0.net31 a_63662_57022# 0.03138f
C2286 VDDD a_61609_60938# 0.20831f
C2287 a_64238_67295# a_64888_67630# 0.07298f
C2288 a_61358_58354# sar10b_0.net4 0.07118f
C2289 a_61395_63280# a_61400_63620# 0.44098f
C2290 a_60945_63273# a_61086_63306# 0.27388f
C2291 m3_n1472_84492# VDDR 0.02674f
C2292 sar10b_0.clk_div_0.COUNT\[0\] sar10b_0.clk_div_0.COUNT\[2\] 0.85964f
C2293 m3_n1472_92332# VCM 0.01412f
C2294 DATA[4] a_68946_56639# 0.14366f
C2295 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 1.73977f
C2296 CLK a_51861_60437# 0.01174f
C2297 c1_n1140_30578# c1_n1140_29458# 0.13255f
C2298 sar10b_0._01_ a_65188_51977# 0.05333f
C2299 sar10b_0.net3 sar10b_0.net39 0.13353f
C2300 sar10b_0.clk_div_0.COUNT\[0\] a_66865_49412# 0.121f
C2301 c1_35572_97972# VCM 0.01358f
C2302 sar10b_0._03_ a_66762_50329# 0.04284f
C2303 sar10b_0.net10 sar10b_0.net38 0.05981f
C2304 sar10b_0.net33 sar10b_0.net16 0.77742f
C2305 m3_n1472_31658# m3_n1472_30538# 0.29566f
C2306 tdc_0.RDY tdc_0.OUTP 0.78763f
C2307 VSSR c1_n1140_69972# 0.04956f
C2308 sar10b_0.net38 sar10b_0.net13 0.02538f
C2309 sar10b_0.net41 VSSD 3.07089f
C2310 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 sar10b_0.SWN[7] 0.38458f
C2311 m3_16884_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26806f
C2312 a_66080_53027# a_65861_51977# 0.01198f
C2313 sar10b_0.CF[6] sar10b_0.CF[8] 0.1211f
C2314 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 2.77569f
C2315 c1_39808_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C2316 a_60969_51311# a_62181_51440# 0.07766f
C2317 a_61153_51603# a_61493_51596# 0.24088f
C2318 sar10b_0.SWN[1] sar10b_0.CF[8] 0.13825f
C2319 a_61929_67295# a_62527_67630# 0.06623f
C2320 c1_15804_21618# m3_16884_21578# 0.15596f
C2321 m3_45124_46218# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C2322 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 sar10b_0.CF[8] 0.26243f
C2323 sar10b_0.clk_div_0.COUNT\[0\] VSSD 1.70912f
C2324 sar10b_0.SWN[2] VSSA 0.24827f
C2325 m3_18296_97932# c1_18628_97972# 1.74381f
C2326 VSSD a_61737_56343# 0.54914f
C2327 a_64533_65967# a_64809_65963# 0.1263f
C2328 VDDR sar10b_0.SWN[0] 3.77806f
C2329 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A 0.68875f
C2330 VSSR m3_45124_36138# 0.63261f
C2331 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y VDDR 0.31995f
C2332 sar10b_0.net3 a_67209_65667# 0.17888f
C2333 a_66593_50645# a_66785_50875# 0.33658f
C2334 a_44345_110521# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A 0.01247f
C2335 sar10b_0.CF[5] sar10b_0.net10 0.01296f
C2336 a_67502_56024# VSSD 0.13717f
C2337 sar10b_0.net4 a_61395_60616# 0.21755f
C2338 VSSR c1_34160_21618# 0.05923f
C2339 VDDA tdc_0.phase_detector_0.pd_out_0.B 1.23572f
C2340 a_41284_8700# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01076f
C2341 a_65865_57675# a_66049_57307# 0.44098f
C2342 th_dif_sw_0.VCP sar10b_0.CF[0] 0.2858f
C2343 m3_n1472_72172# m3_n1472_71052# 0.29566f
C2344 VSSR m3_45124_76652# 0.63305f
C2345 sar10b_0.net33 a_65733_59432# 0.01049f
C2346 VDDD a_61491_52222# 0.78542f
C2347 a_68479_59984# sar10b_0.net21 0.26912f
C2348 sar10b_0.net17 sar10b_0.SWN[0] 0.17327f
C2349 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 0.64443f
C2350 sar10b_0.SWP[3] a_29061_108738# 0.75451f
C2351 VDDD a_63045_57628# 0.26987f
C2352 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 sar10b_0.CF[9] 0.26243f
C2353 sar10b_0._01_ a_65765_50645# 0.28699f
C2354 m3_n1472_88972# c1_n1140_87892# 0.01078f
C2355 m3_45124_88972# c1_45456_89012# 1.74381f
C2356 m3_n1472_87852# c1_n1140_89012# 0.01078f
C2357 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN 4.04975f
C2358 a_68946_49747# sar10b_0.SWN[9] 0.14513f
C2359 a_65682_51977# a_66368_52081# 0.27693f
C2360 a_65861_51977# a_66109_51982# 0.05308f
C2361 c1_45456_35058# m3_45124_35018# 1.74381f
C2362 sar10b_0.CF[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17717f
C2363 c1_n1140_33938# m3_n1472_35018# 0.01078f
C2364 c1_n1140_35058# m3_n1472_33898# 0.01078f
C2365 a_68073_56343# a_68671_55988# 0.06623f
C2366 a_62281_52347# sar10b_0.net16 0.29423f
C2367 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSSR 5.64423f
C2368 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 4.92029f
C2369 a_64773_60292# a_65119_59984# 0.07649f
C2370 VSSR sar10b_0.SWN[8] 3.60822f
C2371 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 2.76888f
C2372 a_63849_63299# a_64033_63591# 0.44532f
C2373 a_66885_56768# a_66633_56639# 0.27388f
C2374 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 31.0559f
C2375 a_61035_71265# VSSD 0.31069f
C2376 a_64454_51311# a_64199_50761# 0.01197f
C2377 a_62933_58787# sar10b_0.net39 0.07776f
C2378 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A 0.68875f
C2379 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 sar10b_0.CF[7] 0.26243f
C2380 VSSD a_68946_61735# 0.33464f
C2381 sar10b_0.SWN[4] a_24259_5788# 0.64881f
C2382 sar10b_0._12_ sar10b_0.net35 0.02546f
C2383 a_66254_69344# sar10b_0.net16 0.22699f
C2384 m3_4176_21578# m3_5588_21578# 0.23959f
C2385 sar10b_0.net33 sar10b_0._17_ 0.0251f
C2386 sar10b_0.net40 a_61395_61948# 0.01467f
C2387 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A sar10b_0.CF[8] 0.26294f
C2388 VSSR c1_45456_42898# 0.09348f
C2389 VDDD sar10b_0.net43 1.72453f
C2390 m3_n1472_84492# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C2391 a_60690_54641# sar10b_0.net5 0.01943f
C2392 a_66464_50363# a_66762_50329# 0.02614f
C2393 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C2394 VSSR m3_n1472_97932# 0.71177f
C2395 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 2.53489f
C2396 c1_45456_74452# c1_45456_73332# 0.13255f
C2397 m3_40888_21578# c1_39808_21618# 0.15596f
C2398 a_66368_52081# sar10b_0._07_ 0.04879f
C2399 VSSR sar10b_0.SWN[9] 13.8206f
C2400 a_63273_56639# a_64233_56639# 0.03432f
C2401 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] 1.16488f
C2402 VSSR m3_23944_21578# 0.41298f
C2403 tdc_0.phase_detector_0.INP tdc_0.phase_detector_0.pd_out_0.B 0.06558f
C2404 VSSD a_60747_65563# 0.32267f
C2405 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y VDDR 0.31995f
C2406 VSSD a_62313_61671# 0.50859f
C2407 c1_45456_27218# VDDR 0.01151f
C2408 sar10b_0.net14 sar10b_0.net13 2.42075f
C2409 m3_45124_30538# th_dif_sw_0.VCN 0.17339f
C2410 sar10b_0.clk_div_0.COUNT\[2\] sar10b_0.net37 0.0382f
C2411 a_61929_51311# VSSD 0.26986f
C2412 sar10b_0.net21 a_68421_58960# 0.02929f
C2413 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 1.11457f
C2414 VSSD a_64993_66255# 0.86254f
C2415 VDDR a_38665_5788# 7.21057f
C2416 a_61400_50300# a_61677_50190# 0.09983f
C2417 a_68235_48621# a_68562_48647# 0.08997f
C2418 sar10b_0.cyclic_flag_0.FINAL a_67393_67963# 0.06815f
C2419 tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.pd_out_0.B 2.26706f
C2420 m3_18296_97932# VCM 0.13579f
C2421 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 3.47757f
C2422 a_61400_52964# sar10b_0.net16 0.13915f
C2423 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_39808_21618# 0.0106f
C2424 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] c1_22864_21618# 0.02548f
C2425 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] a_33863_5788# 2.38822f
C2426 a_68767_54656# VSSD 0.26653f
C2427 th_dif_sw_0.VCP VSSA 10.337f
C2428 c1_n1140_38418# c1_n1140_37298# 0.13255f
C2429 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.60057f
C2430 c1_24276_97972# th_dif_sw_0.VCP 0.13255f
C2431 VDDD a_64888_67630# 0.32273f
C2432 m3_22532_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.02509f
C2433 m3_43712_21578# VCM 0.15231f
C2434 m3_n1472_39498# m3_n1472_38378# 0.29566f
C2435 VSSR c1_n1140_85652# 0.04956f
C2436 sar10b_0.net46 sar10b_0.net14 0.15104f
C2437 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 0.19757f
C2438 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 0.02638f
C2439 sar10b_0.CF[4] sar10b_0.CF[7] 0.11432f
C2440 VSSD sar10b_0.net37 1.84864f
C2441 c1_272_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.01819f
C2442 a_65385_64631# a_65983_64966# 0.06623f
C2443 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 0.12357f
C2444 sar10b_0.CF[6] sar10b_0.SWN[0] 0.13195f
C2445 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y sar10b_0.CF[6] 0.12541f
C2446 sar10b_0.SWN[1] sar10b_0.SWN[0] 7.35755f
C2447 VDDD a_66785_50875# 0.62894f
C2448 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] sar10b_0.CF[9] 0.01482f
C2449 m3_n1472_97932# c1_n1140_97972# 1.74381f
C2450 VSSR m3_45124_51818# 0.63261f
C2451 a_69003_48621# sar10b_0.net36 0.25239f
C2452 VSSD a_62702_61352# 0.13843f
C2453 a_65301_57975# a_65577_57971# 0.1263f
C2454 sar10b_0.net16 a_65865_57675# 0.18368f
C2455 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 0.24788f
C2456 c1_n1140_28338# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C2457 sar10b_0.net9 a_63169_62635# 0.02029f
C2458 m3_8412_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C2459 sar10b_0.net22 a_68946_56639# 0.26111f
C2460 sar10b_0.net17 a_61419_48621# 0.24707f
C2461 sar10b_0.SWN[7] VSSD 1.18682f
C2462 a_64609_64923# sar10b_0.net11 0.01549f
C2463 sar10b_0.CF[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y 0.12541f
C2464 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 sar10b_0.SWN[7] 0.2638f
C2465 VSSR c1_7332_21618# 0.05923f
C2466 DATA[4] sar10b_0.net36 0.10523f
C2467 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.36778f
C2468 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] a_29061_5788# 2.08782f
C2469 sar10b_0.net14 a_62997_67299# 0.17301f
C2470 a_61833_57675# a_62222_57356# 0.05462f
C2471 a_61557_57735# a_62017_57307# 0.26257f
C2472 a_64188_51135# a_64199_50761# 0.54361f
C2473 a_66865_49412# sar10b_0.SWN[6] 0.05597f
C2474 VDDD a_67393_66631# 0.25319f
C2475 m3_n1472_80012# m3_n1472_78892# 0.29566f
C2476 a_63573_63303# sar10b_0.net16 0.29524f
C2477 VSSR m3_45124_92332# 0.63305f
C2478 VDDA sar10b_0.SWP[2] 0.2491f
C2479 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A 1.29717f
C2480 a_65961_68627# sar10b_0.net16 0.3256f
C2481 m3_45124_36138# VDDR 0.0103f
C2482 a_65394_52643# a_65928_53032# 0.35097f
C2483 a_61400_64952# a_62185_64695# 0.26257f
C2484 a_61609_64934# a_61677_64842# 0.35559f
C2485 VSSR c1_36984_97972# 0.05923f
C2486 a_62985_63003# VSSD 0.51405f
C2487 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_29592_21578# 0.03017f
C2488 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_12648_21578# 0.0162f
C2489 sar10b_0.SWN[6] VSSD 0.99419f
C2490 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A sar10b_0.CF[7] 0.06369f
C2491 c1_n1140_41778# m3_n1472_42858# 0.01078f
C2492 c1_45456_42898# m3_45124_42858# 1.74381f
C2493 c1_n1140_42898# m3_n1472_41738# 0.01078f
C2494 VDDD a_61609_50282# 0.21022f
C2495 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A 0.42509f
C2496 VSSD a_62185_64695# 0.15819f
C2497 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VSSR 4.36931f
C2498 sar10b_0.clk_div_0.COUNT\[2\] sar10b_0._03_ 0.22057f
C2499 m3_45124_76652# VDDR 0.01034f
C2500 m3_45124_73292# th_dif_sw_0.VCP 0.17339f
C2501 sar10b_0._07_ sar10b_0.clknet_1_0__leaf_CLK 0.14216f
C2502 c1_24276_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 0.01078f
C2503 sar10b_0.SWP[1] a_39543_110941# 0.71842f
C2504 m3_16884_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.19074f
C2505 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 1.79797f
C2506 VDDD a_62185_66027# 0.30535f
C2507 a_61153_58263# sar10b_0.net2 0.01484f
C2508 a_63369_59007# a_63621_58960# 0.27388f
C2509 a_61400_50300# a_60690_49683# 0.01135f
C2510 a_65021_50292# a_64818_49979# 0.06657f
C2511 a_67393_65299# a_67733_65447# 0.24088f
C2512 a_67209_65667# a_68169_65667# 0.03471f
C2513 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A 1.34718f
C2514 m3_45124_64332# c1_45456_65492# 0.01078f
C2515 m3_n1472_64332# c1_n1140_64372# 1.74381f
C2516 m3_45124_65452# c1_45456_64372# 0.01078f
C2517 VSSR c1_45456_62132# 0.12325f
C2518 sar10b_0.SWN[7] sar10b_0.CF[8] 0.12093f
C2519 a_68767_63980# VSSD 0.26642f
C2520 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 2.37545f
C2521 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VDDR 3.23491f
C2522 m3_38064_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.53746f
C2523 a_43467_5788# sar10b_0.SWN[0] 1.0688f
C2524 m3_14060_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.54821f
C2525 m3_39476_97932# m3_40888_97932# 0.23959f
C2526 c1_45456_82292# c1_45456_81172# 0.13255f
C2527 sar10b_0.net34 a_65957_50273# 0.02134f
C2528 m3_21120_21578# c1_20040_21618# 0.15596f
C2529 a_61249_53311# a_62025_53679# 0.3578f
C2530 m3_n1472_37258# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C2531 VDDR sar10b_0.SWN[8] 1.15764f
C2532 m3_23944_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.09358f
C2533 VSSD a_62185_60699# 0.15219f
C2534 sar10b_0._03_ VSSD 0.32905f
C2535 sar10b_0.net33 a_65682_51977# 0.03159f
C2536 a_60969_56639# a_61929_56639# 0.03432f
C2537 a_61153_56931# a_62181_56768# 0.07826f
C2538 m3_29592_97932# c1_28512_97972# 0.15596f
C2539 VSSD sar10b_0.CF[7] 0.7935f
C2540 VSSR m3_n1472_27178# 0.66371f
C2541 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 sar10b_0.CF[7] 0.40665f
C2542 sar10b_0._10_ sar10b_0._00_ 0.20507f
C2543 a_249_5788# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 0.02167f
C2544 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP sar10b_0.SWP[4] 0.26591f
C2545 c1_45456_42898# VDDR 0.01151f
C2546 m3_45124_46218# th_dif_sw_0.VCN 0.17339f
C2547 CLK a_51861_59345# 0.01174f
C2548 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 a_29939_5779# 0.51724f
C2549 sar10b_0.SWN[6] sar10b_0.CF[8] 0.12306f
C2550 sar10b_0.SWN[1] a_38665_5788# 0.96592f
C2551 a_n8277_54565# a_n9133_57045# 0.11069f
C2552 a_67393_62635# a_67733_62783# 0.24088f
C2553 a_67209_63003# a_68421_62956# 0.07766f
C2554 sar10b_0._05_ a_65821_53072# 0.1422f
C2555 a_61358_51694# CLK 0.01556f
C2556 a_61400_60956# a_62185_60699# 0.26257f
C2557 a_61609_60938# a_61677_60846# 0.35559f
C2558 m3_n1472_97932# VDDR 0.02674f
C2559 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 3.67813f
C2560 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C2561 a_66825_57675# a_67077_57628# 0.27388f
C2562 sar10b_0.net7 a_60690_54641# 0.01796f
C2563 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_12980_21618# 0.0106f
C2564 sar10b_0.net16 a_60969_56639# 0.1872f
C2565 sar10b_0.net1 a_61921_55975# 0.01927f
C2566 VDDR sar10b_0.SWN[9] 0.83216f
C2567 VSSR m3_n1472_67692# 0.66316f
C2568 sar10b_0.net10 a_63525_61624# 0.01302f
C2569 c1_n1140_46258# c1_n1140_45138# 0.13255f
C2570 VDDA a_n8277_66083# 1.54045f
C2571 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 0.02632f
C2572 a_60945_52617# VSSD 0.28664f
C2573 sar10b_0.net2 a_61461_56403# 0.22499f
C2574 m3_4176_21578# VCM 0.15231f
C2575 sar10b_0.net32 a_64485_56768# 0.02697f
C2576 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.41429f
C2577 sar10b_0.net39 th_dif_sw_0.CK 0.12018f
C2578 VDDD a_67077_57628# 0.31918f
C2579 c1_n1140_69972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C2580 m3_n1472_47338# m3_n1472_46218# 0.29566f
C2581 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.40207f
C2582 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.38262f
C2583 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C2584 sar10b_0.net33 sar10b_0._07_ 0.02973f
C2585 VDDD a_62187_48621# 0.26907f
C2586 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.95194f
C2587 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A sar10b_0.CF[1] 0.02149f
C2588 sar10b_0.net3 a_67209_68331# 0.17459f
C2589 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 2.67074f
C2590 sar10b_0.SWN[5] VSSD 1.36336f
C2591 VDDD a_60693_57975# 0.33881f
C2592 sar10b_0.SWN[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 0.44188f
C2593 sar10b_0._01_ sar10b_0.net16 0.3025f
C2594 sar10b_0.CF[1] VCM 3.52651f
C2595 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.72402f
C2596 sar10b_0.CF[3] sar10b_0.CF[9] 0.10503f
C2597 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.02632f
C2598 a_249_113874# sar10b_0.SWP[9] 0.11779f
C2599 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.1659f
C2600 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 0.02632f
C2601 th_dif_sw_0.VCP th_dif_sw_0.VCN 0.41613f
C2602 sar10b_0.CF[8] sar10b_0.CF[7] 60.8468f
C2603 c1_n1140_44018# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C2604 a_66921_61671# a_67445_61451# 0.04522f
C2605 sar10b_0.clk_div_0.COUNT\[1\] a_66961_50219# 0.11955f
C2606 a_66645_61731# a_67310_61352# 0.19065f
C2607 sar10b_0.net38 a_62181_56768# 0.02764f
C2608 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 17.3154f
C2609 sar10b_0.net40 sar10b_0.net8 0.08669f
C2610 VSSR c1_n1140_33938# 0.04956f
C2611 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] 2.33263f
C2612 a_61249_50647# a_62025_51015# 0.3578f
C2613 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[0] 0.05999f
C2614 a_65673_56639# a_66062_57022# 0.06034f
C2615 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[7] 0.01887f
C2616 VSSD a_61395_65944# 0.51728f
C2617 m3_45124_76652# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C2618 m3_n1472_87852# m3_n1472_86732# 0.29566f
C2619 VSSR m3_19708_97932# 0.40111f
C2620 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A 0.02842f
C2621 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP 3.06947f
C2622 m3_19708_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26144f
C2623 m3_45124_51818# VDDR 0.0103f
C2624 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 1.30896f
C2625 a_62185_50043# sar10b_0.net6 0.05284f
C2626 VDDD sar10b_0.clknet_1_1__leaf_CLK 2.49187f
C2627 a_63273_61671# a_63871_61316# 0.06623f
C2628 sar10b_0.net1 a_61833_57675# 0.01448f
C2629 VSSR m3_45124_21578# 0.68122f
C2630 VSSD sar10b_0.net25 0.62653f
C2631 VDDD a_63339_71265# 0.25557f
C2632 a_61131_70891# sar10b_0.net16 0.01551f
C2633 sar10b_0.net2 sar10b_0.net39 0.07102f
C2634 a_65525_68912# VSSD 0.08464f
C2635 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.22192f
C2636 a_66464_50363# VSSD 0.14475f
C2637 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.59327f
C2638 sar10b_0.net39 a_61609_66266# 0.01413f
C2639 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A 0.68875f
C2640 a_66933_64395# sar10b_0.cyclic_flag_0.FINAL 0.06705f
C2641 c1_n1140_49618# m3_n1472_50698# 0.01078f
C2642 c1_n1140_50738# m3_n1472_49578# 0.01078f
C2643 c1_45456_50738# m3_45124_50698# 1.74381f
C2644 c1_n1140_96852# c1_n1140_95732# 0.13255f
C2645 tdc_0.RDY sar10b_0.CF[1] 0.14529f
C2646 sar10b_0.net33 a_66103_50668# 0.02888f
C2647 a_61065_51015# a_61395_49960# 0.19391f
C2648 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[9] 0.17717f
C2649 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A a_6634_111636# 0.01076f
C2650 m3_45124_88972# th_dif_sw_0.VCP 0.17339f
C2651 m3_45124_92332# VDDR 0.01034f
C2652 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.12357f
C2653 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A VDDR 0.7488f
C2654 VDDD a_60747_56239# 0.29855f
C2655 sar10b_0.SWN[5] sar10b_0.CF[8] 0.12386f
C2656 m3_39476_97932# VCM 0.15231f
C2657 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A 0.42509f
C2658 a_66825_69663# sar10b_0.net44 0.02376f
C2659 sar10b_0.net22 sar10b_0.net36 0.16991f
C2660 a_68235_71265# sar10b_0.net15 0.01149f
C2661 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A 0.11547f
C2662 a_65394_52643# a_66378_52993# 0.08669f
C2663 sar10b_0.clknet_1_1__leaf_CLK sar10b_0._08_ 0.03013f
C2664 VDDD a_67297_55975# 0.26179f
C2665 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN 0.01239f
C2666 c1_17216_97972# VCM 0.01358f
C2667 m3_43712_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C2668 sar10b_0.SWN[8] DATA[0] 0.93863f
C2669 VDDA a_51345_58977# 0.6608f
C2670 sar10b_0.net3 a_66921_61671# 0.19361f
C2671 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN 0.12367f
C2672 m3_45124_72172# c1_45456_73332# 0.01078f
C2673 m3_45124_73292# c1_45456_72212# 0.01078f
C2674 m3_n1472_72172# c1_n1140_72212# 1.74381f
C2675 VSSR c1_45456_77812# 0.0935f
C2676 sar10b_0.net2 a_62037_61731# 0.17582f
C2677 sar10b_0.net13 a_60945_65937# 0.01361f
C2678 sar10b_0.net14 sar10b_0.net42 0.0641f
C2679 a_65577_51311# CLK 0.46794f
C2680 sar10b_0.net38 sar10b_0.net8 0.05984f
C2681 a_5929_5779# sar10b_0.SWN[8] 0.17051f
C2682 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VDDR 4.94582f
C2683 c1_21452_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.01302f
C2684 m3_19708_97932# m3_21120_97932# 0.23959f
C2685 c1_45456_90132# c1_45456_89012# 0.13255f
C2686 c1_7332_21618# m3_7000_21578# 1.74381f
C2687 m3_n1472_52938# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C2688 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A 0.11547f
C2689 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 sar10b_0.SWN[8] 0.37025f
C2690 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A 0.07418f
C2691 sar10b_0.SWP[0] sar10b_0.CF[0] 4.2293f
C2692 sar10b_0.net12 a_64533_65967# 0.05516f
C2693 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A 0.68875f
C2694 m3_9824_97932# c1_8744_97972# 0.15596f
C2695 VSSR m3_n1472_42858# 0.66365f
C2696 a_62277_53632# sar10b_0.net6 0.01042f
C2697 sar10b_0.clknet_0_CLK sar10b_0.clk_div_0.COUNT\[0\] 1.05131f
C2698 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A VDDR 0.74806f
C2699 sar10b_0.net16 sar10b_0.net35 0.05103f
C2700 a_61491_52222# a_61496_52091# 0.44532f
C2701 c1_3096_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26825f
C2702 sar10b_0.SWN[9] DATA[0] 0.06877f
C2703 c1_45456_62132# VDDR 0.01153f
C2704 m3_29592_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C2705 sar10b_0.net9 sar10b_0.net40 0.39399f
C2706 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.02638f
C2707 a_67209_55011# a_67393_54643# 0.43491f
C2708 VDDD a_64761_51028# 0.01371f
C2709 VDDD DATA[7] 0.4141f
C2710 a_63045_57628# a_63391_57320# 0.07649f
C2711 a_64199_50761# a_64356_51029# 0.21226f
C2712 a_64773_60292# sar10b_0.net12 0.02763f
C2713 VSSR m3_n1472_83372# 0.66316f
C2714 a_61929_57971# sar10b_0.net16 0.272f
C2715 a_67105_59971# a_67881_60339# 0.3578f
C2716 VDDD a_65821_53072# 0.0122f
C2717 c1_n1140_54098# c1_n1140_52978# 0.13255f
C2718 sar10b_0.net38 a_65673_56639# 0.02504f
C2719 sar10b_0.net40 a_61395_64612# 0.01738f
C2720 m3_n1472_27178# VDDR 0.02681f
C2721 VDDD a_68479_61316# 0.20677f
C2722 m3_n1472_35018# VCM 0.01415f
C2723 c1_n1140_85652# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C2724 m3_n1472_55178# m3_n1472_54058# 0.29566f
C2725 a_66933_63063# VSSD 0.13693f
C2726 a_60690_70625# sar10b_0.SWP[0] 0.1355f
C2727 VDDD a_67733_58787# 0.20874f
C2728 VDDD tdc_0.RDY 0.27371f
C2729 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_33828_21578# 0.0162f
C2730 sar10b_0.SWN[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.33822f
C2731 sar10b_0.net33 a_65394_52643# 0.02868f
C2732 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C2733 c1_35572_21618# VCM 0.01358f
C2734 VDDD a_61400_63620# 0.25201f
C2735 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP sar10b_0.CF[2] 0.10522f
C2736 m3_n1472_67692# VDDR 0.02674f
C2737 VDDD a_67890_69727# 0.2725f
C2738 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.26364f
C2739 sar10b_0.net10 a_64033_63591# 0.01551f
C2740 a_62409_59007# sar10b_0.net16 0.18184f
C2741 m3_n1472_75532# VCM 0.01412f
C2742 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38768f
C2743 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] m3_22532_21578# 0.24105f
C2744 sar10b_0.net30 a_62185_50043# 0.02044f
C2745 a_62527_58306# sar10b_0.net8 0.29066f
C2746 VDDD a_62181_51440# 0.26957f
C2747 VDDD a_61358_67678# 0.28627f
C2748 sar10b_0.net16 a_61395_49960# 0.17746f
C2749 a_67393_54643# sar10b_0.net35 0.01569f
C2750 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP 3.31931f
C2751 sar10b_0._02_ a_65682_49313# 0.10813f
C2752 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A 0.03718f
C2753 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_22076_8700# 0.01076f
C2754 c1_15804_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.01532f
C2755 sar10b_0.SWN[0] sar10b_0.CF[7] 0.14646f
C2756 a_62709_63063# sar10b_0.net2 0.2598f
C2757 m3_45124_23818# m3_45124_22698# 0.29566f
C2758 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 0.12068f
C2759 sar10b_0.clk_div_0.COUNT\[2\] sar10b_0._13_ 0.18202f
C2760 sar10b_0.net4 sar10b_0.net16 4.39867f
C2761 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A sar10b_0.CF[9] 0.03041f
C2762 VSSR c1_n1140_49618# 0.04956f
C2763 sar10b_0.net9 sar10b_0.net38 0.06034f
C2764 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A 0.28117f
C2765 VDDD a_68421_54964# 0.27498f
C2766 m3_45124_92332# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C2767 sar10b_0.net2 sar10b_0.net11 0.64152f
C2768 m3_n1472_95692# m3_n1472_94572# 0.29566f
C2769 m3_31004_21578# c1_31336_21618# 1.74381f
C2770 sar10b_0.net16 a_62126_56024# 0.20518f
C2771 m3_45124_29418# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C2772 a_62185_50043# VSSD 0.15433f
C2773 sar10b_0.net32 sar10b_0.net1 0.04449f
C2774 sar10b_0.net10 sar10b_0.net42 0.03955f
C2775 sar10b_0.net15 VSSD 0.95127f
C2776 VSSR a_29939_5779# 2.46707f
C2777 c1_36984_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26825f
C2778 sar10b_0.net13 sar10b_0.net42 0.05687f
C2779 m3_39476_97932# c1_39808_97972# 1.74381f
C2780 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 1.39288f
C2781 a_62133_59067# sar10b_0.net8 0.01826f
C2782 VSSR m3_5588_21578# 0.54637f
C2783 VDDD a_67231_56974# 0.24848f
C2784 c1_22864_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.01237f
C2785 VSSD EN 0.97579f
C2786 sar10b_0.net3 a_65861_49313# 0.04769f
C2787 a_64521_59303# VSSD 0.50558f
C2788 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 sar10b_0.CF[0] 0.40695f
C2789 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP a_25137_5779# 0.01111f
C2790 sar10b_0._13_ VSSD 0.67456f
C2791 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A sar10b_0.SWN[1] 0.02058f
C2792 sar10b_0.clk_div_0.COUNT\[0\] a_68178_51635# 0.10732f
C2793 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 0.51491f
C2794 m3_n60_97932# VCM 0.15231f
C2795 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A 0.68875f
C2796 a_54660_59599# tdc_0.OUTN 0.01287f
C2797 VDDD a_62497_61303# 0.22368f
C2798 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_21452_21618# 0.01302f
C2799 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN sar10b_0.SWP[8] 0.1944f
C2800 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C2801 m3_45124_64332# m3_45124_63212# 0.29566f
C2802 a_n8277_54565# th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 1.59491f
C2803 sar10b_0.net41 a_64533_65967# 0.0119f
C2804 sar10b_0.net4 a_60969_67295# 0.22614f
C2805 a_60693_67299# a_61153_67587# 0.26257f
C2806 m3_45124_21578# VDDR 0.0103f
C2807 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A 0.42509f
C2808 a_60747_61941# a_60945_61941# 0.06623f
C2809 a_65928_53032# VSSD 0.12206f
C2810 VDDD a_69003_48621# 0.26823f
C2811 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP 3.9628f
C2812 m3_25356_21578# VCM 0.13579f
C2813 m3_4176_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C2814 VCM sar10b_0.CF[2] 3.51908f
C2815 sar10b_0._10_ sar10b_0._09_ 0.96152f
C2816 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.88327f
C2817 sar10b_0.CF[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP 0.18426f
C2818 m3_n1472_80012# c1_n1140_80052# 1.74381f
C2819 m3_45124_81132# c1_45456_80052# 0.01078f
C2820 m3_45124_80012# c1_45456_81172# 0.01078f
C2821 VSSR c1_45456_93492# 0.0935f
C2822 sar10b_0.SWP[4] sar10b_0.CF[9] 0.18445f
C2823 a_61833_57675# a_62527_56974# 0.0165f
C2824 sar10b_0.clk_div_0.COUNT\[1\] sar10b_0.net35 0.14462f
C2825 sar10b_0.SWP[9] CKO 0.06745f
C2826 th_dif_sw_0.CK th_dif_sw_0.th_sw_1.CKB 0.02097f
C2827 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 0.19711f
C2828 m3_n60_97932# m3_1352_97932# 0.23959f
C2829 VDDD a_64814_65014# 0.26071f
C2830 VDDD DATA[4] 0.33066f
C2831 c1_45456_26098# m3_45124_27178# 0.01078f
C2832 c1_45456_27218# m3_45124_26058# 0.01078f
C2833 c1_n1140_26098# m3_n1472_26058# 1.74381f
C2834 sar10b_0.net40 a_62222_57356# 0.03105f
C2835 sar10b_0.net20 sar10b_0._13_ 0.02199f
C2836 a_64773_60292# sar10b_0.net41 0.07202f
C2837 sar10b_0.net14 a_65673_56639# 0.22299f
C2838 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 0.02632f
C2839 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP sar10b_0.SWP[0] 0.35086f
C2840 a_62277_53632# VSSD 0.27176f
C2841 VDDD sar10b_0.SWP[3] 0.36357f
C2842 sar10b_0.net8 a_63457_56931# 0.01765f
C2843 sar10b_0.net16 a_61557_57735# 0.23044f
C2844 c1_45456_77812# VDDR 0.01153f
C2845 sar10b_0.net34 sar10b_0._10_ 0.02593f
C2846 sar10b_0.net27 DATA[9] 0.04878f
C2847 a_68133_61624# a_68479_61316# 0.07649f
C2848 m3_25356_21578# m3_26768_21578# 0.23959f
C2849 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y 0.32324f
C2850 sar10b_0.net38 a_64485_56768# 0.02972f
C2851 VSSR c1_45456_26098# 0.09348f
C2852 a_62277_50968# sar10b_0.net30 0.02773f
C2853 sar10b_0._01_ a_65682_51977# 0.04049f
C2854 a_62185_63363# sar10b_0.net16 0.29833f
C2855 VDDD a_61705_51992# 0.20713f
C2856 m3_n1472_67692# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C2857 a_65682_49313# a_66865_49412# 0.0649f
C2858 a_65861_49313# a_66666_49313# 0.29221f
C2859 a_66109_49318# a_66216_49358# 0.14439f
C2860 sar10b_0.clknet_1_0__leaf_CLK sar10b_0._02_ 0.19317f
C2861 a_64725_68631# sar10b_0.net16 0.22244f
C2862 VSSR m3_40888_97932# 0.54637f
C2863 c1_n1140_65492# c1_n1140_64372# 0.13255f
C2864 tdc_0.RDY sar10b_0.CF[2] 0.13655f
C2865 VDDD a_63967_58652# 0.20924f
C2866 m3_40888_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.53746f
C2867 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP a_19457_110450# 0.11862f
C2868 m3_n1472_42858# VDDR 0.02681f
C2869 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP 0.10502f
C2870 m3_n1472_50698# VCM 0.01415f
C2871 a_66368_52081# VSSD 0.14369f
C2872 a_62133_59067# sar10b_0.net9 0.03041f
C2873 a_61493_58256# VSSD 0.09866f
C2874 a_67598_58688# a_67733_58787# 0.35559f
C2875 VDDD a_68421_64288# 0.27523f
C2876 sar10b_0.net1 a_65589_57735# 0.17188f
C2877 VSSR c1_18628_97972# 0.05435f
C2878 a_55282_59893# tdc_0.RDY 0.06067f
C2879 sar10b_0.net16 sar10b_0.net44 0.05713f
C2880 VDDD a_65589_69723# 0.30005f
C2881 a_62277_50968# VSSD 0.26908f
C2882 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45324f
C2883 a_60789_53739# sar10b_0.net16 0.22304f
C2884 a_65682_49313# VSSD 1.14236f
C2885 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_11236_21578# 0.03017f
C2886 m3_19708_21578# th_dif_sw_0.VCN 0.01078f
C2887 c1_8744_21618# VCM 0.01358f
C2888 sar10b_0.net28 sar10b_0.net6 0.02005f
C2889 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A 0.04073f
C2890 sar10b_0.net34 sar10b_0.net39 0.03645f
C2891 a_61086_63306# a_61400_63620# 0.07826f
C2892 a_61395_63280# a_61609_63602# 0.04522f
C2893 sar10b_0.clknet_0_CLK sar10b_0.SWN[6] 0.08077f
C2894 m3_n1472_83372# VDDR 0.02674f
C2895 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 0.73278f
C2896 a_5051_5788# VSSR 0.06023f
C2897 c1_18628_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 0.02099f
C2898 m3_n1472_91212# VCM 0.01412f
C2899 a_61395_65944# a_61677_66174# 0.05462f
C2900 sar10b_0.net9 a_60747_60609# 0.30099f
C2901 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.94823f
C2902 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.44217f
C2903 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.41774f
C2904 sar10b_0.net46 CKO 0.04461f
C2905 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_7670_111642# 0.01076f
C2906 sar10b_0._01_ sar10b_0._07_ 0.09277f
C2907 c1_45456_30578# c1_45456_29458# 0.13255f
C2908 a_62409_59007# a_62798_58688# 0.05462f
C2909 a_62133_59067# a_62593_58639# 0.26257f
C2910 c1_38396_97972# VCM 0.01358f
C2911 m3_45124_31658# m3_45124_30538# 0.29566f
C2912 sar10b_0.SWN[7] sar10b_0.SWN[8] 19.5411f
C2913 VSSR c1_n1140_68852# 0.04956f
C2914 VDDD sar10b_0.net27 0.35269f
C2915 sar10b_0.CF[5] sar10b_0.SWN[2] 0.12161f
C2916 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C2917 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP 5.56715f
C2918 VDDA a_53564_59480# 0.51472f
C2919 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 2.75475f
C2920 m3_19708_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26144f
C2921 c1_42632_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C2922 a_68421_58960# sar10b_0.net3 0.1775f
C2923 a_61153_51603# a_61929_51311# 0.3578f
C2924 c1_17216_21618# m3_18296_21578# 0.15596f
C2925 VDDD a_61395_52624# 0.77345f
C2926 m3_45124_45098# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C2927 sar10b_0.net16 a_63273_61671# 0.26588f
C2928 a_60693_56643# a_60969_56639# 0.1263f
C2929 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A sar10b_0.CF[0] 0.06396f
C2930 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 2.75442f
C2931 a_68133_60292# VSSD 0.27172f
C2932 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] sar10b_0.SWP[5] 0.07355f
C2933 m3_19708_97932# c1_20040_97972# 1.74381f
C2934 sar10b_0.net16 a_63273_67295# 0.1707f
C2935 a_64533_65967# a_64993_66255# 0.26257f
C2936 VSSR m3_45124_35018# 0.63261f
C2937 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN sar10b_0.SWN[6] 0.20927f
C2938 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP 0.02666f
C2939 sar10b_0.clknet_0_CLK sar10b_0._03_ 0.33316f
C2940 sar10b_0.net43 sar10b_0.net12 0.10909f
C2941 a_68178_51635# sar10b_0.net37 0.01151f
C2942 sar10b_0.net33 sar10b_0._02_ 0.01596f
C2943 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A sar10b_0.CF[8] 0.06369f
C2944 VDDD a_66153_48647# 1.47329f
C2945 VSSR c1_36984_21618# 0.05923f
C2946 sar10b_0.net21 DATA[3] 0.0128f
C2947 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A sar10b_0.CF[8] 0.03041f
C2948 a_68169_55011# a_68421_54964# 0.27388f
C2949 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR 0.41774f
C2950 a_65865_57675# a_66389_57455# 0.04522f
C2951 a_65589_57735# a_66254_57356# 0.19065f
C2952 m3_45124_72172# m3_45124_71052# 0.29566f
C2953 VSSR m3_45124_75532# 0.63305f
C2954 VDDD a_61773_52237# 0.26254f
C2955 sar10b_0.net33 a_66079_59638# 0.02667f
C2956 sar10b_0.net7 a_61086_52650# 0.01476f
C2957 sar10b_0.CF[0] th_dif_sw_0.CK 0.08524f
C2958 a_63374_62684# sar10b_0.net16 0.21402f
C2959 a_61921_55975# a_62949_56296# 0.07826f
C2960 VSSD a_63273_56639# 0.52997f
C2961 sar10b_0.net27 a_68767_67976# 0.27724f
C2962 a_64199_50761# sar10b_0.net16 0.03369f
C2963 m3_n1472_87852# c1_n1140_87892# 1.74381f
C2964 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP sar10b_0.CF[4] 0.10502f
C2965 m3_45124_87852# c1_45456_89012# 0.01078f
C2966 m3_45124_88972# c1_45456_87892# 0.01078f
C2967 VDDD a_60747_65937# 0.21802f
C2968 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP 2.62898f
C2969 sar10b_0.CF[3] sar10b_0.SWP[2] 0.12013f
C2970 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A 1.11457f
C2971 sar10b_0._04_ a_66109_51982# 0.14027f
C2972 a_65861_51977# a_66216_52022# 0.18752f
C2973 c1_n1140_33938# m3_n1472_33898# 1.74381f
C2974 c1_45456_33938# m3_45124_35018# 0.01078f
C2975 c1_45456_35058# m3_45124_33898# 0.01078f
C2976 a_n4470_65264# a_n8277_66083# 0.01412f
C2977 sar10b_0._11_ sar10b_0.net16 0.21012f
C2978 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN sar10b_0.CF[7] 0.06929f
C2979 sar10b_0.net1 a_61153_56931# 0.05242f
C2980 sar10b_0.net10 sar10b_0.net9 0.05934f
C2981 a_65577_51311# a_65586_50645# 0.01255f
C2982 VSSR VCM 0.18541p
C2983 VDDD a_65185_68919# 0.2203f
C2984 sar10b_0.clknet_1_0__leaf_CLK VSSD 1.3617f
C2985 a_67393_66631# a_67598_66680# 0.09983f
C2986 sar10b_0.net33 a_65857_56931# 0.02463f
C2987 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP 4.32584f
C2988 a_63849_63299# a_65061_63428# 0.07766f
C2989 a_66633_56639# a_67231_56974# 0.06623f
C2990 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.01212f
C2991 a_62281_52347# sar10b_0.net6 0.18495f
C2992 VDDD a_65957_50273# 0.84404f
C2993 tdc_0.phase_detector_0.INP a_53564_59480# 0.01732f
C2994 a_66378_52993# VSSD 0.20797f
C2995 sar10b_0.net40 sar10b_0.net1 0.09483f
C2996 c1_45456_93492# VDDR 0.01153f
C2997 sar10b_0._00_ a_65021_50292# 0.13368f
C2998 sar10b_0._07_ sar10b_0.net35 0.06831f
C2999 m3_5588_21578# m3_7000_21578# 0.23959f
C3000 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A 0.03718f
C3001 VSSR c1_45456_41778# 0.09348f
C3002 sar10b_0.net32 a_64338_52411# 0.01926f
C3003 sar10b_0.SWN[0] EN 0.17151f
C3004 th_dif_sw_0.VCP CLK 3.60859f
C3005 sar10b_0.net28 sar10b_0.net30 0.16046f
C3006 a_68169_59007# VSSD 0.29116f
C3007 m3_n1472_83372# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C3008 a_66961_50219# a_66762_50329# 0.29821f
C3009 VDDD a_64910_59686# 0.26589f
C3010 sar10b_0.net40 a_61400_66284# 0.02782f
C3011 tdc_0.phase_detector_0.pd_out_0.A a_53564_59480# 0.48002f
C3012 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 3.70212f
C3013 VSSR m3_1352_97932# 0.54637f
C3014 c1_n1140_73332# c1_n1140_72212# 0.13255f
C3015 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 2.76569f
C3016 m3_42300_21578# c1_41220_21618# 0.15596f
C3017 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A 0.45324f
C3018 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A a_21040_111636# 0.01076f
C3019 VDDA tdc_0.phase_detector_0.INP 0.58279f
C3020 m3_1352_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.53746f
C3021 a_61677_63510# VSSD 0.1344f
C3022 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y sar10b_0.CF[8] 0.12541f
C3023 tdc_0.RDY tdc_0.OUTN 1.78771f
C3024 a_63457_56931# a_64485_56768# 0.07826f
C3025 a_64033_63591# sar10b_0.net42 0.01613f
C3026 VDDD a_68562_71291# 0.22501f
C3027 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[9] 0.05939f
C3028 VDDD sar10b_0.net22 1.09741f
C3029 VSSA tdc_0.phase_detector_0.INN 1.76841f
C3030 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN sar10b_0.CF[9] 0.12367f
C3031 VSSR m3_26768_21578# 0.44047f
C3032 VSSD a_66933_65727# 0.13622f
C3033 a_51345_58977# tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A 0.14814f
C3034 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y 0.32264f
C3035 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y 0.31983f
C3036 c1_45456_26098# VDDR 0.01151f
C3037 sar10b_0.CF[5] th_dif_sw_0.VCP 0.28799f
C3038 m3_45124_29418# th_dif_sw_0.VCN 0.17339f
C3039 sar10b_0.net28 VSSD 0.91414f
C3040 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSSR 41.7127f
C3041 VDDA tdc_0.phase_detector_0.pd_out_0.A 1.7275f
C3042 a_68946_53975# VSSD 0.33131f
C3043 VSSD a_66021_66092# 0.27245f
C3044 m3_n1472_57418# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24058f
C3045 sar10b_0.clknet_0_CLK a_66464_50363# 0.03367f
C3046 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_46086_8700# 0.01076f
C3047 a_66049_69295# sar10b_0.net45 0.01542f
C3048 a_61400_50300# a_62185_50043# 0.26257f
C3049 a_61609_50282# a_61677_50190# 0.35559f
C3050 a_68235_48621# sar10b_0.SWN[7] 0.15191f
C3051 a_68562_48647# a_69003_48621# 0.02339f
C3052 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.36422f
C3053 m3_21120_97932# VCM 0.6299f
C3054 a_61609_52946# sar10b_0.net16 0.18087f
C3055 c1_45456_57458# m3_45124_57418# 1.74381f
C3056 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_42632_21618# 0.0106f
C3057 a_68562_49747# sar10b_0.net37 0.26095f
C3058 c1_45456_38418# c1_45456_37298# 0.13255f
C3059 sar10b_0.SWP[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 0.29562f
C3060 c1_27100_97972# th_dif_sw_0.VCP 0.13255f
C3061 a_66645_60399# sar10b_0.cyclic_flag_0.FINAL 0.06403f
C3062 th_dif_sw_0.CK VSSA 6.89816f
C3063 VDDA th_dif_sw_0.CKB 5.37713f
C3064 m3_25356_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C3065 sar10b_0.net41 sar10b_0.net43 0.12975f
C3066 c1_n1140_97972# VCM 0.01358f
C3067 sar10b_0.net32 sar10b_0.net3 0.16133f
C3068 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 0.01239f
C3069 m3_45124_39498# m3_45124_38378# 0.29566f
C3070 sar10b_0.net38 sar10b_0.net1 0.14816f
C3071 VSSR c1_n1140_84532# 0.04956f
C3072 sar10b_0.net33 VSSD 1.4639f
C3073 a_60690_70625# sar10b_0.net2 0.23844f
C3074 CLK sar10b_0.net1 0.14098f
C3075 c1_3096_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C3076 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 2.80665f
C3077 a_64725_68631# a_65390_69010# 0.19065f
C3078 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 0.1659f
C3079 tdc_0.RDY a_60747_52617# 0.01224f
C3080 a_5051_5788# VDDR 1.62771f
C3081 sar10b_0.net40 a_66254_57356# 0.0337f
C3082 a_62185_66027# sar10b_0.net12 0.17711f
C3083 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.10847f
C3084 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38377f
C3085 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VSSR 2.16373f
C3086 sar10b_0.net20 a_68946_53975# 0.0227f
C3087 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 0.13856p
C3088 th_dif_sw_0.th_sw_1.CK th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 0.22595f
C3089 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.43221f
C3090 VDDD a_67209_63003# 0.89591f
C3091 DATA[6] sar10b_0.net22 0.02281f
C3092 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A 0.68875f
C3093 m3_n60_97932# c1_272_97972# 1.74381f
C3094 m3_n1472_57418# m3_n1472_56298# 0.29566f
C3095 VSSR m3_45124_50698# 0.63261f
C3096 c1_27100_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.02009f
C3097 a_67209_68331# a_68169_68331# 0.03471f
C3098 a_67393_67963# a_67733_68111# 0.24088f
C3099 c1_n1140_27218# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C3100 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] m3_21120_97932# 0.59034f
C3101 m3_11236_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C3102 sar10b_0.net17 a_62187_48621# 0.05539f
C3103 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP 6.77343f
C3104 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C3105 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A 0.10815f
C3106 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A VSSR 0.43773f
C3107 VSSR c1_10156_21618# 0.06746f
C3108 a_5051_113018# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 0.18139f
C3109 sar10b_0.net46 a_67055_68689# 0.01267f
C3110 a_64188_51135# a_64356_51029# 0.27693f
C3111 sar10b_0.net41 a_64888_67630# 0.02621f
C3112 VDDD a_67733_66779# 0.21283f
C3113 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y VSSR 0.32296f
C3114 a_66577_52883# sar10b_0.clk_div_0.COUNT\[3\] 0.12998f
C3115 m3_21120_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 0.59034f
C3116 m3_45124_80012# m3_45124_78892# 0.29566f
C3117 VSSR m3_45124_91212# 0.63305f
C3118 sar10b_0.net4 a_63457_67583# 0.01542f
C3119 VDDD a_65966_58354# 0.26916f
C3120 sar10b_0.cyclic_flag_0.FINAL sar10b_0.net16 0.13672f
C3121 m3_45124_35018# VDDR 0.0103f
C3122 tdc_0.phase_detector_0.pd_out_0.A tdc_0.phase_detector_0.INP 0.03298f
C3123 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN sar10b_0.CF[8] 0.05164f
C3124 a_68767_58652# sar10b_0.net19 0.27351f
C3125 VSSR c1_39808_97972# 0.05923f
C3126 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.11547f
C3127 sar10b_0.net4 a_60693_56643# 0.01673f
C3128 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_32416_21578# 0.03017f
C3129 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_15472_21578# 0.0162f
C3130 a_61491_52222# a_61929_51311# 0.01304f
C3131 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR 0.38377f
C3132 c1_45456_42898# m3_45124_41738# 0.01078f
C3133 c1_n1140_41778# m3_n1472_41738# 1.74381f
C3134 c1_45456_41778# m3_45124_42858# 0.01078f
C3135 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 1.70485f
C3136 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 0.20503f
C3137 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.4249f
C3138 a_67209_59007# sar10b_0.cyclic_flag_0.FINAL 0.24084f
C3139 m3_45124_75532# VDDR 0.01034f
C3140 m3_45124_72172# th_dif_sw_0.VCP 0.17339f
C3141 sar10b_0.CF[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP 0.10502f
C3142 m3_19708_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.18393f
C3143 sar10b_0.net7 sar10b_0.CF[0] 0.1925f
C3144 sar10b_0.clk_div_0.COUNT\[0\] a_66785_50875# 0.13658f
C3145 a_63285_60399# sar10b_0.net11 0.01461f
C3146 a_62281_52347# VSSD 0.13819f
C3147 sar10b_0.net9 a_61395_61948# 0.07277f
C3148 VSSR sar10b_0.SWP[3] 5.13254f
C3149 a_63621_58960# a_63967_58652# 0.07649f
C3150 VDDD a_64245_59307# 0.28924f
C3151 a_65778_49979# a_66762_50329# 0.08669f
C3152 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 2.45542f
C3153 sar10b_0._05_ sar10b_0._10_ 0.0829f
C3154 VDDD a_68331_52243# 0.24598f
C3155 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VSSR 2.9143f
C3156 m3_45124_64332# c1_45456_64372# 1.74381f
C3157 m3_n1472_64332# c1_n1140_63252# 0.01078f
C3158 m3_n1472_63212# c1_n1140_64372# 0.01078f
C3159 VSSR c1_45456_57458# 0.12458f
C3160 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VDDR 0.95194f
C3161 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A sar10b_0.CF[9] 0.03041f
C3162 sar10b_0.net19 sar10b_0.net18 0.44772f
C3163 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] th_dif_sw_0.VCN 2.24218f
C3164 a_66254_69344# VSSD 0.13583f
C3165 VDDD a_60690_54641# 0.44488f
C3166 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 sar10b_0.CF[3] 0.26289f
C3167 m3_40888_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.53746f
C3168 m3_16884_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.19074f
C3169 m3_40888_97932# m3_42300_97932# 0.23959f
C3170 a_68169_64335# a_68421_64288# 0.27388f
C3171 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C3172 c1_n1140_81172# c1_n1140_80052# 0.13255f
C3173 m3_22532_21578# c1_21452_21618# 0.15596f
C3174 sar10b_0.net34 a_66312_50368# 0.01418f
C3175 VDDR VCM 0.27737p
C3176 a_61589_53459# a_62025_53679# 0.16939f
C3177 m3_n1472_36138# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C3178 VDDD a_66080_53027# 0.10902f
C3179 a_51345_58977# sar10b_0.CF[3] 0.02111f
C3180 m3_26768_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.33071f
C3181 a_62133_59067# sar10b_0.net1 0.1682f
C3182 a_60789_51075# CLK 0.01125f
C3183 sar10b_0.cyclic_flag_0.FINAL a_67393_54643# 0.07077f
C3184 a_61493_56924# a_61929_56639# 0.16939f
C3185 a_60969_56639# a_61358_57022# 0.06034f
C3186 a_65865_69663# a_65589_69723# 0.1263f
C3187 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C3188 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A 0.02149f
C3189 m3_31004_97932# c1_29924_97972# 0.15596f
C3190 VSSR m3_n1472_26058# 0.66371f
C3191 sar10b_0.net14 sar10b_0.net1 0.1157f
C3192 a_61395_49960# a_60945_49953# 0.03529f
C3193 a_60747_49953# a_61086_49986# 0.07649f
C3194 a_67209_66999# a_68421_66952# 0.07766f
C3195 c1_45456_41778# VDDR 0.01151f
C3196 m3_45124_45098# th_dif_sw_0.VCN 0.17339f
C3197 sar10b_0.net43 a_64993_66255# 0.01008f
C3198 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A sar10b_0.CF[3] 0.03041f
C3199 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A 0.10815f
C3200 sar10b_0.net3 a_67439_50041# 0.09794f
C3201 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 3.50692f
C3202 sar10b_0.net4 a_61400_62288# 0.01899f
C3203 m3_9824_97932# th_dif_sw_0.VCP 0.01078f
C3204 VDDD a_62025_53679# 0.36509f
C3205 a_67209_68331# sar10b_0.net45 0.01455f
C3206 a_67077_57628# a_67423_57320# 0.07649f
C3207 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_15804_21618# 0.0106f
C3208 sar10b_0.net16 a_61493_56924# 0.15138f
C3209 VSSR m3_n1472_66572# 0.66316f
C3210 c1_45456_46258# c1_45456_45138# 0.13255f
C3211 th_dif_sw_0.VCP a_51861_60437# 0.06955f
C3212 VCM sar10b_0.SWP[7] 0.13075f
C3213 a_61400_52964# VSSD 0.84845f
C3214 sar10b_0.net2 a_61921_55975# 0.04149f
C3215 sar10b_0.net32 a_64831_56974# 0.01202f
C3216 m3_7000_21578# VCM 0.15231f
C3217 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y VDDR 0.3196f
C3218 c1_n1140_68852# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C3219 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[7] 0.01887f
C3220 m3_45124_47338# m3_45124_46218# 0.29566f
C3221 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VDDR 9.88107f
C3222 sar10b_0.clknet_1_1__leaf_CLK a_65573_52937# 0.05024f
C3223 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN 5.64431f
C3224 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26364f
C3225 a_5051_5788# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 0.18139f
C3226 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.59835f
C3227 a_66762_50329# sar10b_0.net35 0.01114f
C3228 VDDD a_66109_51982# 0.01215f
C3229 VDDD a_61153_58263# 0.2711f
C3230 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A 0.05472f
C3231 a_61496_52091# a_61705_51992# 0.24088f
C3232 VDDD a_62025_51015# 0.35139f
C3233 a_60693_57975# a_60969_57971# 0.1263f
C3234 VDDD a_65068_49569# 0.34685f
C3235 c1_n1140_42898# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C3236 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y sar10b_0.CF[0] 0.12541f
C3237 a_16238_111636# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A 0.01076f
C3238 sar10b_0.CF[4] sar10b_0.CF[9] 0.1099f
C3239 sar10b_0.SWN[8] EN 0.86532f
C3240 a_61065_53679# sar10b_0.net5 0.01672f
C3241 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C3242 VSSD a_65865_57675# 0.46984f
C3243 sar10b_0.net38 a_62527_56974# 0.28463f
C3244 VSSR c1_n1140_32818# 0.04956f
C3245 a_61589_50795# a_62025_51015# 0.16939f
C3246 a_64780_52239# sar10b_0._01_ 0.03706f
C3247 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VDDR 2.47806f
C3248 a_64454_51311# sar10b_0.net16 0.21416f
C3249 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.02842f
C3250 VSSD DATA[8] 0.6719f
C3251 sar10b_0._16_ sar10b_0._14_ 0.04736f
C3252 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.95198f
C3253 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.11339f
C3254 m3_45124_75532# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C3255 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VDDR 2.57696f
C3256 a_61153_67587# sar10b_0.net40 0.01105f
C3257 m3_45124_87852# m3_45124_86732# 0.29566f
C3258 VSSR m3_22532_97932# 0.34286f
C3259 m3_22532_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.21489f
C3260 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] a_9853_5788# 0.88621f
C3261 a_64425_64631# sar10b_0.net42 0.02343f
C3262 m3_45124_50698# VDDR 0.0103f
C3263 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A 0.11547f
C3264 a_63573_63303# VSSD 0.16268f
C3265 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A 0.01751f
C3266 sar10b_0.net39 a_61677_62178# 0.01946f
C3267 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_22076_111642# 0.01076f
C3268 VDDD a_68276_50645# 0.27392f
C3269 VSSR c1_272_97972# 0.05576f
C3270 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[9] 0.05939f
C3271 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.02632f
C3272 a_65961_68627# VSSD 0.26016f
C3273 a_64705_59595# sar10b_0.net16 0.11098f
C3274 sar10b_0._09_ a_65021_50292# 0.17409f
C3275 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.11339f
C3276 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[5] 0.01887f
C3277 sar10b_0.SWN[9] EN 8.61858f
C3278 a_67393_62635# sar10b_0.net3 0.13196f
C3279 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 3.24826f
C3280 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A VDDR 0.38472f
C3281 a_66961_50219# VSSD 0.33699f
C3282 sar10b_0.net3 sar10b_0.net40 0.13267f
C3283 sar10b_0.net2 a_61833_57675# 0.01757f
C3284 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP sar10b_0.SWP[1] 0.32962f
C3285 a_67393_63967# sar10b_0.cyclic_flag_0.FINAL 0.02261f
C3286 c1_45456_49618# m3_45124_50698# 0.01078f
C3287 c1_45456_50738# m3_45124_49578# 0.01078f
C3288 c1_n1140_49618# m3_n1472_49578# 1.74381f
C3289 c1_45456_96852# c1_45456_95732# 0.13255f
C3290 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26364f
C3291 a_63273_67295# a_63457_67583# 0.44457f
C3292 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 0.21389f
C3293 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y VDDR 0.31995f
C3294 sar10b_0.clknet_0_CLK a_65682_49313# 0.03011f
C3295 sar10b_0.net10 sar10b_0.net1 0.01389f
C3296 m3_45124_91212# VDDR 0.01034f
C3297 m3_45124_87852# th_dif_sw_0.VCP 0.17339f
C3298 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VCM 6.3144f
C3299 VDDD a_67881_60339# 0.3686f
C3300 VDDD a_61461_56403# 0.30866f
C3301 m3_42300_97932# VCM 0.15231f
C3302 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A 0.39707f
C3303 sar10b_0.net13 sar10b_0.net1 0.17065f
C3304 sar10b_0.net3 a_68421_66952# 0.17732f
C3305 VDDD a_67637_56123# 0.21257f
C3306 a_65573_52937# a_65821_53072# 0.05308f
C3307 m3_n1472_57418# th_dif_sw_0.VCN 0.12457f
C3308 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A sar10b_0.SWN[1] 0.01417f
C3309 sar10b_0.net28 a_61400_50300# 0.02214f
C3310 c1_20040_97972# VCM 0.01358f
C3311 sar10b_0._13_ a_68178_51635# 0.01037f
C3312 a_63745_59971# sar10b_0.net16 0.12981f
C3313 VDDA tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A 0.44525f
C3314 sar10b_0.net16 a_65397_56643# 0.22618f
C3315 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A 0.41861f
C3316 m3_45124_72172# c1_45456_72212# 1.74381f
C3317 m3_n1472_71052# c1_n1140_72212# 0.01078f
C3318 m3_n1472_72172# c1_n1140_71092# 0.01078f
C3319 VSSR c1_45456_76692# 0.0935f
C3320 sar10b_0.CF[6] VCM 3.50537f
C3321 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C3322 m3_1352_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.53746f
C3323 sar10b_0.SWN[1] VCM 0.13076f
C3324 a_66933_68391# VSSD 0.13445f
C3325 c1_24276_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C3326 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN 0.01131f
C3327 m3_21120_97932# m3_22532_97932# 0.23959f
C3328 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y 0.07418f
C3329 VDDD sar10b_0._10_ 0.80548f
C3330 c1_n1140_89012# c1_n1140_87892# 0.13255f
C3331 c1_8744_21618# m3_8412_21578# 1.74381f
C3332 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VCM 0.1236f
C3333 m3_n1472_51818# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C3334 a_63339_71265# sar10b_0.net41 0.25532f
C3335 VDDD a_62997_56643# 0.27772f
C3336 sar10b_0.net3 a_64339_51661# 0.14299f
C3337 a_64705_59595# a_65733_59432# 0.07826f
C3338 sar10b_0.net4 a_60690_53975# 0.37735f
C3339 VDDD sar10b_0.net24 0.48926f
C3340 m3_11236_97932# c1_10156_97972# 0.15596f
C3341 VDDR sar10b_0.SWP[3] 2.86289f
C3342 VSSR m3_n1472_41738# 0.66371f
C3343 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR 2.61522f
C3344 tdc_0.OUTP a_60690_70625# 0.29632f
C3345 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN 6.45047f
C3346 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VDDR 2.62902f
C3347 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.39589f
C3348 c1_5920_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26825f
C3349 a_61496_52091# a_61773_52237# 0.09983f
C3350 a_65586_50645# a_66255_50749# 0.27709f
C3351 c1_45456_57458# VDDR 0.01151f
C3352 m3_32416_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C3353 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A sar10b_0.CF[3] 0.26294f
C3354 a_63169_62635# a_64197_62956# 0.07826f
C3355 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 0.02632f
C3356 sar10b_0.net34 a_66577_52883# 0.02519f
C3357 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] th_dif_sw_0.VCN 0.27764p
C3358 sar10b_0.net38 sar10b_0.net3 0.15334f
C3359 a_64149_64635# sar10b_0.net16 0.24657f
C3360 a_67209_55011# a_67733_54791# 0.04522f
C3361 a_66933_55071# a_67598_54692# 0.19065f
C3362 sar10b_0._10_ sar10b_0._08_ 0.06035f
C3363 sar10b_0.SWN[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A 0.02025f
C3364 VINP a_n8277_66083# 0.64084f
C3365 a_55121_59650# VSSA 0.22099f
C3366 VSSD sar10b_0.CF[9] 0.65311f
C3367 sar10b_0.net3 CLK 0.08752f
C3368 VSSR m3_n1472_82252# 0.66316f
C3369 a_61358_58354# sar10b_0.net16 0.21268f
C3370 VDDD sar10b_0.net39 2.58664f
C3371 a_67445_60119# a_67881_60339# 0.16939f
C3372 c1_45456_54098# c1_45456_52978# 0.13255f
C3373 sar10b_0.net3 a_66933_55071# 0.22571f
C3374 VDDA a_n4470_65264# 1.65073f
C3375 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[0] 0.05999f
C3376 m3_n1472_26058# VDDR 0.02681f
C3377 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.02632f
C3378 a_64188_51135# sar10b_0.net16 0.10645f
C3379 VSSD a_60969_56639# 0.52879f
C3380 m3_n1472_33898# VCM 0.01415f
C3381 sar10b_0.net3 sar10b_0._14_ 0.03168f
C3382 c1_n1140_84532# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C3383 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN 0.01103f
C3384 m3_45124_55178# m3_45124_54058# 0.29566f
C3385 a_65577_57971# a_65966_58354# 0.06034f
C3386 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.02632f
C3387 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] m3_21120_21578# 0.26476f
C3388 a_62187_71265# VSSD 0.35653f
C3389 a_61065_53679# a_61249_53311# 0.43491f
C3390 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_36652_21578# 0.0162f
C3391 sar10b_0.net16 a_65761_58263# 0.12137f
C3392 sar10b_0.net32 sar10b_0._00_ 0.07229f
C3393 c1_38396_21618# VCM 0.01358f
C3394 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.01212f
C3395 VDDD a_61609_63602# 0.2072f
C3396 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 0.1901f
C3397 a_67297_55975# a_67502_56024# 0.09983f
C3398 a_67113_56343# a_68073_56343# 0.03471f
C3399 sar10b_0.SWN[3] sar10b_0.CF[3] 2.41793f
C3400 m3_n1472_66572# VDDR 0.02674f
C3401 tdc_0.OUTP VSSA 0.48683f
C3402 m3_n1472_74412# VCM 0.01412f
C3403 VDDD a_67209_65667# 0.9124f
C3404 a_63745_59971# a_64085_60119# 0.24088f
C3405 VDDD a_62037_61731# 0.30224f
C3406 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C3407 VSSD a_68169_66999# 0.29048f
C3408 sar10b_0.net9 sar10b_0.net8 0.3224f
C3409 VDDD a_62527_51646# 0.20742f
C3410 sar10b_0._01_ VSSD 0.31035f
C3411 a_64814_65014# sar10b_0.net12 0.02574f
C3412 sar10b_0.clknet_0_CLK sar10b_0.clknet_1_0__leaf_CLK 0.10604f
C3413 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A 1.29878f
C3414 VSSD a_66645_61731# 0.13981f
C3415 sar10b_0.net7 a_61833_57675# 0.23819f
C3416 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN 3.23431f
C3417 a_63169_62635# sar10b_0.net2 0.02592f
C3418 a_65001_68627# a_65185_68919# 0.44532f
C3419 VDDD a_65333_66248# 0.20416f
C3420 m3_n1472_22698# m3_n1472_21578# 0.29566f
C3421 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 a_5929_5779# 0.12755f
C3422 VSSR c1_n1140_48498# 0.04956f
C3423 sar10b_0.net34 a_66216_52022# 0.01157f
C3424 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 0.02632f
C3425 sar10b_0.CF[5] sar10b_0.SWP[0] 0.12716f
C3426 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 6.79685f
C3427 VSSR a_33863_5788# 0.06033f
C3428 a_61395_49960# sar10b_0.net6 0.21549f
C3429 sar10b_0.net16 a_61395_60616# 0.1993f
C3430 m3_45124_91212# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C3431 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VCM 0.12564f
C3432 sar10b_0.SWP[4] a_64491_71265# 0.1431f
C3433 m3_45124_95692# m3_45124_94572# 0.29566f
C3434 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 2.74732f
C3435 sar10b_0.CF[9] sar10b_0.CF[8] 65.7246f
C3436 sar10b_0.net4 sar10b_0.net6 0.05438f
C3437 sar10b_0.net34 a_65861_49313# 0.03738f
C3438 m3_32416_21578# c1_32748_21618# 1.74381f
C3439 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 sar10b_0.CF[2] 0.40679f
C3440 m3_45124_28298# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C3441 a_65778_49979# VSSD 1.1423f
C3442 a_65525_68912# sar10b_0.net43 0.01115f
C3443 a_249_5788# VSSR 0.06021f
C3444 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A 0.39559f
C3445 c1_39808_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26825f
C3446 m3_40888_97932# c1_41220_97972# 1.74381f
C3447 sar10b_0._15_ a_68276_50645# 0.09557f
C3448 a_62593_58639# sar10b_0.net8 0.02952f
C3449 VSSR m3_8412_21578# 0.53625f
C3450 sar10b_0.net6 a_62126_56024# 0.073f
C3451 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C3452 c1_25688_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.26825f
C3453 sar10b_0.net3 a_63918_50969# 0.02204f
C3454 VSSR a_44345_110521# 3.47951f
C3455 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y 0.12541f
C3456 sar10b_0.net3 a_66109_49318# 0.02012f
C3457 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] a_25137_112201# 0.68523f
C3458 a_61131_70891# VSSD 0.31867f
C3459 sar10b_0.net47 sar10b_0.net15 0.09931f
C3460 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 1.98252f
C3461 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.02632f
C3462 m3_2764_97932# VCM 0.15231f
C3463 a_65481_59303# sar10b_0.net14 0.01866f
C3464 sar10b_0.net16 a_63797_56924# 0.14316f
C3465 c1_32748_21618# th_dif_sw_0.VCN 0.13255f
C3466 VDDA sar10b_0.CF[3] 0.53372f
C3467 VDDD a_62837_61451# 0.20415f
C3468 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_24276_21618# 0.0106f
C3469 a_67209_55011# VSSD 0.51749f
C3470 m3_n1472_63212# m3_n1472_62092# 0.29566f
C3471 sar10b_0.net4 a_61493_67580# 0.05154f
C3472 a_61395_61948# a_61086_61974# 0.07766f
C3473 a_67372_52833# VSSD 0.21271f
C3474 a_68946_68627# VSSD 0.33163f
C3475 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A 0.02842f
C3476 m3_28180_21578# VCM 0.13579f
C3477 m3_7000_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C3478 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26364f
C3479 a_60690_54641# tdc_0.OUTN 0.28109f
C3480 sar10b_0.CF[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP 0.19336f
C3481 sar10b_0.clk_div_0.COUNT\[2\] sar10b_0.net35 0.02642f
C3482 m3_45124_80012# c1_45456_80052# 1.74381f
C3483 m3_n1472_78892# c1_n1140_80052# 0.01078f
C3484 m3_n1472_80012# c1_n1140_78932# 0.01078f
C3485 VSSR c1_45456_92372# 0.0935f
C3486 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A 0.04073f
C3487 a_67209_64335# sar10b_0.net3 0.1932f
C3488 sar10b_0.net3 sar10b_0.net29 0.01804f
C3489 m3_1352_97932# m3_2764_97932# 0.23959f
C3490 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A 0.60057f
C3491 c1_45456_26098# m3_45124_26058# 1.74381f
C3492 c1_n1140_24978# m3_n1472_26058# 0.01078f
C3493 c1_n1140_26098# m3_n1472_24938# 0.01078f
C3494 a_60945_65937# a_61400_66284# 0.3578f
C3495 a_66865_49412# sar10b_0.net35 0.02871f
C3496 sar10b_0.net33 sar10b_0.clknet_0_CLK 0.72841f
C3497 sar10b_0.CF[6] sar10b_0.SWP[3] 0.12147f
C3498 a_61677_52854# sar10b_0.net1 0.01783f
C3499 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 sar10b_0.CF[5] 0.40665f
C3500 VDDD a_62709_63063# 0.28745f
C3501 sar10b_0.net16 a_62017_57307# 0.11207f
C3502 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.04562f
C3503 c1_45456_76692# VDDR 0.01153f
C3504 VDDD sar10b_0.net11 2.38059f
C3505 m3_26768_21578# m3_28180_21578# 0.23959f
C3506 sar10b_0.net3 a_68325_56296# 0.17851f
C3507 VSSD sar10b_0.net35 1.12162f
C3508 sar10b_0.net38 a_64831_56974# 0.02492f
C3509 VSSR c1_45456_24978# 0.09348f
C3510 sar10b_0.net6 a_61557_57735# 0.02023f
C3511 a_63339_48621# VSSD 0.34105f
C3512 sar10b_0.SWP[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A 0.01506f
C3513 m3_n1472_66572# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C3514 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y 0.32264f
C3515 VSSR m3_43712_97932# 0.54637f
C3516 c1_45456_65492# c1_45456_64372# 0.13255f
C3517 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP a_14655_111306# 0.09439f
C3518 m3_43712_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.33071f
C3519 m3_n1472_41738# VDDR 0.02681f
C3520 VCM cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 4.06768f
C3521 a_61677_52854# a_62185_52707# 0.19065f
C3522 m3_n1472_49578# VCM 0.01415f
C3523 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN 3.77743f
C3524 a_61929_57971# VSSD 0.28605f
C3525 a_62593_58639# sar10b_0.net9 0.02511f
C3526 a_67393_58639# a_68169_59007# 0.3578f
C3527 a_60747_64605# a_60945_64605# 0.06623f
C3528 VSSR c1_21452_97972# 0.0466f
C3529 a_64814_65014# sar10b_0.net41 0.01424f
C3530 VDDD a_66049_69295# 0.23374f
C3531 a_63810_50901# VSSD 0.38398f
C3532 a_65761_58263# a_66789_58100# 0.07826f
C3533 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_14060_21578# 0.03017f
C3534 m3_22532_21578# th_dif_sw_0.VCN 0.01078f
C3535 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSSR 5.24147f
C3536 c1_11568_21618# VCM 0.01358f
C3537 sar10b_0.net30 a_61395_49960# 0.02544f
C3538 sar10b_0.net16 sar10b_0._12_ 0.02465f
C3539 a_65188_51977# sar10b_0.net16 0.08468f
C3540 m3_n1472_82252# VDDR 0.02674f
C3541 m3_n1472_90092# VCM 0.01412f
C3542 a_61395_65944# a_62185_66027# 0.1263f
C3543 sar10b_0.CF[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN 0.12367f
C3544 c1_n1140_29458# c1_n1140_28338# 0.13255f
C3545 a_63849_63299# sar10b_0.net2 0.01323f
C3546 a_62409_59007# VSSD 0.50378f
C3547 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A 0.42509f
C3548 sar10b_0.net4 a_61400_64952# 0.01899f
C3549 c1_41220_97972# VCM 0.01358f
C3550 m3_n1472_30538# m3_n1472_29418# 0.29566f
C3551 sar10b_0.SWN[7] VCM 0.13075f
C3552 sar10b_0.net13 a_61153_67587# 0.01352f
C3553 VSSR c1_n1140_67732# 0.04956f
C3554 a_60747_69559# VSSD 0.32872f
C3555 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 a_25137_112201# 0.4393f
C3556 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C3557 a_60747_64231# VSSD 0.32267f
C3558 a_65481_59303# sar10b_0.net13 0.0266f
C3559 a_61395_49960# VSSD 0.48695f
C3560 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.38072f
C3561 a_63339_48621# sar10b_0.net31 0.25741f
C3562 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 0.02632f
C3563 m3_22532_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.21489f
C3564 a_61358_51694# sar10b_0.net1 0.06982f
C3565 c1_45456_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C3566 sar10b_0.net4 VSSD 3.5209f
C3567 a_66795_71265# sar10b_0.net45 0.01175f
C3568 a_67209_64335# a_67598_64016# 0.05462f
C3569 a_62181_51440# a_61929_51311# 0.27388f
C3570 a_61153_51603# sar10b_0.net28 0.03795f
C3571 sar10b_0._07_ a_64454_51311# 0.16465f
C3572 a_66933_64395# a_67393_63967# 0.26257f
C3573 c1_18628_21618# m3_19708_21578# 0.15596f
C3574 th_dif_sw_0.CKB sar10b_0.CF[3] 0.17526f
C3575 VDDD a_61086_52650# 0.31199f
C3576 m3_45124_43978# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C3577 sar10b_0.net5 a_61153_56931# 0.02898f
C3578 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSSR 27.5188f
C3579 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] 1.04257f
C3580 sar10b_0.SWN[0] sar10b_0.CF[9] 0.84219f
C3581 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[1] 0.17717f
C3582 c1_272_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26825f
C3583 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] sar10b_0.SWP[6] 0.22722f
C3584 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A 0.74888f
C3585 m3_21120_97932# c1_21452_97972# 1.74381f
C3586 VSSD a_62126_56024# 0.13428f
C3587 VSSR m3_45124_33898# 0.63261f
C3588 a_64809_65963# a_65333_66248# 0.05022f
C3589 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR 2.50957f
C3590 sar10b_0.net3 a_67598_65348# 0.25604f
C3591 a_64910_59686# sar10b_0.net12 0.02444f
C3592 sar10b_0.SWN[6] VCM 0.13076f
C3593 a_68073_56343# VSSD 0.29128f
C3594 sar10b_0.net4 a_61400_60956# 0.01875f
C3595 VDDR a_33863_5788# 6.41271f
C3596 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSSR 6.85451f
C3597 VSSR c1_39808_21618# 0.05923f
C3598 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 3.28979f
C3599 a_60747_60609# a_61086_60642# 0.07649f
C3600 a_61395_60616# a_60945_60609# 0.03471f
C3601 a_68421_54964# a_68767_54656# 0.07649f
C3602 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN 0.01165f
C3603 m3_n1472_71052# m3_n1472_69932# 0.29566f
C3604 a_19457_5788# VSSR 0.06033f
C3605 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A 0.60057f
C3606 a_249_5788# VDDR 0.82898f
C3607 VSSR m3_45124_74412# 0.63305f
C3608 a_65765_50645# sar10b_0.net16 0.04396f
C3609 sar10b_0.net3 a_67564_50907# 0.02389f
C3610 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSSR 1.11457f
C3611 sar10b_0.net46 sar10b_0.net3 0.13252f
C3612 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP a_33863_107882# 0.19132f
C3613 m3_45124_87852# c1_45456_87892# 1.74381f
C3614 m3_n1472_86732# c1_n1140_87892# 0.01078f
C3615 m3_n1472_87852# c1_n1140_86772# 0.01078f
C3616 a_62313_61671# a_62497_61303# 0.44098f
C3617 a_68421_54964# sar10b_0.net37 0.02393f
C3618 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 2.66562f
C3619 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VDDR 2.56591f
C3620 VDDD sar10b_0.SWP[8] 0.41984f
C3621 sar10b_0._04_ a_66216_52022# 0.07634f
C3622 a_65682_51977# a_66865_52076# 0.0649f
C3623 a_65861_51977# a_66666_51977# 0.29221f
C3624 sar10b_0.net23 a_68169_63003# 0.01663f
C3625 c1_45456_33938# m3_45124_33898# 1.74381f
C3626 c1_n1140_33938# m3_n1472_32778# 0.01078f
C3627 c1_n1140_32818# m3_n1472_33898# 0.01078f
C3628 sar10b_0.net39 a_61677_64842# 0.02955f
C3629 sar10b_0.CF[4] sar10b_0.SWP[2] 0.12174f
C3630 sar10b_0.CF[5] sar10b_0.SWP[1] 0.12273f
C3631 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 3.25674f
C3632 CLK tdc_0.phase_detector_0.INN 0.03583f
C3633 VSSR a_33863_107882# 0.06033f
C3634 sar10b_0.SWP[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 0.42754f
C3635 sar10b_0.net1 a_62181_56768# 0.06421f
C3636 c1_24276_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.01445f
C3637 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.12068f
C3638 VDDD a_66213_68756# 0.27396f
C3639 a_67598_66680# a_67733_66779# 0.35559f
C3640 VCM sar10b_0.CF[7] 3.5074f
C3641 a_64033_63591# a_65061_63428# 0.07826f
C3642 a_63573_63303# a_64238_63682# 0.19065f
C3643 a_67231_56974# sar10b_0.net37 0.27502f
C3644 a_30644_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A 0.01076f
C3645 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 2.9143f
C3646 sar10b_0.net2 a_61153_56931# 0.03377f
C3647 VDDD a_66312_50368# 0.13937f
C3648 c1_45456_92372# VDDR 0.01153f
C3649 a_63621_58960# sar10b_0.net39 0.0805f
C3650 sar10b_0._11_ a_64780_52239# 0.12171f
C3651 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y 0.07183f
C3652 a_66825_69663# sar10b_0.net16 0.266f
C3653 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.36778f
C3654 m3_7000_21578# m3_8412_21578# 0.23959f
C3655 VSSD a_61557_57735# 0.13613f
C3656 VSSR c1_45456_40658# 0.09348f
C3657 sar10b_0.net2 sar10b_0.net40 0.99203f
C3658 CLK sar10b_0.net5 0.01289f
C3659 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR 0.36333f
C3660 VSSR a_39543_110941# 3.14203f
C3661 a_68767_58652# VSSD 0.26921f
C3662 m3_n1472_82252# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C3663 VSSR m3_4176_97932# 0.54637f
C3664 th_dif_sw_0.CK CLK 0.11183f
C3665 c1_45456_73332# c1_45456_72212# 0.13255f
C3666 sar10b_0.net16 a_60945_61941# 0.26608f
C3667 m3_43712_21578# c1_42632_21618# 0.15596f
C3668 m3_4176_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.53746f
C3669 sar10b_0.CF[1] sar10b_0.CF[0] 39.8486f
C3670 a_62185_63363# VSSD 0.15732f
C3671 sar10b_0.net39 a_61677_60846# 0.01935f
C3672 sar10b_0.clk_div_0.COUNT\[1\] sar10b_0._12_ 0.21887f
C3673 a_66865_52076# sar10b_0._07_ 0.04846f
C3674 a_64725_68631# VSSD 0.13754f
C3675 a_63797_56924# a_64233_56639# 0.16939f
C3676 a_62497_61303# a_62702_61352# 0.09983f
C3677 VSSR m3_29592_21578# 0.49843f
C3678 sar10b_0.net16 a_61086_65970# 0.18334f
C3679 sar10b_0._07_ a_64188_51135# 0.01836f
C3680 VSSD a_67393_65299# 0.8514f
C3681 sar10b_0.SWP[4] VDDA 0.2491f
C3682 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] sar10b_0.SWP[2] 0.23418f
C3683 VDDD a_67209_68331# 0.8941f
C3684 c1_45456_24978# VDDR 0.01151f
C3685 m3_45124_28298# th_dif_sw_0.VCN 0.17339f
C3686 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP 0.02666f
C3687 sar10b_0.net44 VSSD 1.74731f
C3688 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] a_5929_113881# 0.22044f
C3689 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A 0.05472f
C3690 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y 0.3196f
C3691 sar10b_0.CF[5] th_dif_sw_0.CK 0.17586f
C3692 VSSD a_66367_66298# 0.27123f
C3693 a_60789_53739# VSSD 0.13736f
C3694 sar10b_0.CF[1] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.01368f
C3695 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A 0.26294f
C3696 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C3697 sar10b_0.SWN[5] VCM 0.13075f
C3698 m3_23944_97932# VCM 0.13579f
C3699 c1_45456_56338# m3_45124_57418# 0.01078f
C3700 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_45456_21618# 0.0106f
C3701 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP a_5051_113018# 0.04592f
C3702 sar10b_0.net8 sar10b_0.net1 0.45568f
C3703 sar10b_0.net18 VSSD 0.89477f
C3704 sar10b_0.net19 a_68671_55988# 0.01991f
C3705 sar10b_0.SWP[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 0.27668f
C3706 c1_n1140_37298# c1_n1140_36178# 0.13255f
C3707 a_60747_60235# sar10b_0.CF[3] 0.14607f
C3708 a_69003_71265# VSSD 0.33076f
C3709 sar10b_0.clk_div_0.COUNT\[0\] a_65957_50273# 0.0645f
C3710 m3_28180_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C3711 c1_1684_97972# VCM 0.01358f
C3712 m3_n1472_38378# m3_n1472_37258# 0.29566f
C3713 a_65045_59588# sar10b_0.net1 0.05003f
C3714 VSSR c1_n1140_83412# 0.04956f
C3715 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR 2.96457f
C3716 sar10b_0.cyclic_flag_0.FINAL a_67113_56343# 0.23922f
C3717 sar10b_0.cyclic_flag_0.FINAL a_66933_67059# 0.05303f
C3718 sar10b_0.net38 sar10b_0.net2 0.53673f
C3719 c1_5920_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C3720 c1_n1140_21618# m3_n60_21578# 0.15596f
C3721 sar10b_0.net38 a_61609_66266# 0.0226f
C3722 a_64245_59307# sar10b_0.net12 0.01064f
C3723 VDDD sar10b_0.SWN[4] 0.19275f
C3724 VDDA VINP 0.87608f
C3725 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 0.38263f
C3726 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 5.16397f
C3727 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C3728 tdc_0.phase_detector_0.INN a_52417_59293# 0.10585f
C3729 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A 0.07418f
C3730 m3_1352_97932# c1_1684_97972# 1.74381f
C3731 VSSR m3_45124_49578# 0.63261f
C3732 c1_29924_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.26825f
C3733 VSSD a_63273_61671# 0.29931f
C3734 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A sar10b_0.SWN[0] 0.01417f
C3735 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] a_44345_110521# 1.14986f
C3736 sar10b_0.net16 a_66049_57307# 0.11922f
C3737 sar10b_0.net20 sar10b_0.net18 0.61871f
C3738 c1_n1140_26098# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C3739 VSSD sar10b_0.SWP[2] 0.98111f
C3740 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A 0.68875f
C3741 m3_14060_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C3742 VSSD a_63273_67295# 0.52636f
C3743 sar10b_0.net39 a_63391_57320# 0.02391f
C3744 VSSR c1_12980_21618# 0.05685f
C3745 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP 3.13736f
C3746 a_61833_57675# a_62793_57675# 0.03471f
C3747 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A 0.05472f
C3748 a_62017_57307# a_62357_57455# 0.24088f
C3749 VDDD sar10b_0.CF[0] 0.48185f
C3750 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VDDR 6.76175f
C3751 sar10b_0._14_ sar10b_0.clk_div_0.COUNT\[3\] 0.42361f
C3752 m3_n1472_78892# m3_n1472_77772# 0.29566f
C3753 a_64373_63584# sar10b_0.net16 0.17657f
C3754 VSSR m3_45124_90092# 0.63305f
C3755 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP a_34741_5779# 0.01488f
C3756 m3_45124_33898# VDDR 0.0103f
C3757 VDDD a_66921_61671# 0.8853f
C3758 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.38263f
C3759 a_61065_51015# sar10b_0.net16 0.19025f
C3760 sar10b_0.CF[1] VSSA 0.38195f
C3761 DATA[7] sar10b_0.net25 0.02654f
C3762 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR 3.26488f
C3763 a_65573_52937# a_66080_53027# 0.21226f
C3764 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 1.78633f
C3765 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 0.01132f
C3766 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.07418f
C3767 VSSR c1_42632_97972# 0.05923f
C3768 a_63374_62684# VSSD 0.14243f
C3769 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_18296_21578# 0.0162f
C3770 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_35240_21578# 0.03017f
C3771 m3_43712_21578# th_dif_sw_0.VCN 0.01078f
C3772 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VDDR 4.04887f
C3773 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A 0.03718f
C3774 a_64199_50761# VSSD 0.63836f
C3775 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 2.6566f
C3776 c1_20040_21618# VCM 0.01358f
C3777 c1_n1140_40658# m3_n1472_41738# 0.01078f
C3778 c1_n1140_41778# m3_n1472_40618# 0.01078f
C3779 c1_45456_41778# m3_45124_41738# 1.74381f
C3780 VDDD a_65021_50292# 0.22479f
C3781 a_19457_5788# VDDR 4.02021f
C3782 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A 0.01751f
C3783 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A 0.07183f
C3784 m3_45124_71052# th_dif_sw_0.VCP 0.17339f
C3785 m3_45124_74412# VDDR 0.01034f
C3786 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A 0.41861f
C3787 m3_22532_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.15113f
C3788 sar10b_0.net9 sar10b_0.net1 0.05521f
C3789 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VDDR 0.95194f
C3790 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN sar10b_0.CF[3] 0.10416f
C3791 sar10b_0._11_ VSSD 0.38537f
C3792 a_67084_53565# sar10b_0._16_ 0.2071f
C3793 sar10b_0.SWP[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.32591f
C3794 VDDD a_60690_70625# 0.40882f
C3795 a_67393_65299# a_68421_65620# 0.07826f
C3796 sar10b_0.SWP[3] sar10b_0.CF[7] 0.12518f
C3797 sar10b_0.SWP[2] sar10b_0.CF[8] 0.13046f
C3798 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VDDR 4.31516f
C3799 m3_45124_64332# c1_45456_63252# 0.01078f
C3800 m3_n1472_63212# c1_n1140_63252# 1.74381f
C3801 m3_45124_63212# c1_45456_64372# 0.01078f
C3802 VSSR c1_45456_56338# 0.09348f
C3803 sar10b_0.clknet_0_CLK sar10b_0._01_ 0.05362f
C3804 sar10b_0.net23 VSSD 0.88093f
C3805 a_51345_60437# a_51603_61205# 0.06738f
C3806 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A 0.10815f
C3807 a_68946_61735# sar10b_0.net22 0.01815f
C3808 m3_43712_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.33071f
C3809 VDDR a_33863_107882# 6.41271f
C3810 a_66837_56403# sar10b_0.net40 0.17432f
C3811 sar10b_0._08_ a_65021_50292# 0.0923f
C3812 m3_19708_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.18393f
C3813 sar10b_0.SWN[8] sar10b_0.CF[9] 0.13258f
C3814 m3_42300_97932# m3_43712_97932# 0.23959f
C3815 a_68421_64288# a_68767_63980# 0.07649f
C3816 c1_45456_81172# c1_45456_80052# 0.13255f
C3817 m3_23944_21578# c1_22864_21618# 0.15596f
C3818 VINN th_dif_sw_0.th_sw_1.CK 0.32523f
C3819 m3_n1472_35018# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C3820 VDDD a_66577_52883# 0.39116f
C3821 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 1.77469f
C3822 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 2.62902f
C3823 a_61249_50647# CLK 0.02421f
C3824 sar10b_0.CF[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 0.16034f
C3825 a_62181_56768# a_62527_56974# 0.07649f
C3826 a_61493_56924# a_61358_57022# 0.35559f
C3827 a_65865_69663# a_66049_69295# 0.43491f
C3828 VSSD a_60747_61941# 0.2587f
C3829 a_66153_48647# sar10b_0.SWN[7] 0.02069f
C3830 m3_32416_97932# c1_31336_97972# 0.15596f
C3831 VSSR m3_n1472_24938# 0.66371f
C3832 sar10b_0.clknet_0_CLK a_65778_49979# 0.05485f
C3833 a_61395_49960# a_61400_50300# 0.43491f
C3834 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.59327f
C3835 c1_35572_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26825f
C3836 c1_45456_40658# VDDR 0.01151f
C3837 sar10b_0.net7 sar10b_0.net38 0.0467f
C3838 m3_45124_43978# th_dif_sw_0.VCN 0.17339f
C3839 sar10b_0.SWP[5] a_65643_71265# 0.1431f
C3840 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR 0.59846f
C3841 a_67393_62635# a_68421_62956# 0.07826f
C3842 sar10b_0.net2 sar10b_0.net14 0.06252f
C3843 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.12357f
C3844 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN 3.06947f
C3845 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C3846 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.28117f
C3847 sar10b_0.net7 CLK 0.05137f
C3848 VDDD a_62623_53324# 0.21258f
C3849 sar10b_0.SWN[9] sar10b_0.CF[9] 2.43858f
C3850 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 0.24774f
C3851 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_18628_21618# 0.0106f
C3852 sar10b_0.net16 a_61929_56639# 0.32351f
C3853 a_65188_51977# sar10b_0._07_ 0.0214f
C3854 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A 0.43651f
C3855 VSSR m3_n1472_65452# 0.66316f
C3856 c1_n1140_45138# c1_n1140_44018# 0.13255f
C3857 sar10b_0.CF[8] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 0.01331f
C3858 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C3859 a_61609_52946# VSSD 0.09801f
C3860 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 a_44345_110521# 0.75105f
C3861 sar10b_0.SWN[6] a_66153_48647# 0.09312f
C3862 m3_9824_21578# VCM 0.13573f
C3863 sar10b_0.net6 a_61493_56924# 0.02599f
C3864 c1_n1140_67732# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C3865 sar10b_0.net3 sar10b_0.net42 0.13229f
C3866 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.1066f
C3867 m3_n1472_46218# m3_n1472_45098# 0.29566f
C3868 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN 0.01183f
C3869 m3_19708_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 0.48426f
C3870 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN sar10b_0.CF[7] 0.06919f
C3871 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y sar10b_0.CF[2] 0.12541f
C3872 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A 0.10815f
C3873 sar10b_0.net3 a_67598_68012# 0.23749f
C3874 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.22192f
C3875 sar10b_0.net38 a_66837_56403# 0.02722f
C3876 VDDD a_66216_52022# 0.1367f
C3877 VDDD a_68946_63299# 0.27896f
C3878 VDDD a_62181_58100# 0.27078f
C3879 sar10b_0.SWP[8] a_5051_113018# 0.22599f
C3880 a_68767_66644# sar10b_0.net26 0.27142f
C3881 a_61491_52222# a_62281_52347# 0.1263f
C3882 a_66921_60339# sar10b_0.net3 0.1825f
C3883 a_1127_5779# sar10b_0.SWN[9] 0.08773f
C3884 VDDD a_62623_50660# 0.20184f
C3885 a_60969_57971# a_61153_58263# 0.44532f
C3886 sar10b_0.CF[0] sar10b_0.CF[2] 0.12815f
C3887 VDDD a_65861_49313# 0.84101f
C3888 c1_n1140_41778# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C3889 a_61395_63280# sar10b_0.net40 0.01724f
C3890 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A 1.11704f
C3891 VCM EN 2.09751f
C3892 a_66921_61671# a_68133_61624# 0.07766f
C3893 a_67105_61303# a_67445_61451# 0.24088f
C3894 VSSR c1_n1140_31698# 0.04956f
C3895 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] a_10731_5779# 0.3365f
C3896 sar10b_0.net4 a_61454_53360# 0.07375f
C3897 a_66197_56924# a_66062_57022# 0.35559f
C3898 a_64583_51628# sar10b_0.net16 0.01266f
C3899 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] a_9853_112162# 0.88621f
C3900 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 2.48625f
C3901 sar10b_0.clknet_0_CLK sar10b_0.net35 0.17355f
C3902 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.02842f
C3903 m3_45124_74412# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C3904 a_62181_67424# sar10b_0.net40 0.02383f
C3905 m3_n1472_86732# m3_n1472_85612# 0.29566f
C3906 VSSR m3_25356_97932# 0.44647f
C3907 sar10b_0.net34 sar10b_0.net40 0.37914f
C3908 sar10b_0._10_ a_65573_52937# 0.01418f
C3909 sar10b_0.cyclic_flag_0.FINAL a_67135_58306# 0.01523f
C3910 m3_25356_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.27266f
C3911 a_64609_64923# sar10b_0.net42 0.01976f
C3912 m3_45124_49578# VDDR 0.0103f
C3913 a_60747_52617# a_61086_52650# 0.07649f
C3914 sar10b_0.net29 a_61035_48621# 0.28332f
C3915 a_61395_52624# a_60945_52617# 0.03529f
C3916 VDDD a_68946_71059# 0.2715f
C3917 a_60969_67295# sar10b_0.net16 0.17797f
C3918 VDDD a_60747_49953# 0.22619f
C3919 VSSR c1_3096_97972# 0.05923f
C3920 a_65733_59432# sar10b_0.net16 0.21131f
C3921 sar10b_0.cyclic_flag_0.FINAL VSSD 3.91093f
C3922 a_67733_62783# sar10b_0.net3 0.16914f
C3923 VDDD a_60693_67299# 0.33734f
C3924 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A sar10b_0.CF[3] 0.06369f
C3925 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VDDR 3.03881f
C3926 sar10b_0.net39 sar10b_0.net12 0.06377f
C3927 sar10b_0.SWP[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 0.48483f
C3928 a_62997_56643# a_63662_57022# 0.19065f
C3929 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26364f
C3930 c1_n1140_48498# m3_n1472_49578# 0.01078f
C3931 c1_n1140_49618# m3_n1472_48458# 0.01078f
C3932 c1_45456_49618# m3_45124_49578# 1.74381f
C3933 c1_n1140_95732# c1_n1140_94612# 0.13255f
C3934 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A sar10b_0.CF[5] 0.02149f
C3935 a_63273_67295# a_64492_67433# 0.07276f
C3936 VSSR sar10b_0.SWP[8] 3.53937f
C3937 m3_45124_90092# VDDR 0.01034f
C3938 m3_45124_86732# th_dif_sw_0.VCP 0.17339f
C3939 VDDD a_68479_59984# 0.21268f
C3940 VDDD a_61921_55975# 0.2263f
C3941 m3_45124_97932# VCM 0.15686f
C3942 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 0.02632f
C3943 a_67890_69727# sar10b_0.net15 0.14196f
C3944 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] m3_22532_21578# 0.53272f
C3945 sar10b_0.net10 sar10b_0.net2 0.53489f
C3946 sar10b_0._09_ CLK 0.05323f
C3947 a_65928_53032# a_65821_53072# 0.14439f
C3948 sar10b_0.net2 sar10b_0.net13 0.03037f
C3949 sar10b_0.CF[1] th_dif_sw_0.VCN 0.28956f
C3950 a_64491_71265# VSSD 0.36767f
C3951 c1_22864_97972# VCM 0.01162f
C3952 sar10b_0._03_ a_65957_50273# 0.3098f
C3953 sar10b_0.net28 a_61609_50282# 0.01541f
C3954 a_64085_60119# sar10b_0.net16 0.14879f
C3955 w_n9655_63119# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 0.99238f
C3956 sar10b_0.net3 a_67105_61303# 0.13379f
C3957 m3_45124_72172# c1_45456_71092# 0.01078f
C3958 m3_n1472_71052# c1_n1140_71092# 1.74381f
C3959 m3_45124_71052# c1_45456_72212# 0.01078f
C3960 VSSR c1_45456_75572# 0.0935f
C3961 a_19457_110450# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 0.4985f
C3962 m3_4176_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.53746f
C3963 sar10b_0.net39 a_63662_57022# 0.01259f
C3964 sar10b_0.CF[4] a_60747_61567# 0.14807f
C3965 c1_27100_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C3966 a_67393_67963# VSSD 0.85045f
C3967 m3_22532_97932# m3_23944_97932# 0.23959f
C3968 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 0.02666f
C3969 c1_10156_21618# m3_9824_21578# 1.74381f
C3970 c1_45456_89012# c1_45456_87892# 0.13255f
C3971 m3_n1472_50698# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C3972 a_65045_59588# a_65481_59303# 0.16939f
C3973 sar10b_0.net34 sar10b_0.net38 0.23791f
C3974 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.36779f
C3975 m3_12648_97932# c1_11568_97972# 0.15596f
C3976 a_60969_51311# CLK 0.01964f
C3977 m3_45124_57418# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C3978 VSSR m3_n1472_40618# 0.66371f
C3979 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 0.01864f
C3980 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_26878_111642# 0.01076f
C3981 sar10b_0.net47 a_66933_68391# 0.22592f
C3982 sar10b_0.clk_div_0.COUNT\[0\] a_68276_50645# 0.11059f
C3983 c1_8744_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.28115f
C3984 a_65765_50645# a_66103_50668# 0.21601f
C3985 a_65586_50645# a_65996_50650# 0.07154f
C3986 c1_45456_56338# VDDR 0.01151f
C3987 VSSA sar10b_0.CF[2] 0.36958f
C3988 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[2] 0.05939f
C3989 m3_35240_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C3990 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 0.62612f
C3991 VSSR c1_21452_21618# 0.0466f
C3992 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26364f
C3993 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] c1_22864_97972# 0.01334f
C3994 sar10b_0.clk_div_0.COUNT\[1\] sar10b_0.net16 0.0192f
C3995 VSSR m3_n1472_81132# 0.66316f
C3996 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] a_29061_108738# 2.08782f
C3997 c1_n1140_52978# c1_n1140_51858# 0.13255f
C3998 sar10b_0.net38 a_66197_56924# 0.02083f
C3999 a_68331_52243# sar10b_0.net37 0.02342f
C4000 m3_n1472_24938# VDDR 0.02681f
C4001 a_61737_56343# a_61461_56403# 0.1263f
C4002 VSSD a_61493_56924# 0.09868f
C4003 m3_n1472_32778# VCM 0.01415f
C4004 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A 0.11547f
C4005 VDDD a_61833_57675# 0.84068f
C4006 c1_n1140_83412# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C4007 m3_n1472_54058# m3_n1472_52938# 0.29566f
C4008 sar10b_0.CF[5] tdc_0.OUTP 0.15687f
C4009 a_67598_62684# VSSD 0.13556f
C4010 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSSR 2.45476f
C4011 VDDD a_68421_58960# 0.27526f
C4012 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A 0.07418f
C4013 sar10b_0.net16 a_60945_64605# 0.29236f
C4014 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A VSSR 0.39674f
C4015 a_60789_53739# a_61454_53360# 0.19065f
C4016 a_61065_53679# a_61589_53459# 0.04522f
C4017 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_39476_21578# 0.0162f
C4018 sar10b_0.net16 a_66789_58100# 0.17399f
C4019 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[2] 0.17717f
C4020 c1_41220_21618# VCM 0.01358f
C4021 a_67502_56024# a_67637_56123# 0.35559f
C4022 m3_n1472_65452# VDDR 0.02674f
C4023 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A 0.38427f
C4024 m3_n1472_62092# th_dif_sw_0.VCP 0.12457f
C4025 sar10b_0._04_ a_68943_51605# 0.01727f
C4026 a_43467_5788# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 1.02702f
C4027 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VCM 0.12358f
C4028 c1_18628_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.02523f
C4029 m3_n1472_73292# VCM 0.01412f
C4030 a_62798_58688# sar10b_0.net16 0.22368f
C4031 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.43651f
C4032 sar10b_0.net28 a_62187_48621# 0.03427f
C4033 sar10b_0.SWN[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP 0.28712f
C4034 a_65407_63634# sar10b_0.net13 0.01616f
C4035 a_65397_56643# a_65857_56931# 0.26257f
C4036 sar10b_0.CF[4] sar10b_0.SWN[3] 0.11956f
C4037 VSSD a_68767_66644# 0.26637f
C4038 VSSR sar10b_0.SWN[4] 4.86208f
C4039 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR 0.95734f
C4040 c1_n1140_57458# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C4041 sar10b_0.clknet_1_1__leaf_CLK sar10b_0.clknet_1_0__leaf_CLK 0.07504f
C4042 a_67696_52265# a_67651_51991# 0.01224f
C4043 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.32324f
C4044 sar10b_0.CF[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP 0.1053f
C4045 VDDD a_66795_71265# 0.26692f
C4046 a_63509_62783# sar10b_0.net2 0.0256f
C4047 sar10b_0.CF[0] tdc_0.OUTN 0.2561f
C4048 a_65001_68627# a_66213_68756# 0.07766f
C4049 VDDD a_65769_65963# 0.36939f
C4050 a_65185_68919# a_65525_68912# 0.24088f
C4051 VDDD a_61065_53679# 0.82448f
C4052 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A 0.01751f
C4053 sar10b_0.SWP[5] VDDD 0.47059f
C4054 VSSR c1_n1140_47378# 0.04956f
C4055 sar10b_0.net34 a_66666_51977# 0.01385f
C4056 sar10b_0.net16 a_60945_60609# 0.26406f
C4057 m3_45124_90092# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C4058 a_65957_50273# a_66464_50363# 0.21226f
C4059 m3_n1472_94572# m3_n1472_93452# 0.29566f
C4060 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 sar10b_0.CF[4] 0.26311f
C4061 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.12357f
C4062 sar10b_0.net16 a_62697_56343# 0.26291f
C4063 m3_33828_21578# c1_34160_21618# 1.74381f
C4064 a_64454_51311# VSSD 0.41349f
C4065 m3_45124_27178# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C4066 VSSR sar10b_0.CF[0] 16.8353f
C4067 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN 3.19421f
C4068 c1_42632_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26825f
C4069 a_66825_69663# a_67423_69308# 0.06623f
C4070 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VDDR 0.95141f
C4071 m3_42300_97932# c1_42632_97972# 1.74381f
C4072 sar10b_0.net3 a_67372_52243# 0.01678f
C4073 VSSD a_60747_61567# 0.32213f
C4074 a_n8277_65767# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 1.59491f
C4075 a_62933_58787# sar10b_0.net8 0.01008f
C4076 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.43651f
C4077 VSSR m3_11236_21578# 0.49843f
C4078 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C4079 a_65390_69010# sar10b_0.net16 0.22679f
C4080 sar10b_0.net3 a_66216_49358# 0.04082f
C4081 a_64705_59595# VSSD 0.86334f
C4082 c1_n1140_57458# m3_n1472_56298# 0.01078f
C4083 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 3.04082f
C4084 VSSR cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.31308p
C4085 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.40463f
C4086 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.41774f
C4087 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y sar10b_0.CF[1] 0.12541f
C4088 a_68235_48621# sar10b_0.net35 0.30633f
C4089 m3_5588_97932# VCM 0.15231f
C4090 sar10b_0.net16 a_64233_56639# 0.26f
C4091 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_27100_21618# 0.0106f
C4092 m3_45124_63212# m3_45124_62092# 0.29566f
C4093 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] sar10b_0.SWP[9] 0.22372f
C4094 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN sar10b_0.SWN[7] 0.20215f
C4095 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A sar10b_0.CF[8] 0.02149f
C4096 sar10b_0.net4 a_61929_67295# 0.09064f
C4097 a_60945_61941# a_61400_62288# 0.3578f
C4098 sar10b_0.CF[4] VDDA 0.50636f
C4099 m3_31004_21578# VCM 0.13579f
C4100 m3_9824_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C4101 m3_n1472_78892# c1_n1140_78932# 1.74381f
C4102 m3_45124_80012# c1_45456_78932# 0.01078f
C4103 m3_45124_78892# c1_45456_80052# 0.01078f
C4104 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y 0.32296f
C4105 VSSR c1_45456_91252# 0.0935f
C4106 a_68331_52243# sar10b_0._03_ 0.14196f
C4107 sar10b_0.net24 a_68946_61735# 0.26084f
C4108 sar10b_0.SWP[8] VDDR 1.22823f
C4109 a_63745_59971# VSSD 0.883f
C4110 VSSD a_65397_56643# 0.14151f
C4111 m3_2764_97932# m3_4176_97932# 0.23959f
C4112 a_64425_64631# a_64609_64923# 0.44532f
C4113 c1_45456_26098# m3_45124_24938# 0.01078f
C4114 c1_45456_24978# m3_45124_26058# 0.01078f
C4115 c1_n1140_24978# m3_n1472_24938# 1.74381f
C4116 sar10b_0.net40 a_62793_57675# 0.0546f
C4117 a_60945_65937# a_61609_66266# 0.16939f
C4118 sar10b_0.net33 sar10b_0.clknet_1_1__leaf_CLK 0.20395f
C4119 a_63745_59971# a_63561_60339# 0.44098f
C4120 a_62185_52707# sar10b_0.net1 0.013f
C4121 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 a_1127_114301# 0.04962f
C4122 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C4123 a_66865_52076# sar10b_0.clk_div_0.COUNT\[2\] 0.12382f
C4124 a_67372_52243# a_67798_52206# 0.16025f
C4125 sar10b_0.clk_div_0.COUNT\[1\] a_67696_52265# 0.01064f
C4126 VDDD a_63169_62635# 0.22075f
C4127 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 3.62378f
C4128 sar10b_0.net21 sar10b_0.net3 0.22182f
C4129 VSSR m3_n1472_56298# 0.66371f
C4130 sar10b_0.net16 a_62357_57455# 0.14709f
C4131 sar10b_0.CF[6] sar10b_0.net11 0.01224f
C4132 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A 0.05472f
C4133 a_61035_71265# sar10b_0.net39 0.25439f
C4134 c1_45456_75572# VDDR 0.01153f
C4135 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A 1.11704f
C4136 m3_28180_21578# m3_29592_21578# 0.23959f
C4137 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 0.62612f
C4138 VSSA tdc_0.OUTN 1.44534f
C4139 VSSR c1_45456_23858# 0.09348f
C4140 sar10b_0.SWN[3] VSSD 1.61912f
C4141 sar10b_0.SWP[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A 0.01453f
C4142 m3_n1472_65452# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C4143 sar10b_0.SWP[8] sar10b_0.SWP[7] 19.5366f
C4144 VSSR m3_n1472_96812# 0.66316f
C4145 sar10b_0.net18 sar10b_0.SWN[8] 0.0794f
C4146 c1_n1140_64372# c1_n1140_63252# 0.13255f
C4147 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.59327f
C4148 a_64149_64635# VSSD 0.18148f
C4149 a_65643_71265# sar10b_0.SWP[6] 0.01261f
C4150 VDDD sar10b_0.net32 2.01563f
C4151 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.36422f
C4152 m3_n1472_40618# VDDR 0.02681f
C4153 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM 3.13305f
C4154 VSSR VSSA 30.3976f
C4155 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.10847f
C4156 m3_n1472_48458# VCM 0.01415f
C4157 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 0.22396f
C4158 a_66865_52076# VSSD 0.33239f
C4159 a_60747_62899# VSSD 0.32267f
C4160 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A 0.39674f
C4161 a_61358_58354# VSSD 0.13462f
C4162 a_67733_58787# a_68169_59007# 0.16939f
C4163 a_65637_64760# sar10b_0.net14 0.0247f
C4164 a_61395_64612# a_61086_64638# 0.07766f
C4165 VSSR c1_24276_97972# 0.05929f
C4166 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A 0.10815f
C4167 a_65861_51977# a_65577_51311# 0.01795f
C4168 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] sar10b_0.SWN[6] 0.22719f
C4169 a_64188_51135# VSSD 1.172f
C4170 a_64197_62956# sar10b_0.net42 0.01341f
C4171 VDDD a_66389_69443# 0.20837f
C4172 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A VSSR 0.39656f
C4173 a_66101_58256# a_66537_57971# 0.16939f
C4174 a_68946_52411# DATA[2] 0.14249f
C4175 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_n60_21578# 0.01492f
C4176 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_16884_21578# 0.03017f
C4177 th_dif_sw_0.VCN sar10b_0.CF[2] 0.29716f
C4178 a_66368_49417# VSSD 0.14034f
C4179 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C4180 c1_14392_21618# VCM 0.01358f
C4181 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN sar10b_0.CF[7] 0.12367f
C4182 VSSD a_60747_64605# 0.2587f
C4183 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM 2.04843f
C4184 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] a_39543_110941# 1.0337f
C4185 a_61400_63620# a_61677_63510# 0.09983f
C4186 m3_n1472_81132# VDDR 0.02674f
C4187 sar10b_0._07_ sar10b_0.net16 0.40533f
C4188 VSSD a_65761_58263# 0.85595f
C4189 m3_n1472_88972# VCM 0.01412f
C4190 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 0.24771f
C4191 sar10b_0.net18 sar10b_0.SWN[9] 0.03171f
C4192 sar10b_0.net9 a_61086_60642# 0.04521f
C4193 sar10b_0.net32 sar10b_0._08_ 0.03114f
C4194 c1_45456_29458# c1_45456_28338# 0.13255f
C4195 a_60789_51075# sar10b_0.net1 0.17638f
C4196 a_62409_59007# a_63369_59007# 0.03471f
C4197 a_62593_58639# a_62933_58787# 0.24088f
C4198 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VDDR 2.40255f
C4199 c1_44044_97972# VCM 0.01358f
C4200 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.36778f
C4201 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A VDDR 0.60103f
C4202 m3_45124_30538# m3_45124_29418# 0.29566f
C4203 a_64780_52239# a_65188_51977# 0.08493f
C4204 DATA[3] sar10b_0.net36 0.10413f
C4205 VSSR c1_n1140_66612# 0.04956f
C4206 a_66933_64395# VSSD 0.13693f
C4207 a_62313_61671# a_62037_61731# 0.1263f
C4208 sar10b_0.SWN[3] sar10b_0.net31 0.01009f
C4209 sar10b_0.SWN[3] sar10b_0.CF[8] 0.12682f
C4210 m3_25356_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.27266f
C4211 sar10b_0._14_ sar10b_0._04_ 0.47505f
C4212 a_61929_51311# a_62527_51646# 0.06623f
C4213 a_62181_51440# sar10b_0.net28 0.04563f
C4214 m3_45124_42858# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C4215 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.38427f
C4216 VSSD a_61395_60616# 0.49262f
C4217 VDDR sar10b_0.SWN[4] 2.46652f
C4218 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] sar10b_0.CF[7] 0.01386f
C4219 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 6.30914f
C4220 c1_3096_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26825f
C4221 m3_22532_97932# c1_22864_97972# 1.74381f
C4222 m3_n1472_96812# c1_n1140_97972# 0.01078f
C4223 sar10b_0.CF[4] th_dif_sw_0.CKB 0.08567f
C4224 m3_n1472_97932# c1_n1140_96852# 0.01078f
C4225 a_64993_66255# a_65333_66248# 0.24088f
C4226 sar10b_0.net16 a_63457_67583# 0.10758f
C4227 a_64809_65963# a_65769_65963# 0.03432f
C4228 VSSR m3_45124_32778# 0.63261f
C4229 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.31983f
C4230 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] 3.24823f
C4231 sar10b_0.net2 sar10b_0.net42 2.44266f
C4232 sar10b_0.net46 sar10b_0.net45 0.72044f
C4233 a_68562_71291# sar10b_0.net15 0.25929f
C4234 sar10b_0.CF[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 0.26311f
C4235 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A sar10b_0.CF[1] 0.26294f
C4236 a_64521_59303# a_64910_59686# 0.06034f
C4237 a_68671_55988# VSSD 0.26806f
C4238 a_67209_63003# a_66933_63063# 0.1263f
C4239 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.38989f
C4240 VSSR c1_42632_21618# 0.05923f
C4241 m3_45124_57418# th_dif_sw_0.VCN 0.34926f
C4242 a_61395_60616# a_61400_60956# 0.44098f
C4243 sar10b_0.net16 a_60693_56643# 0.20257f
C4244 a_66049_57307# a_66389_57455# 0.24088f
C4245 a_65865_57675# a_67077_57628# 0.07766f
C4246 VDDR sar10b_0.CF[0] 1.6915f
C4247 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_272_21618# 0.01819f
C4248 a_61419_71265# th_dif_sw_0.CK 0.1421f
C4249 sar10b_0.SWP[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.01506f
C4250 m3_45124_71052# m3_45124_69932# 0.29566f
C4251 VSSR m3_45124_73292# 0.63305f
C4252 m3_18296_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 0.32786f
C4253 a_66103_50668# sar10b_0.net16 0.0276f
C4254 a_63945_63003# sar10b_0.net16 0.29525f
C4255 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.38427f
C4256 VSSD a_63797_56924# 0.11274f
C4257 VDDD a_65589_57735# 0.30352f
C4258 a_33863_5788# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.81562f
C4259 m3_45124_86732# c1_45456_87892# 0.01078f
C4260 m3_n1472_86732# c1_n1140_86772# 1.74381f
C4261 m3_45124_87852# c1_45456_86772# 0.01078f
C4262 a_62313_61671# a_62837_61451# 0.04522f
C4263 a_62037_61731# a_62702_61352# 0.19065f
C4264 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VSSR 1.99065f
C4265 sar10b_0.CF[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP 0.16026f
C4266 VDDR cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 16.0474f
C4267 sar10b_0._04_ a_66666_51977# 0.02332f
C4268 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38377f
C4269 sar10b_0.net23 a_68767_62648# 0.02711f
C4270 c1_45456_33938# m3_45124_32778# 0.01078f
C4271 c1_n1140_32818# m3_n1472_32778# 1.74381f
C4272 c1_45456_32818# m3_45124_33898# 0.01078f
C4273 VDDA sar10b_0.CF[8] 0.39322f
C4274 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A 0.06369f
C4275 th_dif_sw_0.th_sw_1.CK a_n8277_66083# 0.05367f
C4276 a_68671_55988# sar10b_0.net20 0.27386f
C4277 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 31.0559f
C4278 VDDD a_63849_63299# 0.84598f
C4279 a_249_113874# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.28719f
C4280 a_65637_64760# sar10b_0.net13 0.01959f
C4281 sar10b_0.net1 a_62527_56974# 0.05836f
C4282 c1_27100_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.01078f
C4283 VDDD a_66559_68962# 0.20582f
C4284 a_67393_66631# a_68169_66999# 0.3578f
C4285 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[0] 0.01902f
C4286 a_64373_63584# a_64809_63299# 0.16939f
C4287 sar10b_0.net2 a_62181_56768# 0.0162f
C4288 VDDD a_67439_50041# 0.34648f
C4289 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR 1.10847f
C4290 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y 0.31995f
C4291 c1_45456_91252# VDDR 0.01153f
C4292 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A VSSR 0.43773f
C4293 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] th_dif_sw_0.VCP 35.0616f
C4294 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26364f
C4295 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 0.02632f
C4296 m3_8412_21578# m3_9824_21578# 0.23959f
C4297 VSSD a_62017_57307# 0.82881f
C4298 VSSR c1_45456_39538# 0.09348f
C4299 sar10b_0.net34 a_65586_50645# 0.01632f
C4300 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 a_39543_110941# 0.67311f
C4301 a_19457_5788# sar10b_0.SWN[5] 0.5431f
C4302 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[7] 0.17717f
C4303 sar10b_0.net16 a_60945_49953# 0.27325f
C4304 c1_n1140_57458# th_dif_sw_0.VCN 0.02482f
C4305 m3_n1472_81132# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C4306 sar10b_0.net4 a_61491_52222# 0.2442f
C4307 VSSR m3_7000_97932# 0.54637f
C4308 c1_n1140_72212# c1_n1140_71092# 0.13255f
C4309 sar10b_0.net16 a_61400_62288# 0.10356f
C4310 m3_45124_21578# c1_44044_21618# 0.15596f
C4311 m3_7000_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.53769f
C4312 m3_n1472_56298# VDDR 0.02681f
C4313 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C4314 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.42811f
C4315 a_64485_56768# a_64831_56974# 0.07649f
C4316 a_63797_56924# sar10b_0.net31 0.03921f
C4317 a_62702_61352# a_62837_61451# 0.35559f
C4318 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A 0.9514f
C4319 VSSR m3_32416_21578# 0.49843f
C4320 VSSD a_67733_65447# 0.09956f
C4321 sar10b_0.net10 a_63285_60399# 0.05049f
C4322 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN 0.0121f
C4323 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.38218f
C4324 c1_45456_23858# VDDR 0.01151f
C4325 m3_45124_27178# th_dif_sw_0.VCN 0.17339f
C4326 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 30.4789f
C4327 th_dif_sw_0.CKB VSSD 0.93771f
C4328 sar10b_0.clknet_0_CLK a_66205_50408# 0.01988f
C4329 m3_n1472_96812# VDDR 0.02674f
C4330 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A 1.33999f
C4331 VDDD a_66062_57022# 0.26152f
C4332 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.59835f
C4333 m3_26768_97932# VCM 0.13579f
C4334 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A 0.39674f
C4335 VDDR VSSA 0.30426f
C4336 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.95198f
C4337 sar10b_0._12_ VSSD 0.2965f
C4338 c1_45456_37298# c1_45456_36178# 0.13255f
C4339 a_65188_51977# VSSD 0.02184f
C4340 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A 0.60103f
C4341 c1_32748_97972# th_dif_sw_0.VCP 0.13255f
C4342 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 0.20254f
C4343 a_67310_60020# sar10b_0.cyclic_flag_0.FINAL 0.05298f
C4344 sar10b_0.net47 sar10b_0.net44 0.0384f
C4345 VSSR th_dif_sw_0.VCN 0.11976p
C4346 sar10b_0.clk_div_0.COUNT\[0\] a_66312_50368# 0.03147f
C4347 c1_4508_97972# VCM 0.01358f
C4348 sar10b_0.net2 sar10b_0.net8 0.06408f
C4349 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 0.02632f
C4350 sar10b_0.SWN[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 0.35085f
C4351 m3_31004_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C4352 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A VDDR 0.6007f
C4353 m3_45124_38378# m3_45124_37258# 0.29566f
C4354 VSSR c1_n1140_82292# 0.04956f
C4355 m3_16884_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.66386f
C4356 a_66785_50875# sar10b_0.net35 0.03184f
C4357 VCM cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 7.03045f
C4358 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.02638f
C4359 sar10b_0.SWP[5] VSSR 4.48811f
C4360 c1_8744_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C4361 sar10b_0.clknet_1_0__leaf_CLK a_66153_48647# 1.88869f
C4362 a_62702_61352# sar10b_0.net11 0.01244f
C4363 sar10b_0.CF[6] sar10b_0.SWN[4] 0.12042f
C4364 sar10b_0.CF[1] CLK 0.18347f
C4365 c1_272_21618# m3_1352_21578# 0.15596f
C4366 sar10b_0.net40 a_66825_57675# 0.047f
C4367 VDDD a_61153_56931# 0.26578f
C4368 a_64245_59307# a_64521_59303# 0.1263f
C4369 VDDD sar10b_0.SWP[6] 2.02726f
C4370 a_68331_52243# sar10b_0._13_ 0.26661f
C4371 sar10b_0.SWP[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.47058f
C4372 VDDD a_67393_62635# 0.24951f
C4373 m3_2764_97932# c1_3096_97972# 1.74381f
C4374 VSSR m3_45124_48458# 0.63261f
C4375 c1_32748_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.01078f
C4376 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.59327f
C4377 VSSD a_63871_61316# 0.29132f
C4378 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN 0.01212f
C4379 a_67393_67963# a_68421_68284# 0.07826f
C4380 VDDD sar10b_0.net40 2.23413f
C4381 sar10b_0.net16 a_66389_57455# 0.15565f
C4382 c1_n1140_24978# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C4383 m3_16884_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C4384 a_62985_63003# a_62709_63063# 0.1263f
C4385 sar10b_0.CF[6] sar10b_0.CF[0] 0.11672f
C4386 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN 0.02638f
C4387 sar10b_0.CF[5] sar10b_0.CF[1] 0.1135f
C4388 VSSR c1_15804_21618# 0.06681f
C4389 th_dif_sw_0.CKB sar10b_0.CF[8] 0.08862f
C4390 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A 0.05472f
C4391 VDDD a_68421_66952# 0.27523f
C4392 a_62985_63003# sar10b_0.net11 0.01652f
C4393 a_64809_63299# sar10b_0.net16 0.27209f
C4394 m3_45124_78892# m3_45124_77772# 0.29566f
C4395 VSSR m3_45124_88972# 0.63305f
C4396 a_66921_60339# a_67105_59971# 0.44098f
C4397 tdc_0.phase_detector_0.INN a_53564_60302# 0.01732f
C4398 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 8.01941f
C4399 sar10b_0.SWN[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN 0.22816f
C4400 m3_45124_32778# VDDR 0.0103f
C4401 a_66080_53027# a_65928_53032# 0.22517f
C4402 a_65573_52937# a_66577_52883# 0.06302f
C4403 a_65765_50645# VSSD 0.55875f
C4404 VSSR c1_45456_97972# 0.11546f
C4405 sar10b_0.clknet_1_0__leaf_CLK a_65957_50273# 0.01206f
C4406 a_62185_64695# sar10b_0.net11 0.17016f
C4407 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR 1.10847f
C4408 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_21120_21578# 0.0162f
C4409 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_38064_21578# 0.03017f
C4410 a_64356_51029# VSSD 0.18166f
C4411 VDDD a_64339_51661# 0.24865f
C4412 c1_22864_21618# VCM 0.01162f
C4413 c1_45456_41778# m3_45124_40618# 0.01078f
C4414 c1_n1140_40658# m3_n1472_40618# 1.74381f
C4415 c1_45456_40658# m3_45124_41738# 0.01078f
C4416 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP 0.02666f
C4417 a_67393_58639# sar10b_0.cyclic_flag_0.FINAL 0.08047f
C4418 m3_45124_69932# th_dif_sw_0.VCP 0.17339f
C4419 m3_45124_73292# VDDR 0.01034f
C4420 m3_25356_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.19539f
C4421 a_64425_64631# sar10b_0.net2 0.01178f
C4422 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 a_34741_5779# 0.59518f
C4423 sar10b_0.net9 sar10b_0.net2 0.78215f
C4424 sar10b_0.net33 a_66153_48647# 0.01691f
C4425 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VDDR 2.56431f
C4426 VDDD sar10b_0.net38 5.52904f
C4427 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 2.76511f
C4428 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP 5.97231f
C4429 m3_n1472_63212# c1_n1140_62132# 0.01078f
C4430 m3_45124_63212# c1_45456_63252# 1.74381f
C4431 m3_n1472_62092# c1_n1140_63252# 0.01078f
C4432 sar10b_0.clknet_1_1__leaf_CLK sar10b_0._01_ 0.19733f
C4433 VSSR c1_45456_55218# 0.09226f
C4434 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 0.68875f
C4435 a_65682_51977# sar10b_0._07_ 0.17031f
C4436 VDDD CLK 1.14499f
C4437 sar10b_0._08_ a_64339_51661# 0.03659f
C4438 VDDD a_66933_55071# 0.32719f
C4439 a_66825_69663# VSSD 0.28884f
C4440 m3_n1472_96812# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C4441 m3_22532_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.15113f
C4442 VCM sar10b_0.CF[9] 3.48271f
C4443 m3_43712_97932# m3_45124_97932# 0.23959f
C4444 c1_n1140_80052# c1_n1140_78932# 0.13255f
C4445 m3_25356_21578# c1_24276_21618# 0.15596f
C4446 VSSA a_51345_60437# 0.48384f
C4447 a_62025_53679# a_62277_53632# 0.27388f
C4448 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 4.60179f
C4449 m3_n1472_33898# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C4450 VDDD sar10b_0._14_ 0.648f
C4451 VSSD a_60747_60235# 0.32798f
C4452 a_61589_50795# CLK 0.01091f
C4453 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR 0.95198f
C4454 a_65865_69663# a_66389_69443# 0.04522f
C4455 a_65589_69723# a_66254_69344# 0.19065f
C4456 VSSD a_60945_61941# 0.28764f
C4457 m3_33828_97932# c1_32748_97972# 0.15596f
C4458 VSSR m3_n1472_23818# 0.66371f
C4459 a_60969_51311# a_61358_51694# 0.06034f
C4460 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A VDDR 0.38472f
C4461 a_61395_49960# a_61609_50282# 0.04522f
C4462 sar10b_0.net43 sar10b_0.net44 0.05055f
C4463 c1_38396_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26825f
C4464 c1_45456_39538# VDDR 0.01151f
C4465 sar10b_0.CF[5] VDDD 0.33621f
C4466 m3_45124_42858# th_dif_sw_0.VCN 0.17339f
C4467 VSSD a_61086_65970# 0.27183f
C4468 sar10b_0._08_ CLK 0.20097f
C4469 sar10b_0.CF[6] VSSA 0.11513f
C4470 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 sar10b_0.CF[0] 0.40695f
C4471 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.11339f
C4472 m3_15472_97932# th_dif_sw_0.VCP 0.01078f
C4473 sar10b_0.SWN[1] VSSA 0.24827f
C4474 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y 0.32324f
C4475 sar10b_0.net16 a_61358_57022# 0.20509f
C4476 sar10b_0.net33 a_65957_50273# 0.02852f
C4477 sar10b_0._13_ a_68276_50645# 0.01537f
C4478 sar10b_0._14_ sar10b_0._08_ 0.15399f
C4479 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.05472f
C4480 VSSR m3_n1472_64332# 0.66316f
C4481 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR 0.38366f
C4482 sar10b_0.net4 a_62185_66027# 0.04078f
C4483 c1_45456_45138# c1_45456_44018# 0.13255f
C4484 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y sar10b_0.CF[9] 0.12541f
C4485 a_43467_5788# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 2.98903f
C4486 sar10b_0._06_ a_67055_68689# 0.09554f
C4487 m3_12648_21578# VCM 0.13579f
C4488 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y 0.07183f
C4489 c1_n1140_66612# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C4490 m3_45124_46218# m3_45124_45098# 0.29566f
C4491 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR 0.59284f
C4492 VDDD a_64491_48621# 0.27338f
C4493 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A 0.07418f
C4494 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A VDDR 0.75806f
C4495 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A 0.60103f
C4496 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 5.31293f
C4497 VDDD a_66666_51977# 0.08613f
C4498 VDDD a_62527_58306# 0.20468f
C4499 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 a_25137_5779# 0.4393f
C4500 sar10b_0.net1 a_64831_56974# 0.01355f
C4501 sar10b_0.net16 sar10b_0.net6 1.78172f
C4502 a_61773_52237# a_62281_52347# 0.19065f
C4503 VDDD a_63918_50969# 0.08958f
C4504 VDDR th_dif_sw_0.VCN 0.66161f
C4505 a_60969_57971# a_62181_58100# 0.07766f
C4506 a_61153_58263# a_61493_58256# 0.24088f
C4507 VDDD a_66109_49318# 0.01418f
C4508 c1_n1140_40658# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C4509 a_64780_52239# sar10b_0.net16 0.13564f
C4510 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y sar10b_0.CF[2] 0.12541f
C4511 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP sar10b_0.CF[9] 0.10502f
C4512 sar10b_0.net3 a_67209_66999# 0.18328f
C4513 VSSD a_66049_57307# 0.81881f
C4514 sar10b_0.SWP[5] VDDR 2.22468f
C4515 VSSR c1_n1140_30578# 0.04956f
C4516 a_62025_51015# a_62277_50968# 0.27388f
C4517 m3_45124_73292# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C4518 m3_45124_86732# m3_45124_85612# 0.29566f
C4519 VSSR m3_28180_97932# 0.46562f
C4520 th_dif_sw_0.CKB sar10b_0.SWN[0] 0.13373f
C4521 VDDD a_62133_59067# 0.30196f
C4522 m3_28180_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.30309f
C4523 m3_45124_48458# VDDR 0.0103f
C4524 a_61395_52624# a_61400_52964# 0.43491f
C4525 a_60945_52617# a_61086_52650# 0.27388f
C4526 a_64373_63584# VSSD 0.11846f
C4527 VDDD sar10b_0.net14 4.10525f
C4528 a_60693_51315# sar10b_0.net16 0.22448f
C4529 VDDD a_67209_64335# 0.91f
C4530 a_61493_67580# sar10b_0.net16 0.15781f
C4531 VDDD sar10b_0.net29 0.59403f
C4532 a_6634_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A 0.01076f
C4533 VSSR c1_5920_97972# 0.05923f
C4534 a_66079_59638# sar10b_0.net16 0.04109f
C4535 a_61065_51015# VSSD 0.48932f
C4536 sar10b_0.clknet_0_CLK a_66865_52076# 0.01461f
C4537 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_n1472_21578# 0.03017f
C4538 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 0.24771f
C4539 VDDD DATA[3] 0.36785f
C4540 sar10b_0.net2 a_62222_57356# 0.01316f
C4541 c1_45456_49618# m3_45124_48458# 0.01078f
C4542 c1_45456_95732# c1_45456_94612# 0.13255f
C4543 c1_n1140_48498# m3_n1472_48458# 1.74381f
C4544 c1_45456_48498# m3_45124_49578# 0.01078f
C4545 VDDD a_60747_60609# 0.22622f
C4546 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A 0.01751f
C4547 a_60693_57975# sar10b_0.net4 0.05863f
C4548 sar10b_0.net38 sar10b_0.CF[2] 0.01398f
C4549 sar10b_0.clknet_0_CLK a_66368_49417# 0.01389f
C4550 a_65865_69663# a_66559_68962# 0.0165f
C4551 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VCM 2.64982f
C4552 m3_45124_88972# VDDR 0.01034f
C4553 m3_45124_85612# th_dif_sw_0.VCP 0.17339f
C4554 VDDD a_62261_56123# 0.20552f
C4555 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A 0.45324f
C4556 sar10b_0.net47 sar10b_0.cyclic_flag_0.FINAL 0.40667f
C4557 sar10b_0.net40 a_66633_56639# 0.01977f
C4558 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A sar10b_0.CF[1] 0.26294f
C4559 CLK sar10b_0.CF[2] 0.1796f
C4560 c1_45456_97972# VDDR 0.01153f
C4561 a_66080_53027# a_66378_52993# 0.02614f
C4562 VDDD a_68325_56296# 0.27541f
C4563 sar10b_0.SWN[2] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.23412f
C4564 sar10b_0.net34 a_65577_51311# 0.0635f
C4565 sar10b_0._03_ a_66312_50368# 0.05567f
C4566 c1_25688_97972# VCM 0.01358f
C4567 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR 0.95198f
C4568 sar10b_0.net3 a_67445_61451# 0.16765f
C4569 sar10b_0.net16 a_65857_56931# 0.09855f
C4570 m3_n1472_71052# c1_n1140_69972# 0.01078f
C4571 m3_45124_71052# c1_45456_71092# 1.74381f
C4572 m3_n1472_69932# c1_n1140_71092# 0.01078f
C4573 VSSR a_29061_5788# 0.06033f
C4574 VSSR c1_45456_74452# 0.0935f
C4575 a_14655_111306# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 0.3928f
C4576 m3_7000_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.53769f
C4577 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VSSR 1.33727f
C4578 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 0.20887f
C4579 c1_29924_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C4580 a_67733_68111# VSSD 0.09968f
C4581 sar10b_0.net33 a_65966_58354# 0.0288f
C4582 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.10847f
C4583 m3_23944_97932# m3_25356_97932# 0.23959f
C4584 a_66933_59067# sar10b_0.net3 0.22888f
C4585 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP sar10b_0.CF[3] 0.10517f
C4586 a_60969_67295# a_61493_67580# 0.05022f
C4587 c1_n1140_87892# c1_n1140_86772# 0.13255f
C4588 c1_11568_21618# m3_11236_21578# 1.74381f
C4589 sar10b_0.CF[4] sar10b_0.CF[3] 48.9619f
C4590 sar10b_0.CF[5] sar10b_0.CF[2] 0.106f
C4591 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 17.8827f
C4592 m3_n1472_49578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C4593 sar10b_0._14_ sar10b_0._15_ 0.21891f
C4594 sar10b_0.SWN[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.01417f
C4595 VDDD a_63457_56931# 0.21676f
C4596 a_65733_59432# a_66079_59638# 0.07649f
C4597 th_dif_sw_0.VCP th_dif_sw_0.CK 17.2624f
C4598 sar10b_0.SWP[3] sar10b_0.CF[9] 0.20205f
C4599 a_66645_60399# VSSD 0.1394f
C4600 m3_14060_97932# c1_12980_97972# 0.15596f
C4601 a_61493_51596# CLK 0.01417f
C4602 VSSR m3_n1472_39498# 0.66371f
C4603 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN sar10b_0.SWP[4] 0.22155f
C4604 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP 7.39338f
C4605 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 1.72813f
C4606 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VCM 10.6522f
C4607 sar10b_0.net47 a_67393_67963# 0.04316f
C4608 a_65586_50645# a_66593_50645# 0.08338f
C4609 c1_45456_55218# VDDR 0.01151f
C4610 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A 1.37832f
C4611 VDDD sar10b_0.SWP[9] 0.45048f
C4612 m3_38064_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C4613 VSSR c1_24276_21618# 0.05929f
C4614 sar10b_0.net4 a_60747_56239# 0.03584f
C4615 a_64949_64916# sar10b_0.net16 0.1551f
C4616 a_67393_54643# a_67733_54791# 0.24088f
C4617 a_67209_55011# a_68421_54964# 0.07766f
C4618 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 0.21251f
C4619 a_19457_5788# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 0.4985f
C4620 VSSR m3_n1472_80012# 0.66316f
C4621 VDDD a_67843_52961# 0.01015f
C4622 c1_45456_52978# c1_45456_51858# 0.13255f
C4623 a_67881_60339# a_68133_60292# 0.27388f
C4624 sar10b_0.net3 a_67598_54692# 0.25847f
C4625 sar10b_0.net38 a_66633_56639# 0.06774f
C4626 VDDA th_dif_sw_0.th_sw_1.CK 2.05852f
C4627 th_dif_sw_0.VCN a_51345_60437# 0.11478f
C4628 sar10b_0.net40 a_61677_64842# 0.01034f
C4629 a_61737_56343# a_61921_55975# 0.43491f
C4630 m3_n1472_23818# VDDR 0.02681f
C4631 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 0.02632f
C4632 sar10b_0.net30 sar10b_0.net16 0.03689f
C4633 VSSD a_61929_56639# 0.27663f
C4634 m3_n1472_31658# VCM 0.01415f
C4635 c1_n1140_82292# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C4636 m3_45124_54058# m3_45124_52938# 0.29566f
C4637 sar10b_0.SWP[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A 0.01082f
C4638 sar10b_0.clknet_1_0__leaf_CLK a_65068_49569# 0.01539f
C4639 sar10b_0.CF[3] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.0136f
C4640 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 3.00838f
C4641 sar10b_0.net16 a_61400_64952# 0.12472f
C4642 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_42300_21578# 0.0162f
C4643 sar10b_0.CF[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A 0.03041f
C4644 sar10b_0.net33 a_66080_53027# 0.01995f
C4645 c1_44044_21618# VCM 0.01358f
C4646 VDDD sar10b_0.net10 1.51432f
C4647 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y 0.31983f
C4648 a_67297_55975# a_68073_56343# 0.3578f
C4649 sar10b_0.net1 sar10b_0.net5 0.30965f
C4650 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A 0.26364f
C4651 m3_n1472_64332# VDDR 0.02674f
C4652 sar10b_0.CF[6] th_dif_sw_0.VCN 0.28584f
C4653 VDDD sar10b_0.net13 3.42434f
C4654 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A sar10b_0.CF[2] 0.26294f
C4655 sar10b_0.net32 sar10b_0.net17 0.0776f
C4656 sar10b_0.net16 VSSD 20.4398f
C4657 m3_n1472_72172# VCM 0.01412f
C4658 VDDD a_67598_65348# 0.27471f
C4659 a_63745_59971# a_64773_60292# 0.07826f
C4660 a_65673_56639# a_66197_56924# 0.05022f
C4661 VSSR sar10b_0.SWP[6] 4.17357f
C4662 th_dif_sw_0.th_sw_1.CKB th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 0.35456f
C4663 c1_n1140_56338# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C4664 sar10b_0.SWN[4] sar10b_0.CF[7] 0.12407f
C4665 sar10b_0.net16 a_63561_60339# 0.2664f
C4666 sar10b_0.CF[6] sar10b_0.SWP[5] 0.1186f
C4667 th_dif_sw_0.CKB a_61419_48621# 0.14263f
C4668 VSSD a_67310_61352# 0.13042f
C4669 VDDD a_65198_66346# 0.2676f
C4670 a_65185_68919# a_65961_68627# 0.3578f
C4671 VSSR c1_n1140_46258# 0.04956f
C4672 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A 0.03718f
C4673 sar10b_0.net28 a_62025_51015# 0.02238f
C4674 sar10b_0.net16 a_61400_60956# 0.10092f
C4675 a_67209_59007# VSSD 0.55806f
C4676 m3_45124_88972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C4677 a_33863_107882# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.81562f
C4678 a_66464_50363# a_66312_50368# 0.22517f
C4679 a_65957_50273# a_66961_50219# 0.06302f
C4680 VDDD a_67564_50907# 0.2329f
C4681 m3_45124_94572# m3_45124_93452# 0.29566f
C4682 VDDD a_68946_52411# 0.27099f
C4683 VDDD sar10b_0.net46 1.27375f
C4684 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN 1.63976f
C4685 m3_35240_21578# c1_35572_21618# 1.74381f
C4686 m3_45124_26058# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C4687 sar10b_0.CF[0] sar10b_0.CF[7] 0.11657f
C4688 sar10b_0.cyclic_flag_0.FINAL sar10b_0.net43 0.04781f
C4689 sar10b_0.net3 a_67798_52206# 0.02392f
C4690 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSSR 4.82113f
C4691 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.32324f
C4692 a_64521_59303# sar10b_0.net11 0.21361f
C4693 a_62997_56643# a_63273_56639# 0.1263f
C4694 m3_43712_97932# c1_44044_97972# 1.74381f
C4695 sar10b_0.net34 a_66101_58256# 0.01136f
C4696 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VCM 1.46158f
C4697 VSSR m3_14060_21578# 0.49683f
C4698 sar10b_0.net6 a_62697_56343# 0.05181f
C4699 tdc_0.RDY sar10b_0.net4 0.27726f
C4700 VSSD sar10b_0.CF[3] 0.81437f
C4701 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.24774f
C4702 a_61400_63620# sar10b_0.net4 0.01892f
C4703 a_60969_67295# VSSD 0.51558f
C4704 sar10b_0.SWN[7] VSSA 0.24841f
C4705 sar10b_0.net32 sar10b_0.net12 0.16929f
C4706 sar10b_0.net3 a_66666_49313# 0.05009f
C4707 sar10b_0.net33 a_66109_51982# 0.01341f
C4708 a_65733_59432# VSSD 0.27321f
C4709 c1_n1140_56338# m3_n1472_56298# 1.74381f
C4710 c1_45456_57458# m3_45124_56298# 0.01078f
C4711 tdc_0.RDY tdc_0.phase_detector_0.pd_out_0.B 0.0472f
C4712 sar10b_0.net14 a_62527_67630# 0.28647f
C4713 m3_8412_97932# VCM 0.15231f
C4714 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A 0.68875f
C4715 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A 0.26294f
C4716 sar10b_0.net16 sar10b_0.net31 0.1871f
C4717 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_29924_21618# 0.0106f
C4718 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 0.39671f
C4719 sar10b_0.SWN[4] sar10b_0.SWN[5] 14.3558f
C4720 sar10b_0.SWP[5] a_19457_110450# 0.5431f
C4721 VDDD a_63525_61624# 0.27236f
C4722 a_67393_54643# VSSD 0.85357f
C4723 sar10b_0.net4 a_61358_67678# 0.06841f
C4724 sar10b_0.net2 sar10b_0.net1 1.71563f
C4725 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 0.21212f
C4726 a_61395_61948# a_61677_62178# 0.05462f
C4727 VDDD a_62997_67299# 0.29209f
C4728 a_60945_61941# a_61609_62270# 0.16939f
C4729 sar10b_0.net39 a_63273_56639# 0.02396f
C4730 a_60747_68227# VSSD 0.32809f
C4731 m3_12648_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C4732 m3_33828_21578# VCM 0.15071f
C4733 m3_45124_78892# c1_45456_78932# 1.74381f
C4734 m3_n1472_78892# c1_n1140_77812# 0.01078f
C4735 m3_n1472_77772# c1_n1140_78932# 0.01078f
C4736 VSSR c1_45456_90132# 0.0935f
C4737 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.41774f
C4738 a_67598_64016# sar10b_0.net3 0.25664f
C4739 sar10b_0.SWN[6] VSSA 0.24837f
C4740 sar10b_0.cyclic_flag_0.FINAL a_64888_67630# 0.11798f
C4741 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A 0.10815f
C4742 a_64085_60119# VSSD 0.14672f
C4743 m3_4176_97932# m3_5588_97932# 0.23959f
C4744 a_64425_64631# a_65637_64760# 0.07766f
C4745 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VSSR 22.8984f
C4746 c1_45456_24978# m3_45124_24938# 1.74381f
C4747 c1_n1140_24978# m3_n1472_23818# 0.01078f
C4748 c1_n1140_23858# m3_n1472_24938# 0.01078f
C4749 VSSR CLK 12.9516f
C4750 sar10b_0.net40 a_63391_57320# 0.30426f
C4751 a_61400_66284# a_61609_66266# 0.24088f
C4752 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[4] 0.05939f
C4753 a_67696_52265# sar10b_0.clk_div_0.COUNT\[2\] 0.23978f
C4754 a_67055_68689# sar10b_0.net45 0.02418f
C4755 a_63950_60020# a_63285_60399# 0.19065f
C4756 a_64085_60119# a_63561_60339# 0.04522f
C4757 VDDD a_65586_50645# 0.45483f
C4758 a_61041_52340# sar10b_0.net16 0.28706f
C4759 sar10b_0.clk_div_0.COUNT\[1\] sar10b_0.clk_div_0.COUNT\[2\] 0.26026f
C4760 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A 0.11547f
C4761 VDDD a_63509_62783# 0.20261f
C4762 sar10b_0._17_ VSSD 0.39479f
C4763 VSSR m3_n1472_55178# 0.66371f
C4764 VDDD a_64428_50947# 0.14215f
C4765 VDDR a_29061_5788# 5.61521f
C4766 c1_45456_74452# VDDR 0.01153f
C4767 sar10b_0.CF[3] sar10b_0.CF[8] 0.10869f
C4768 m3_n1472_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C4769 sar10b_0.net42 a_64238_67295# 0.02167f
C4770 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y 0.32408f
C4771 m3_29592_21578# m3_31004_21578# 0.23959f
C4772 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VDDR 0.74952f
C4773 sar10b_0.CF[5] VSSR 21.8281f
C4774 VSSR c1_45456_22738# 0.09348f
C4775 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.95198f
C4776 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A 0.41861f
C4777 a_14655_5788# VSSR 0.06033f
C4778 sar10b_0.net4 a_62497_61303# 0.01947f
C4779 sar10b_0.net27 a_68946_68627# 0.26211f
C4780 m3_n1472_64332# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C4781 a_61249_53311# sar10b_0.net1 0.02325f
C4782 a_65861_49313# sar10b_0.SWN[6] 0.06243f
C4783 a_65301_57975# a_65761_58263# 0.26257f
C4784 VSSR m3_n1472_95692# 0.66316f
C4785 c1_45456_64372# c1_45456_63252# 0.13255f
C4786 sar10b_0._09_ a_64924_52385# 0.1415f
C4787 a_61677_63510# sar10b_0.net39 0.0216f
C4788 a_67696_52265# VSSD 0.20527f
C4789 m3_n1472_39498# VDDR 0.02681f
C4790 m3_n1472_47338# VCM 0.01415f
C4791 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A 0.41861f
C4792 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 0.19508f
C4793 sar10b_0.clk_div_0.COUNT\[1\] VSSD 1.95435f
C4794 VSSA sar10b_0.CF[7] 0.11513f
C4795 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.02638f
C4796 a_60747_68227# sar10b_0.CF[8] 0.14211f
C4797 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A 0.83558f
C4798 sar10b_0.cyclic_flag_0.FINAL a_67393_66631# 0.08f
C4799 a_65983_64966# sar10b_0.net14 0.01756f
C4800 a_60945_64605# a_61400_64952# 0.3578f
C4801 VSSR c1_27100_97972# 0.06179f
C4802 sar10b_0.net33 sar10b_0._10_ 0.06066f
C4803 a_66789_58100# a_67135_58306# 0.07649f
C4804 sar10b_0.net8 a_62793_57675# 0.0293f
C4805 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A sar10b_0.CF[7] 0.03041f
C4806 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_19708_21578# 0.03017f
C4807 a_65577_57971# sar10b_0.net14 0.02053f
C4808 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_2764_21578# 0.0162f
C4809 sar10b_0.clknet_0_CLK a_65765_50645# 0.01168f
C4810 c1_17216_21618# VCM 0.01358f
C4811 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP a_29061_108738# 0.16709f
C4812 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN sar10b_0.CF[2] 0.12381f
C4813 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45324f
C4814 VSSD a_60945_64605# 0.28758f
C4815 a_61609_63602# a_61677_63510# 0.35559f
C4816 a_61400_63620# a_62185_63363# 0.26257f
C4817 m3_n1472_80012# VDDR 0.02674f
C4818 sar10b_0.net12 a_65589_57735# 0.05234f
C4819 VSSD a_66789_58100# 0.26904f
C4820 VDDD a_61395_61948# 0.85895f
C4821 m3_n1472_87852# VCM 0.01412f
C4822 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.41774f
C4823 c1_n1140_28338# c1_n1140_27218# 0.13255f
C4824 VSSR cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 58.0445f
C4825 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A 0.11547f
C4826 a_61249_50647# sar10b_0.net1 0.02399f
C4827 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR 0.4143f
C4828 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A 0.39707f
C4829 sar10b_0.SWP[4] sar10b_0.CF[4] 2.39963f
C4830 VDDD a_60945_65937# 0.40355f
C4831 a_62798_58688# VSSD 0.12948f
C4832 VCM sar10b_0.SWP[2] 0.13074f
C4833 a_24259_109594# VSSR 0.06033f
C4834 a_65778_49979# a_65957_50273# 0.54361f
C4835 a_67209_65667# a_66933_65727# 0.1263f
C4836 a_n4470_53722# th_dif_sw_0.th_sw_1.CKB 2.27999f
C4837 m3_n1472_29418# m3_n1472_28298# 0.29566f
C4838 a_64780_52239# sar10b_0._07_ 0.02606f
C4839 VSSR c1_n1140_65492# 0.04956f
C4840 a_67393_63967# VSSD 0.85606f
C4841 sar10b_0.net4 a_61705_51992# 0.0342f
C4842 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 1.37832f
C4843 sar10b_0.net33 sar10b_0.net39 0.02767f
C4844 m3_28180_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.30309f
C4845 sar10b_0.net21 sar10b_0.net36 0.02682f
C4846 a_62527_51646# sar10b_0.net28 0.29855f
C4847 a_67209_64335# a_68169_64335# 0.03471f
C4848 a_67393_63967# a_67733_64115# 0.24088f
C4849 sar10b_0.net7 sar10b_0.net1 0.1961f
C4850 sar10b_0._07_ sar10b_0._02_ 0.1287f
C4851 VDDD a_61677_52854# 0.27046f
C4852 m3_45124_41738# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C4853 sar10b_0.SWN[5] VSSA 0.24829f
C4854 a_60693_56643# a_61358_57022# 0.19065f
C4855 sar10b_0.net14 a_65865_69663# 0.22895f
C4856 VSSD a_60945_60609# 0.26438f
C4857 VDDR sar10b_0.SWP[6] 1.88228f
C4858 c1_5920_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26825f
C4859 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP sar10b_0.CF[8] 0.20882f
C4860 a_64809_65963# a_65198_66346# 0.06034f
C4861 m3_23944_97932# c1_24276_97972# 1.74381f
C4862 VSSD a_62697_56343# 0.29061f
C4863 a_64993_66255# a_65769_65963# 0.3578f
C4864 sar10b_0.net16 a_64492_67433# 0.16808f
C4865 VSSR m3_45124_31658# 0.63261f
C4866 a_66153_48647# sar10b_0.net35 0.04929f
C4867 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A a_30644_111636# 0.01076f
C4868 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] th_dif_sw_0.VCP 2.24218f
C4869 sar10b_0.net3 a_68169_65667# 0.27548f
C4870 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A 0.45324f
C4871 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A 0.03718f
C4872 VSSR c1_45456_21618# 0.11545f
C4873 a_60945_60609# a_61400_60956# 0.3578f
C4874 a_61395_60616# a_61609_60938# 0.04522f
C4875 a_65390_69010# VSSD 0.1245f
C4876 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C4877 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_3096_21618# 0.0106f
C4878 m3_n1472_69932# m3_n1472_68812# 0.29566f
C4879 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR 2.59302f
C4880 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.31983f
C4881 VSSR m3_45124_72172# 0.63305f
C4882 VCM cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 2.58383f
C4883 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A 0.43773f
C4884 a_64543_62648# sar10b_0.net16 0.04218f
C4885 a_62697_56343# a_63295_55988# 0.06623f
C4886 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C4887 VSSD a_64233_56639# 0.30737f
C4888 sar10b_0.SWP[7] sar10b_0.SWP[6] 17.8531f
C4889 m3_n1472_85612# c1_n1140_86772# 0.01078f
C4890 m3_n1472_86732# c1_n1140_85652# 0.01078f
C4891 m3_45124_86732# c1_45456_86772# 1.74381f
C4892 a_64199_50761# a_64761_51028# 0.05308f
C4893 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 sar10b_0.CF[9] 0.40665f
C4894 sar10b_0.cyclic_flag_0.FINAL a_67077_57628# 0.01476f
C4895 sar10b_0.net4 a_61395_52624# 0.20995f
C4896 c1_n1140_32818# m3_n1472_31658# 0.01078f
C4897 VSSA th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 2.12205f
C4898 c1_45456_32818# m3_45124_32778# 1.74381f
C4899 c1_n1140_31698# m3_n1472_32778# 0.01078f
C4900 VDDD a_64033_63591# 0.21793f
C4901 sar10b_0.SWN[4] a_25137_5779# 0.48461f
C4902 a_67733_66779# a_68169_66999# 0.16939f
C4903 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] a_39543_5779# 1.0337f
C4904 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C4905 a_65061_63428# a_65407_63634# 0.07649f
C4906 a_64373_63584# a_64238_63682# 0.35559f
C4907 a_65577_57971# sar10b_0.net13 0.20816f
C4908 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A 1.3479f
C4909 sar10b_0.SWP[0] sar10b_0.SWP[1] 7.30218f
C4910 a_68946_63299# sar10b_0.net25 0.26112f
C4911 a_67552_52656# VSSD 0.01142f
C4912 c1_45456_90132# VDDR 0.01153f
C4913 sar10b_0.net18 a_69003_48621# 0.06223f
C4914 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38377f
C4915 sar10b_0.CF[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05939f
C4916 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 1.05065f
C4917 sar10b_0._16_ sar10b_0.clk_div_0.COUNT\[3\] 0.13158f
C4918 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A sar10b_0.CF[0] 0.02149f
C4919 m3_9824_21578# m3_11236_21578# 0.23959f
C4920 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 11.9058f
C4921 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 18.0458f
C4922 sar10b_0.SWN[4] EN 0.17358f
C4923 VSSD a_62357_57455# 0.08338f
C4924 sar10b_0.net40 a_62185_62031# 0.01351f
C4925 VSSR c1_45456_38418# 0.09348f
C4926 a_60789_51075# a_61249_50647# 0.26257f
C4927 a_61065_51015# a_61454_50696# 0.05462f
C4928 sar10b_0.SWN[0] sar10b_0.CF[3] 0.12398f
C4929 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 4.02253f
C4930 VSSR sar10b_0.SWP[9] 3.2416f
C4931 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VDDR 5.22497f
C4932 VDDR CLK 0.25718f
C4933 sar10b_0.net34 a_66255_50749# 0.01475f
C4934 sar10b_0.net23 a_68479_61316# 0.01327f
C4935 VDDD a_61358_51694# 0.28819f
C4936 a_65682_51977# VSSD 1.14103f
C4937 sar10b_0.net19 VSSD 1.10032f
C4938 sar10b_0.net16 a_61400_50300# 0.09895f
C4939 sar10b_0.SWP[4] VSSD 1.00172f
C4940 m3_n1472_80012# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C4941 VDDD a_68946_59303# 0.27936f
C4942 sar10b_0.net4 a_61773_52237# 0.05765f
C4943 sar10b_0.net40 sar10b_0.net12 0.24431f
C4944 VSSR m3_9824_97932# 0.4731f
C4945 c1_45456_72212# c1_45456_71092# 0.13255f
C4946 sar10b_0.clk_div_0.COUNT\[2\] sar10b_0._07_ 0.28839f
C4947 sar10b_0.net16 a_61609_62270# 0.15837f
C4948 m3_9824_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 1.01327f
C4949 VDDD sar10b_0.net42 1.93252f
C4950 sar10b_0.SWP[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A 0.02059f
C4951 m3_n1472_55178# VDDR 0.02681f
C4952 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 3.10203f
C4953 a_64233_56639# sar10b_0.net31 0.05404f
C4954 a_62497_61303# a_63273_61671# 0.3578f
C4955 sar10b_0.net7 a_60789_51075# 0.04023f
C4956 sar10b_0.net16 a_61677_66174# 0.22665f
C4957 VSSR m3_35240_21578# 0.54637f
C4958 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y 0.31995f
C4959 a_66027_53575# sar10b_0._05_ 0.14263f
C4960 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 4.61508f
C4961 VDDD a_67598_68012# 0.27516f
C4962 c1_45456_22738# VDDR 0.01151f
C4963 sar10b_0.CF[5] VDDR 1.73433f
C4964 m3_45124_26058# th_dif_sw_0.VCN 0.17339f
C4965 a_14655_5788# VDDR 3.22284f
C4966 sar10b_0.net14 a_65001_68627# 0.029f
C4967 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN sar10b_0.CF[3] 0.12378f
C4968 m3_n1472_95692# VDDR 0.02674f
C4969 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP 3.44425f
C4970 VDDD a_66921_60339# 0.89947f
C4971 a_67077_69616# sar10b_0.net45 0.01801f
C4972 m3_29592_97932# VCM 0.13579f
C4973 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A 1.37832f
C4974 sar10b_0.net19 sar10b_0.net20 1.56015f
C4975 sar10b_0.SWP[0] th_dif_sw_0.CK 0.093f
C4976 c1_n1140_36178# c1_n1140_35058# 0.13255f
C4977 sar10b_0._07_ VSSD 1.40814f
C4978 VSSD DATA[5] 0.80661f
C4979 a_66933_64395# sar10b_0.net43 0.17078f
C4980 a_60969_51311# sar10b_0.net1 0.07502f
C4981 c1_7332_97972# VCM 0.01358f
C4982 m3_33828_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C4983 th_dif_sw_0.VCN sar10b_0.CF[7] 0.28585f
C4984 m3_n1472_37258# m3_n1472_36138# 0.29566f
C4985 VSSR c1_n1140_81172# 0.04956f
C4986 VDDD a_67084_53565# 0.41343f
C4987 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 7.22725f
C4988 sar10b_0.SWP[3] sar10b_0.SWP[2] 10.8273f
C4989 m3_19708_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.09361f
C4990 sar10b_0.cyclic_flag_0.FINAL a_67297_55975# 0.08105f
C4991 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] c1_22864_21618# 0.02527f
C4992 sar10b_0.net46 a_65865_69663# 0.01487f
C4993 c1_11568_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C4994 sar10b_0.CF[6] sar10b_0.SWP[6] 2.43565f
C4995 sar10b_0.SWP[4] sar10b_0.CF[8] 0.125f
C4996 sar10b_0.SWP[5] sar10b_0.CF[7] 0.12317f
C4997 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 0.56487f
C4998 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C4999 a_61454_53360# sar10b_0.net16 0.22853f
C5000 c1_1684_21618# m3_2764_21578# 0.15596f
C5001 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 0.26289f
C5002 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38377f
C5003 VDDD a_62181_56768# 0.25683f
C5004 sar10b_0.net38 sar10b_0.net12 0.02547f
C5005 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 0.12068f
C5006 VDDR cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 11.373f
C5007 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR 0.38781f
C5008 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A VDDR 0.60057f
C5009 VDDD a_67733_62783# 0.20874f
C5010 m3_4176_97932# c1_4508_97972# 1.74381f
C5011 a_24259_109594# VDDR 4.81771f
C5012 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.36333f
C5013 VSSR m3_45124_47338# 0.63261f
C5014 a_n8277_54249# EN 0.04264f
C5015 c1_n1140_23858# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C5016 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] sar10b_0.SWN[8] 0.22497f
C5017 c1_n1140_62132# th_dif_sw_0.VCP 0.02482f
C5018 m3_19708_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C5019 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 0.20739f
C5020 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 0.12357f
C5021 VSSD a_63457_67583# 0.91807f
C5022 a_62985_63003# a_63169_62635# 0.43491f
C5023 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.83558f
C5024 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN sar10b_0.CF[1] 0.10492f
C5025 VSSR a_10731_113461# 1.11603f
C5026 VSSR c1_18628_21618# 0.05435f
C5027 sar10b_0.SWN[3] a_29939_5779# 0.56255f
C5028 VDDD a_61419_71265# 0.2904f
C5029 a_n4470_53722# a_n8277_54249# 0.01417f
C5030 a_62017_57307# a_63045_57628# 0.07826f
C5031 VDDD CKO 0.24297f
C5032 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.01239f
C5033 a_64238_63682# sar10b_0.net16 0.27002f
C5034 m3_n1472_77772# m3_n1472_76652# 0.29566f
C5035 VSSR m3_45124_87852# 0.63305f
C5036 sar10b_0.net3 sar10b_0.clk_div_0.COUNT\[3\] 0.27605f
C5037 a_66645_60399# a_67310_60020# 0.19065f
C5038 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 0.24775f
C5039 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C5040 a_66921_60339# a_67445_60119# 0.04522f
C5041 VSSD a_60693_56643# 0.15023f
C5042 sar10b_0.net38 a_63662_57022# 0.04683f
C5043 m3_45124_31658# VDDR 0.0103f
C5044 VDDD a_67105_61303# 0.28269f
C5045 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05939f
C5046 a_61454_50696# sar10b_0.net16 0.24977f
C5047 sar10b_0.net2 sar10b_0.SWP[0] 0.10795f
C5048 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN sar10b_0.CF[4] 0.12375f
C5049 m3_n1472_94572# c1_n1140_93492# 0.01078f
C5050 a_66103_50668# VSSD 0.11822f
C5051 VSSR c1_45456_96852# 0.0935f
C5052 a_63945_63003# VSSD 0.33388f
C5053 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A 0.68875f
C5054 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.10815f
C5055 VSSA EN 3.74536f
C5056 c1_45456_21618# VDDR 0.01151f
C5057 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[7] 0.05939f
C5058 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_23944_21578# 0.0162f
C5059 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_40888_21578# 0.03017f
C5060 CLK a_51345_60437# 0.32634f
C5061 VDDD a_65577_51311# 1.47042f
C5062 w_n9655_56533# a_n4470_53722# 0.01216f
C5063 c1_25688_21618# VCM 0.01358f
C5064 c1_n1140_39538# m3_n1472_40618# 0.01078f
C5065 c1_n1140_40658# m3_n1472_39498# 0.01078f
C5066 c1_45456_40658# m3_45124_40618# 1.74381f
C5067 a_n4470_65264# th_dif_sw_0.th_sw_1.CK 2.27995f
C5068 m3_45124_68812# th_dif_sw_0.VCP 0.17339f
C5069 m3_45124_72172# VDDR 0.01034f
C5070 sar10b_0.net34 a_66254_57356# 0.01981f
C5071 VDDD sar10b_0.net8 1.62633f
C5072 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A 0.38472f
C5073 m3_28180_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.96307f
C5074 a_n4470_53722# VSSA 2.16753f
C5075 a_61153_56931# a_61737_56343# 0.01027f
C5076 sar10b_0.net9 a_61677_62178# 0.01357f
C5077 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A 0.11547f
C5078 sar10b_0.net7 a_60747_57571# 0.08377f
C5079 sar10b_0.clknet_0_CLK sar10b_0.net16 0.02264f
C5080 VDDD a_67543_51991# 0.01122f
C5081 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A sar10b_0.CF[4] 0.06369f
C5082 sar10b_0.net13 a_65001_68627# 0.23862f
C5083 a_64725_68631# a_65185_68919# 0.26257f
C5084 VDDD a_65045_59588# 0.20068f
C5085 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.21001f
C5086 sar10b_0.CF[6] CLK 0.09331f
C5087 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.01212f
C5088 m3_45124_63212# c1_45456_62132# 0.01078f
C5089 m3_45124_62092# c1_45456_63252# 0.01078f
C5090 m3_n1472_62092# c1_n1140_62132# 1.74381f
C5091 VSSR c1_45456_54098# 0.09348f
C5092 a_60969_57971# sar10b_0.net38 0.01007f
C5093 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR 1.10847f
C5094 sar10b_0._08_ a_65577_51311# 0.9102f
C5095 a_67423_69308# VSSD 0.26883f
C5096 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 0.64443f
C5097 m3_n1472_95692# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C5098 sar10b_0.clk_div_0.COUNT\[3\] a_67798_52206# 0.18032f
C5099 m3_25356_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.19539f
C5100 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] sar10b_0.CF[2] 0.01366f
C5101 c1_45456_80052# c1_45456_78932# 0.13255f
C5102 m3_26768_21578# c1_25688_21618# 0.15596f
C5103 VSSA tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A 0.5729f
C5104 a_62277_53632# a_62623_53324# 0.07649f
C5105 m3_n1472_32778# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C5106 a_60945_49953# VSSD 0.28719f
C5107 a_68767_58652# sar10b_0.net22 0.01983f
C5108 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A 0.75026f
C5109 a_66049_69295# a_66254_69344# 0.09983f
C5110 m3_35240_97932# c1_34160_97972# 0.15596f
C5111 sar10b_0.CF[6] sar10b_0.CF[5] 56.9039f
C5112 VSSD a_61400_62288# 0.85195f
C5113 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C5114 VSSR m3_n1472_22698# 0.66371f
C5115 a_61493_51596# a_61358_51694# 0.35559f
C5116 sar10b_0.CF[5] sar10b_0.SWN[1] 0.1227f
C5117 sar10b_0.net47 a_66825_69663# 0.0161f
C5118 sar10b_0.net1 a_63285_60399# 0.16673f
C5119 VDDD a_63950_60020# 0.2669f
C5120 VDDD a_65673_56639# 0.74653f
C5121 c1_45456_38418# VDDR 0.01151f
C5122 c1_41220_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26825f
C5123 a_25842_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A 0.01076f
C5124 m3_45124_41738# th_dif_sw_0.VCN 0.17339f
C5125 sar10b_0.SWP[9] VDDR 11.358f
C5126 VSSR a_249_113874# 0.06021f
C5127 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_31680_111642# 0.01076f
C5128 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 0.12068f
C5129 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.11339f
C5130 m3_18296_97932# th_dif_sw_0.VCP 0.01078f
C5131 a_60747_49953# EN 0.01181f
C5132 sar10b_0.cyclic_flag_0.FINAL a_67231_56974# 0.01687f
C5133 VDDD a_66027_53575# 0.29241f
C5134 sar10b_0.net14 sar10b_0.net12 0.03352f
C5135 sar10b_0.CF[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.26269f
C5136 a_11436_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A 0.01076f
C5137 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 2.64269f
C5138 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 0.41934f
C5139 c1_20040_21618# th_dif_sw_0.VCN 0.13255f
C5140 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_17274_8700# 0.01076f
C5141 VSSR m3_n1472_63212# 0.66316f
C5142 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 1.76305f
C5143 sar10b_0._10_ sar10b_0._01_ 0.02822f
C5144 c1_n1140_44018# c1_n1140_42898# 0.13255f
C5145 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C5146 w_n9655_63119# a_n8277_66083# 68.4698f
C5147 a_65394_52643# VSSD 1.16778f
C5148 m3_15472_21578# VCM 0.13579f
C5149 sar10b_0.net6 a_61358_57022# 0.01896f
C5150 c1_n1140_65492# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C5151 m3_n1472_45098# m3_n1472_43978# 0.29566f
C5152 VSSR a_20335_5779# 1.79211f
C5153 c1_20040_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 0.01078f
C5154 a_68562_71291# a_69003_71265# 0.02339f
C5155 sar10b_0.net4 a_60690_54641# 0.02772f
C5156 sar10b_0.net45 a_67209_66999# 0.01557f
C5157 VDDD a_64425_64631# 0.83186f
C5158 sar10b_0.net3 a_68169_68331# 0.26947f
C5159 m3_22532_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 0.53272f
C5160 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VDDR 0.83558f
C5161 VDDD a_67372_52243# 0.10437f
C5162 VDDD sar10b_0.net9 1.40771f
C5163 a_67105_59971# sar10b_0.net3 0.11549f
C5164 a_66368_52081# a_66216_52022# 0.22338f
C5165 a_60693_57975# a_61358_58354# 0.19065f
C5166 a_61153_58263# a_61929_57971# 0.3578f
C5167 VDDD a_66216_49358# 0.14476f
C5168 c1_n1140_39538# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C5169 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 4.30791f
C5170 sar10b_0.clknet_0_CLK sar10b_0._17_ 0.04451f
C5171 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 0.02632f
C5172 VDDD a_61395_64612# 0.86128f
C5173 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04073f
C5174 m3_45124_22698# m3_45124_21578# 0.29566f
C5175 a_67105_61303# a_68133_61624# 0.07826f
C5176 sar10b_0.net3 a_66837_56403# 0.2177f
C5177 VSSD a_66389_57455# 0.08231f
C5178 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04073f
C5179 VSSR c1_n1140_29458# 0.04956f
C5180 a_62277_50968# a_62623_50660# 0.07649f
C5181 sar10b_0.net4 a_62025_53679# 0.01006f
C5182 VDDD a_66101_58256# 0.20668f
C5183 sar10b_0.net40 a_62313_61671# 0.02019f
C5184 a_60945_63273# sar10b_0.net16 0.29436f
C5185 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.02638f
C5186 m3_45124_72172# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C5187 a_65682_49313# a_65861_49313# 0.54426f
C5188 m3_n1472_85612# m3_n1472_84492# 0.29566f
C5189 VSSR m3_31004_97932# 0.49843f
C5190 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 2.31287f
C5191 VDDD a_62593_58639# 0.22532f
C5192 m3_31004_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.31585f
C5193 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.59846f
C5194 m3_45124_47338# VDDR 0.0103f
C5195 sar10b_0.net29 sar10b_0.SWN[1] 0.07191f
C5196 a_61395_52624# a_61609_52946# 0.04522f
C5197 a_61086_52650# a_61400_52964# 0.07826f
C5198 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 sar10b_0.CF[3] 0.26311f
C5199 a_64809_63299# VSSD 0.29969f
C5200 a_67209_59007# a_67393_58639# 0.43491f
C5201 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] 18.0458f
C5202 a_61153_51603# sar10b_0.net16 0.10625f
C5203 a_61929_67295# sar10b_0.net16 0.30101f
C5204 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A 0.05472f
C5205 VSSR c1_8744_97972# 0.054f
C5206 th_dif_sw_0.CK sar10b_0.SWP[1] 0.26807f
C5207 a_68421_62956# sar10b_0.net3 0.17818f
C5208 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP sar10b_0.CF[9] 0.19147f
C5209 sar10b_0.net16 a_64533_65967# 0.2394f
C5210 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A 0.28117f
C5211 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A 0.42509f
C5212 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_1352_21578# 0.03017f
C5213 m3_9824_21578# th_dif_sw_0.VCN 0.01078f
C5214 a_66762_50329# VSSD 0.19633f
C5215 c1_n1140_21618# VCM 0.01358f
C5216 a_63457_56931# a_63662_57022# 0.09983f
C5217 c1_n1140_47378# m3_n1472_48458# 0.01078f
C5218 c1_n1140_48498# m3_n1472_47338# 0.01078f
C5219 c1_45456_48498# m3_45124_48458# 1.74381f
C5220 a_62997_67299# a_63663_67678# 0.19082f
C5221 a_63457_67583# a_64492_67433# 0.08258f
C5222 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VCM 0.12357f
C5223 a_61153_58263# sar10b_0.net4 0.1163f
C5224 a_67637_56123# sar10b_0.net35 0.01005f
C5225 m3_45124_87852# VDDR 0.01034f
C5226 m3_45124_84492# th_dif_sw_0.VCP 0.17339f
C5227 VDDD sar10b_0.net21 1.06415f
C5228 sar10b_0.net29 a_60690_49683# 0.05917f
C5229 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A 0.43651f
C5230 a_66666_51977# sar10b_0.clk_div_0.COUNT\[0\] 0.02432f
C5231 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 3.21929f
C5232 a_60747_58903# VSSD 0.32513f
C5233 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] a_19457_5788# 1.48701f
C5234 c1_45456_96852# VDDR 0.01153f
C5235 sar10b_0.net46 sar10b_0.SWP[7] 0.0263f
C5236 a_66577_52883# a_66378_52993# 0.29821f
C5237 sar10b_0._03_ a_67439_50041# 0.07854f
C5238 c1_28512_97972# VCM 0.01358f
C5239 a_64773_60292# sar10b_0.net16 0.17376f
C5240 sar10b_0.net16 a_66885_56768# 0.17333f
C5241 m3_45124_71052# c1_45456_69972# 0.01078f
C5242 m3_n1472_69932# c1_n1140_69972# 1.74381f
C5243 m3_45124_69932# c1_45456_71092# 0.01078f
C5244 a_60690_53975# VSSD 0.51889f
C5245 VSSR c1_45456_73332# 0.0935f
C5246 sar10b_0.net13 sar10b_0.net12 0.30118f
C5247 VDDD a_67055_68689# 0.40256f
C5248 sar10b_0.SWN[3] VCM 0.13076f
C5249 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C5250 m3_9824_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 1.01327f
C5251 c1_32748_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C5252 sar10b_0.SWP[7] a_10731_113461# 0.24998f
C5253 sar10b_0.CF[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A 0.06369f
C5254 m3_25356_97932# m3_26768_97932# 0.23959f
C5255 a_61153_67587# a_62181_67424# 0.07826f
C5256 sar10b_0.net23 sar10b_0.net22 0.79994f
C5257 a_60969_67295# a_61929_67295# 0.03432f
C5258 c1_45456_87892# c1_45456_86772# 0.13255f
C5259 c1_12980_21618# m3_12648_21578# 1.74381f
C5260 sar10b_0.net14 sar10b_0.net41 0.0561f
C5261 m3_n1472_48458# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C5262 VDDD a_64485_56768# 0.25955f
C5263 a_n9133_63315# th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 1.06244f
C5264 a_n8277_66083# a_n8277_65767# 0.64152f
C5265 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 1.72813f
C5266 a_51345_60437# a_51861_60437# 0.08876f
C5267 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_52417_60961# 0.09051f
C5268 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP 0.16581f
C5269 a_61929_51311# CLK 0.02727f
C5270 m3_15472_97932# c1_14392_97972# 0.15596f
C5271 VSSR m3_n1472_38378# 0.66371f
C5272 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VCM 0.12358f
C5273 a_65765_50645# a_66785_50875# 0.05416f
C5274 a_66255_50749# a_66593_50645# 0.02853f
C5275 c1_45456_54098# VDDR 0.01151f
C5276 sar10b_0.net3 sar10b_0.net45 0.17132f
C5277 m3_40888_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C5278 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR 0.95198f
C5279 a_67113_56343# VSSD 0.55314f
C5280 VSSD a_66933_67059# 0.13832f
C5281 a_63945_63003# a_64543_62648# 0.06623f
C5282 VSSR cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.16481p
C5283 a_61803_48621# sar10b_0.SWN[2] 0.11484f
C5284 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.39384f
C5285 sar10b_0.net34 sar10b_0.net3 0.29623f
C5286 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A VSSR 0.43651f
C5287 VSSR c1_27100_21618# 0.06179f
C5288 a_65385_64631# sar10b_0.net16 0.27105f
C5289 VDDD sar10b_0.SWN[2] 0.14347f
C5290 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[3] 0.17717f
C5291 VSSR m3_n1472_78892# 0.66316f
C5292 a_65301_57975# sar10b_0.net16 0.22597f
C5293 a_68133_60292# a_68479_59984# 0.07649f
C5294 c1_n1140_51858# c1_n1140_50738# 0.13255f
C5295 sar10b_0.net40 a_62185_64695# 0.0151f
C5296 m3_n1472_22698# VDDR 0.02681f
C5297 a_61737_56343# a_62261_56123# 0.04522f
C5298 a_61461_56403# a_62126_56024# 0.19065f
C5299 VSSD a_61358_57022# 0.13499f
C5300 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] 2.32591f
C5301 VDDD a_62222_57356# 0.26569f
C5302 m3_n1472_30538# VCM 0.01415f
C5303 a_64188_51135# a_64761_51028# 0.04602f
C5304 c1_n1140_81172# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C5305 m3_n1472_52938# m3_n1472_51818# 0.29566f
C5306 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 2.75093f
C5307 sar10b_0.clknet_1_0__leaf_CLK a_65861_49313# 0.0164f
C5308 a_249_113874# VDDR 0.82898f
C5309 a_68169_63003# VSSD 0.29067f
C5310 VDDD a_64924_52385# 0.10598f
C5311 sar10b_0.net16 a_61609_64934# 0.15597f
C5312 sar10b_0.net30 sar10b_0.net6 0.10206f
C5313 a_61065_53679# a_62277_53632# 0.07766f
C5314 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_45124_21578# 0.0162f
C5315 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 2.64509f
C5316 sar10b_0._14_ sar10b_0.net37 0.5604f
C5317 VDDA VCM 0.4431f
C5318 tdc_0.OUTP sar10b_0.SWP[0] 0.13371f
C5319 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 0.73278f
C5320 a_67637_56123# a_68073_56343# 0.16939f
C5321 th_dif_sw_0.VCP sar10b_0.CF[1] 0.28581f
C5322 m3_n1472_63212# VDDR 0.02674f
C5323 sar10b_0.clk_div_0.COUNT\[1\] a_68178_51635# 0.08966f
C5324 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A 0.06369f
C5325 a_63369_59007# sar10b_0.net16 0.26189f
C5326 m3_n1472_71052# VCM 0.01412f
C5327 sar10b_0.net2 sar10b_0.net5 0.01075f
C5328 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C5329 sar10b_0.net7 a_60843_52216# 0.29053f
C5330 a_65673_56639# a_66633_56639# 0.03432f
C5331 VSSD sar10b_0.net26 0.36299f
C5332 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] sar10b_0.SWN[7] 0.22605f
C5333 c1_n1140_55218# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C5334 sar10b_0.CF[7] sar10b_0.SWP[6] 0.12119f
C5335 a_62409_59007# sar10b_0.net39 0.07924f
C5336 sar10b_0.net40 a_62185_60699# 0.01269f
C5337 VSSR cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 58.0445f
C5338 VSSD sar10b_0.net6 1.80537f
C5339 c1_27100_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.02009f
C5340 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C5341 a_66213_68756# a_65961_68627# 0.27388f
C5342 VSSR c1_n1140_45138# 0.04956f
C5343 a_64780_52239# VSSD 0.24016f
C5344 sar10b_0.net16 a_61609_60938# 0.15764f
C5345 m3_45124_87852# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C5346 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A 0.05472f
C5347 sar10b_0.net4 sar10b_0.net39 0.04719f
C5348 a_65957_50273# a_66205_50408# 0.05308f
C5349 m3_n1472_93452# m3_n1472_92332# 0.29566f
C5350 sar10b_0.net34 a_66666_49313# 0.06814f
C5351 m3_36652_21578# c1_36984_21618# 1.74381f
C5352 m3_45124_24938# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C5353 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.10847f
C5354 sar10b_0.SWP[3] a_29939_111781# 0.56255f
C5355 a_60747_63273# VSSD 0.2587f
C5356 sar10b_0._02_ VSSD 0.42785f
C5357 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A sar10b_0.CF[9] 0.02149f
C5358 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[8] 0.01887f
C5359 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.4249f
C5360 sar10b_0.net34 a_66537_57971# 0.03617f
C5361 m3_45124_97932# c1_45456_97972# 1.74381f
C5362 DATA[1] sar10b_0.net36 0.10364f
C5363 VSSR m3_16884_21578# 0.43913f
C5364 c1_21452_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 0.28822f
C5365 sar10b_0.net10 sar10b_0.net41 0.05283f
C5366 a_68235_71265# VSSD 0.31083f
C5367 tdc_0.RDY VDDA 0.23192f
C5368 a_60693_51315# VSSD 0.14646f
C5369 sar10b_0.net13 sar10b_0.net41 0.0609f
C5370 a_61493_67580# VSSD 0.09866f
C5371 sar10b_0.net3 a_67371_49579# 0.07153f
C5372 sar10b_0.net33 a_66216_52022# 0.01877f
C5373 c1_n1140_55218# m3_n1472_56298# 0.01078f
C5374 c1_n1140_56338# m3_n1472_55178# 0.01078f
C5375 a_66079_59638# VSSD 0.26399f
C5376 c1_45456_56338# m3_45124_56298# 1.74381f
C5377 sar10b_0.CF[4] VSSD 0.92424f
C5378 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN 0.01212f
C5379 a_60945_49953# a_61400_50300# 0.3578f
C5380 m3_11236_97932# VCM 0.13579f
C5381 sar10b_0.net3 sar10b_0.net36 0.02826f
C5382 sar10b_0.SWP[6] a_14655_111306# 0.43739f
C5383 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 0.40575f
C5384 sar10b_0.net4 a_62037_61731# 0.01366f
C5385 sar10b_0.net33 a_65861_49313# 0.02484f
C5386 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_32748_21618# 0.0106f
C5387 a_67733_54791# VSSD 0.09761f
C5388 sar10b_0.net14 a_64993_66255# 0.02661f
C5389 a_14655_5788# sar10b_0.SWN[6] 0.43739f
C5390 a_61400_62288# a_61609_62270# 0.24088f
C5391 a_61395_61948# a_62185_62031# 0.1263f
C5392 m3_36652_21578# VCM 0.15231f
C5393 m3_15472_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C5394 sar10b_0.net6 sar10b_0.net31 0.40532f
C5395 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP 0.02666f
C5396 sar10b_0.clknet_0_CLK sar10b_0._07_ 0.02934f
C5397 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VCM 0.12068f
C5398 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP 0.10502f
C5399 a_67564_50907# a_67611_50645# 0.19021f
C5400 m3_n1472_77772# c1_n1140_77812# 1.74381f
C5401 m3_45124_78892# c1_45456_77812# 0.01078f
C5402 m3_45124_77772# c1_45456_78932# 0.01078f
C5403 VSSR c1_45456_89012# 0.0935f
C5404 sar10b_0.SWP[8] sar10b_0.CF[9] 0.13258f
C5405 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VCM 1.23381f
C5406 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 0.95011f
C5407 VSSD a_65857_56931# 0.85545f
C5408 m3_5588_97932# m3_7000_97932# 0.23959f
C5409 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR 0.36778f
C5410 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A 1.11457f
C5411 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A 0.38427f
C5412 a_64149_64635# a_64814_65014# 0.19065f
C5413 a_64609_64923# a_65637_64760# 0.07826f
C5414 c1_n1140_23858# m3_n1472_23818# 1.74381f
C5415 sar10b_0.SWN[4] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 0.2309f
C5416 c1_45456_23858# m3_45124_24938# 0.01078f
C5417 c1_45456_24978# m3_45124_23818# 0.01078f
C5418 sar10b_0.clk_div_0.COUNT\[0\] a_67564_50907# 0.39714f
C5419 CLK sar10b_0.CF[7] 0.09336f
C5420 sar10b_0.net21 a_68169_55011# 0.01543f
C5421 sar10b_0.net40 a_61395_65944# 0.01746f
C5422 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y 0.07418f
C5423 a_61491_52222# sar10b_0.net16 0.19672f
C5424 a_15533_5779# VSSR 1.45369f
C5425 VDDD a_66255_50749# 0.12547f
C5426 VINN th_dif_sw_0.th_sw_1.CKB 0.08416f
C5427 VSSR m3_n1472_54058# 0.66371f
C5428 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05939f
C5429 sar10b_0.SWN[2] sar10b_0.CF[2] 2.49492f
C5430 a_67209_68331# a_66933_68391# 0.1263f
C5431 sar10b_0.net16 a_63045_57628# 0.17449f
C5432 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A 0.03718f
C5433 c1_45456_73332# VDDR 0.01153f
C5434 m3_1352_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C5435 a_67209_63003# sar10b_0.cyclic_flag_0.FINAL 0.24116f
C5436 m3_31004_21578# m3_32416_21578# 0.23959f
C5437 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN 8.07467f
C5438 VSSR c1_272_21618# 0.05576f
C5439 th_dif_sw_0.CKB VCM 0.24229f
C5440 sar10b_0.CF[5] sar10b_0.CF[7] 0.11787f
C5441 sar10b_0.CF[4] sar10b_0.CF[8] 0.1137f
C5442 sar10b_0.net19 sar10b_0.SWN[9] 0.10368f
C5443 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 2.76087f
C5444 sar10b_0.SWN[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A 0.01417f
C5445 VINP th_dif_sw_0.th_sw_1.CK 0.32471f
C5446 m3_n1472_63212# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C5447 a_61589_53459# sar10b_0.net1 0.01211f
C5448 a_65577_57971# a_66101_58256# 0.05022f
C5449 sar10b_0.net7 sar10b_0.net5 0.50726f
C5450 VSSR m3_n1472_94572# 0.66316f
C5451 a_68325_56296# sar10b_0.net37 0.03018f
C5452 c1_n1140_63252# c1_n1140_62132# 0.13255f
C5453 a_64949_64916# VSSD 0.10335f
C5454 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 4.92029f
C5455 sar10b_0.clk_div_0.COUNT\[2\] VSSD 0.8465f
C5456 m3_n1472_38378# VDDR 0.02681f
C5457 m3_n1472_46218# VCM 0.01415f
C5458 a_68169_59007# a_68421_58960# 0.27388f
C5459 VSSR c1_29924_97972# 0.05685f
C5460 a_60945_64605# a_61609_64934# 0.16939f
C5461 a_61395_64612# a_61677_64842# 0.05462f
C5462 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.39589f
C5463 VDDR cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 14.4489f
C5464 sar10b_0.net30 VSSD 0.56949f
C5465 VDDD a_67077_69616# 0.32427f
C5466 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A 0.28117f
C5467 sar10b_0.net8 a_63391_57320# 0.01644f
C5468 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A VDDR 0.38427f
C5469 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_5588_21578# 0.0162f
C5470 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_22532_21578# 0.02509f
C5471 a_66865_49412# VSSD 0.32823f
C5472 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 0.02638f
C5473 sar10b_0.net16 sar10b_0.net43 0.68392f
C5474 VDDD sar10b_0.net1 4.38435f
C5475 VSSD a_61400_64952# 0.85606f
C5476 m3_n1472_78892# VDDR 0.02674f
C5477 VSSD a_67135_58306# 0.2692f
C5478 VDDD a_61086_61974# 0.31749f
C5479 VDDA sar10b_0.SWP[3] 0.2491f
C5480 sar10b_0.net9 a_61677_60846# 0.04206f
C5481 m3_n1472_86732# VCM 0.01412f
C5482 a_60747_64231# sar10b_0.net11 0.28154f
C5483 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A 0.68875f
C5484 sar10b_0.net34 a_65861_51977# 0.02989f
C5485 sar10b_0.SWP[2] a_33863_107882# 0.86021f
C5486 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.72402f
C5487 c1_45456_28338# c1_45456_27218# 0.13255f
C5488 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 sar10b_0.CF[9] 0.26243f
C5489 VDDD a_61400_66284# 0.25364f
C5490 a_62593_58639# a_63621_58960# 0.07826f
C5491 sar10b_0.net4 sar10b_0.net11 0.18203f
C5492 a_65778_49979# a_66312_50368# 0.35097f
C5493 a_67209_65667# a_67393_65299# 0.44098f
C5494 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C5495 sar10b_0.CF[5] sar10b_0.SWN[5] 2.41127f
C5496 m3_45124_29418# m3_45124_28298# 0.29566f
C5497 VSSR c1_n1140_64372# 0.04956f
C5498 a_64033_63591# sar10b_0.net12 0.02042f
C5499 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 4.32122f
C5500 a_67733_64115# VSSD 0.10001f
C5501 VSSD a_63561_60339# 0.55993f
C5502 m3_31004_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.31585f
C5503 sar10b_0.net3 sar10b_0._04_ 0.02764f
C5504 sar10b_0.SWP[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.21523f
C5505 sar10b_0._13_ a_67439_50041# 0.09566f
C5506 VDDD a_62185_52707# 0.30454f
C5507 m3_45124_40618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C5508 sar10b_0.SWN[4] sar10b_0.CF[9] 0.18391f
C5509 m3_16884_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.66386f
C5510 VSSD a_61400_60956# 0.81519f
C5511 c1_8744_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.28115f
C5512 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C5513 sar10b_0.net7 sar10b_0.net2 0.05808f
C5514 VDDR cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 11.373f
C5515 VSSD a_63295_55988# 0.27285f
C5516 a_64993_66255# a_65198_66346# 0.09983f
C5517 m3_25356_97932# c1_25688_97972# 1.74381f
C5518 a_66021_66092# a_65769_65963# 0.27388f
C5519 sar10b_0.net16 a_64888_67630# 0.02008f
C5520 VSSR m3_45124_30538# 0.63261f
C5521 sar10b_0._10_ a_64199_50761# 0.02573f
C5522 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 1.16488f
C5523 sar10b_0.net30 sar10b_0.net31 0.05881f
C5524 VDDA w_n9655_63119# 1.49178f
C5525 a_64705_59595# a_64910_59686# 0.09983f
C5526 sar10b_0.net20 VSSD 0.67263f
C5527 a_67209_63003# a_67598_62684# 0.05462f
C5528 a_66933_63063# a_67393_62635# 0.26257f
C5529 sar10b_0.net42 sar10b_0.net12 0.05359f
C5530 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A a_39543_110941# 0.01247f
C5531 a_60945_60609# a_61609_60938# 0.16939f
C5532 sar10b_0.CF[0] sar10b_0.CF[9] 0.11283f
C5533 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.95198f
C5534 a_66049_57307# a_67077_57628# 0.07826f
C5535 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_5920_21618# 0.0106f
C5536 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 2.56839f
C5537 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y 0.32264f
C5538 m3_45124_69932# m3_45124_68812# 0.29566f
C5539 VSSR m3_45124_71052# 0.63305f
C5540 m3_23944_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 0.3358f
C5541 a_66785_50875# sar10b_0.net16 0.40284f
C5542 th_dif_sw_0.VCP sar10b_0.CF[2] 0.28618f
C5543 VSSD sar10b_0.net31 2.45904f
C5544 VSSD sar10b_0.CF[8] 0.67585f
C5545 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A 0.11547f
C5546 VDDD a_66254_57356# 0.26996f
C5547 m3_45124_85612# c1_45456_86772# 0.01078f
C5548 m3_45124_86732# c1_45456_85652# 0.01078f
C5549 m3_n1472_85612# c1_n1140_85652# 1.74381f
C5550 a_62313_61671# a_63525_61624# 0.07766f
C5551 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A 0.02842f
C5552 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VCM 0.13025f
C5553 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VSSR 4.36957f
C5554 a_44345_5779# sar10b_0.SWN[0] 0.79636f
C5555 sar10b_0.net23 sar10b_0.net24 0.49782f
C5556 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C5557 c1_45456_31698# m3_45124_32778# 0.01078f
C5558 c1_45456_32818# m3_45124_31658# 0.01078f
C5559 c1_n1140_31698# m3_n1472_31658# 1.74381f
C5560 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 0.30288f
C5561 sar10b_0._09_ sar10b_0._00_ 0.02835f
C5562 VDDD a_65061_63428# 0.27504f
C5563 sar10b_0.net19 a_68562_49747# 0.04127f
C5564 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A sar10b_0.CF[8] 0.26294f
C5565 sar10b_0.net32 sar10b_0.clknet_1_0__leaf_CLK 0.03079f
C5566 CKO sar10b_0.SWP[7] 0.07334f
C5567 VDDD a_60789_51075# 0.33537f
C5568 sar10b_0.net10 a_62985_63003# 0.07468f
C5569 sar10b_0.net31 a_63295_55988# 0.01533f
C5570 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] a_5051_5788# 0.58622f
C5571 a_61041_52340# VSSD 0.28622f
C5572 a_60969_51311# sar10b_0.net5 0.21438f
C5573 c1_45456_89012# VDDR 0.01153f
C5574 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 3.44428f
C5575 a_29939_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A 0.01197f
C5576 m3_11236_21578# m3_12648_21578# 0.23959f
C5577 a_66921_61671# a_66645_61731# 0.1263f
C5578 VSSR c1_45456_37298# 0.09348f
C5579 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A 0.95194f
C5580 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR 0.59327f
C5581 sar10b_0.net16 a_61609_50282# 0.15119f
C5582 m3_n1472_78892# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C5583 tdc_0.OUTP th_dif_sw_0.CK 0.07693f
C5584 VSSR m3_12648_97932# 0.49843f
C5585 sar10b_0.CF[4] sar10b_0.SWN[0] 0.12506f
C5586 c1_n1140_71092# c1_n1140_69972# 0.13255f
C5587 VSSR sar10b_0.SWN[2] 5.56887f
C5588 m3_12648_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.31585f
C5589 a_29939_111781# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A 0.01197f
C5590 m3_n1472_54058# VDDR 0.02681f
C5591 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A 0.07418f
C5592 a_61400_50300# sar10b_0.net6 0.01552f
C5593 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A sar10b_0.CF[9] 0.02149f
C5594 a_62837_61451# a_63273_61671# 0.16939f
C5595 sar10b_0.CF[1] a_60747_57571# 0.14313f
C5596 sar10b_0.SWN[1] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.23544f
C5597 sar10b_0.net7 a_61249_50647# 0.02182f
C5598 sar10b_0.net16 a_62185_66027# 0.22592f
C5599 sar10b_0._08_ a_64818_49979# 0.05079f
C5600 VSSR m3_38064_21578# 0.54637f
C5601 VSSD a_68421_65620# 0.27173f
C5602 a_n8277_54249# VINN 0.64084f
C5603 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VDDR 4.85357f
C5604 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 1.16383f
C5605 m3_45124_24938# th_dif_sw_0.VCN 0.17339f
C5606 a_64033_63591# sar10b_0.net41 0.02009f
C5607 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A 0.02842f
C5608 sar10b_0.net14 a_65525_68912# 0.03657f
C5609 sar10b_0.clknet_0_CLK a_66762_50329# 0.03059f
C5610 m3_n1472_94572# VDDR 0.02674f
C5611 a_1127_114301# sar10b_0.SWP[9] 0.08773f
C5612 m3_32416_97932# VCM 0.13579f
C5613 VSSA sar10b_0.CF[9] 0.12636f
C5614 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] m3_9824_21578# 0.0122f
C5615 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 0.01165f
C5616 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN 3.38193f
C5617 c1_45456_36178# c1_45456_35058# 0.13255f
C5618 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN 0.09308f
C5619 a_66049_69295# sar10b_0.net44 0.02553f
C5620 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP 0.02666f
C5621 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 1.70485f
C5622 VDDD a_67209_66999# 0.8965f
C5623 a_61493_51596# sar10b_0.net1 0.0698f
C5624 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A 0.02842f
C5625 w_n9655_56533# VINN 0.08726f
C5626 VDDA a_n8277_65767# 0.05067f
C5627 c1_10156_97972# VCM 0.01358f
C5628 m3_36652_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C5629 m3_45124_37258# m3_45124_36138# 0.29566f
C5630 VDDD sar10b_0._16_ 0.59031f
C5631 VSSR c1_n1140_80052# 0.04956f
C5632 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A 0.28117f
C5633 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.03718f
C5634 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN sar10b_0.SWN[9] 0.18315f
C5635 m3_22532_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.07708f
C5636 sar10b_0.net41 sar10b_0.net42 1.07874f
C5637 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP a_38665_5788# 0.21556f
C5638 VSSA VINN 8.94434f
C5639 sar10b_0.net33 sar10b_0.net32 0.08492f
C5640 a_63339_48621# sar10b_0.SWN[4] 0.01329f
C5641 c1_14392_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C5642 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 4.35595f
C5643 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VSSR 5.18022f
C5644 a_63273_61671# sar10b_0.net11 0.02063f
C5645 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.07183f
C5646 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.01751f
C5647 c1_3096_21618# m3_4176_21578# 0.15596f
C5648 m3_45124_56298# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C5649 VDDD a_62527_56974# 0.18552f
C5650 a_65045_59588# sar10b_0.net12 0.01145f
C5651 tdc_0.OUTP sar10b_0.net2 0.11057f
C5652 a_60690_70625# a_61131_70891# 0.02852f
C5653 a_64245_59307# a_64705_59595# 0.26257f
C5654 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A 0.41861f
C5655 CLK EN 0.50413f
C5656 m3_5588_97932# c1_5920_97972# 1.74381f
C5657 VSSR m3_45124_46218# 0.63261f
C5658 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[7] 0.17717f
C5659 sar10b_0.net16 a_67077_57628# 0.17416f
C5660 sar10b_0.clk_div_0.COUNT\[1\] a_66785_50875# 0.01774f
C5661 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C5662 a_60843_52216# a_61182_52404# 0.07649f
C5663 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VCM 1.23381f
C5664 c1_n1140_22738# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C5665 m3_22532_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.53626f
C5666 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A 1.37544f
C5667 VSSD a_64492_67433# 0.29439f
C5668 a_65390_69010# sar10b_0.net43 0.02184f
C5669 a_62709_63063# a_63374_62684# 0.19065f
C5670 a_62985_63003# a_63509_62783# 0.04522f
C5671 a_n4470_53722# CLK 0.02136f
C5672 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A sar10b_0.CF[0] 0.02149f
C5673 m3_45124_77772# m3_45124_76652# 0.29566f
C5674 VSSR m3_45124_86732# 0.63305f
C5675 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.41496f
C5676 a_60693_57975# sar10b_0.net16 0.21836f
C5677 sar10b_0.CF[1] sar10b_0.SWP[0] 0.12129f
C5678 VDDD a_60747_57571# 0.29517f
C5679 m3_45124_30538# VDDR 0.0103f
C5680 VDDD a_67445_61451# 0.21684f
C5681 a_65861_51977# sar10b_0._04_ 0.36266f
C5682 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C5683 VDDD a_64338_52411# 0.24617f
C5684 m3_n1472_93452# c1_n1140_93492# 1.74381f
C5685 m3_45124_94572# c1_45456_93492# 0.01078f
C5686 VSSR c1_45456_95732# 0.0935f
C5687 a_64543_62648# VSSD 0.27764f
C5688 sar10b_0.SWN[0] VSSD 1.19492f
C5689 VDDD a_66933_59067# 0.32759f
C5690 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_26768_21578# 0.0162f
C5691 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_43712_21578# 0.03017f
C5692 CLK tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A 0.09504f
C5693 a_51603_58977# VSSA 0.06774f
C5694 VDDD a_64667_51628# 0.01557f
C5695 c1_28512_21618# VCM 0.01358f
C5696 c1_45456_39538# m3_45124_40618# 0.01078f
C5697 c1_45456_40658# m3_45124_39498# 0.01078f
C5698 c1_n1140_39538# m3_n1472_39498# 1.74381f
C5699 VDDD a_64907_50292# 0.01693f
C5700 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 4.10362f
C5701 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y 0.3196f
C5702 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 0.02632f
C5703 m3_45124_67692# th_dif_sw_0.VCP 0.17339f
C5704 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 0.02666f
C5705 m3_45124_71052# VDDR 0.01034f
C5706 VSSR th_dif_sw_0.VCP 0.11971p
C5707 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] th_dif_sw_0.VCN 70.5858f
C5708 a_65761_58263# a_65966_58354# 0.09983f
C5709 m3_31004_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.53746f
C5710 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.40249f
C5711 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A 0.03718f
C5712 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A 0.42509f
C5713 sar10b_0.net9 a_62185_62031# 0.22973f
C5714 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 sar10b_0.CF[9] 0.40665f
C5715 sar10b_0.net30 a_61400_50300# 0.01771f
C5716 sar10b_0.clknet_1_1__leaf_CLK sar10b_0.net16 0.05886f
C5717 VDDD a_61153_67587# 0.26824f
C5718 sar10b_0.net13 a_65525_68912# 0.03733f
C5719 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[3] 0.01887f
C5720 VDDD DATA[1] 0.3348f
C5721 VDDD a_65481_59303# 0.35394f
C5722 a_68169_65667# a_68767_65312# 0.06623f
C5723 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 2.7692f
C5724 sar10b_0.cyclic_flag_0.FINAL a_67209_65667# 0.26311f
C5725 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VDDR 4.94629f
C5726 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 2.16373f
C5727 m3_45124_62092# c1_45456_62132# 1.74381f
C5728 VSSR c1_45456_52978# 0.09348f
C5729 a_61493_58256# sar10b_0.net38 0.02118f
C5730 sar10b_0.net4 sar10b_0.CF[0] 0.09104f
C5731 VDDD a_67598_54692# 0.27387f
C5732 m3_n1472_94572# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C5733 m3_28180_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.96307f
C5734 sar10b_0.SWP[8] a_69003_71265# 0.1431f
C5735 sar10b_0._08_ a_64907_50292# 0.01511f
C5736 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.01132f
C5737 c1_n1140_78932# c1_n1140_77812# 0.13255f
C5738 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP sar10b_0.CF[3] 0.16021f
C5739 m3_28180_21578# c1_27100_21618# 0.15596f
C5740 m3_n1472_31658# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C5741 sar10b_0.net33 a_65589_57735# 0.01912f
C5742 VDDD sar10b_0.net3 13.0673f
C5743 a_61400_50300# VSSD 0.84835f
C5744 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN 0.01212f
C5745 a_66254_69344# a_66389_69443# 0.35559f
C5746 a_65865_69663# a_67077_69616# 0.07766f
C5747 m3_36652_97932# c1_35572_97972# 0.15596f
C5748 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 0.24487f
C5749 VSSD a_61609_62270# 0.10001f
C5750 VSSR m3_n1472_21578# 0.71232f
C5751 sar10b_0.net47 a_67423_69308# 0.2891f
C5752 sar10b_0.net1 tdc_0.OUTN 0.11225f
C5753 sar10b_0.net7 a_60969_51311# 0.03679f
C5754 sar10b_0.SWN[0] sar10b_0.CF[8] 0.18518f
C5755 c1_45456_37298# VDDR 0.01151f
C5756 c1_44044_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.01078f
C5757 m3_45124_40618# th_dif_sw_0.VCN 0.17339f
C5758 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 a_1127_5779# 0.04962f
C5759 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45324f
C5760 VSSD a_61677_66174# 0.13539f
C5761 a_68169_63003# a_68767_62648# 0.06623f
C5762 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45324f
C5763 sar10b_0.clk_div_0.COUNT\[0\] a_65577_51311# 0.03775f
C5764 sar10b_0.net29 EN 0.05412f
C5765 VDDR sar10b_0.SWN[2] 3.12286f
C5766 VDDD sar10b_0.SWP[0] 0.33534f
C5767 sar10b_0.net34 a_65355_53949# 0.07741f
C5768 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 0.02632f
C5769 c1_22864_21618# th_dif_sw_0.VCN 0.13255f
C5770 VSSR m3_n1472_62092# 0.74277f
C5771 sar10b_0.net3 sar10b_0._08_ 0.24909f
C5772 c1_45456_44018# c1_45456_42898# 0.13255f
C5773 VSSR a_24259_5788# 0.06033f
C5774 m3_18296_21578# VCM 0.13579f
C5775 sar10b_0.clk_div_0.COUNT\[0\] a_67543_51991# 0.02076f
C5776 c1_n1140_64372# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C5777 m3_45124_45098# m3_45124_43978# 0.29566f
C5778 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A 0.42509f
C5779 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A sar10b_0.CF[9] 0.06369f
C5780 sar10b_0.net17 sar10b_0.SWN[2] 0.06272f
C5781 VDDD a_64609_64923# 0.22523f
C5782 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 0.51491f
C5783 VDDD a_67798_52206# 0.08326f
C5784 th_dif_sw_0.VCN sar10b_0.CF[9] 0.33314f
C5785 a_61454_53360# VSSD 0.13439f
C5786 c1_11568_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.26825f
C5787 a_67445_60119# sar10b_0.net3 0.15999f
C5788 a_66368_52081# a_66666_51977# 0.02614f
C5789 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A 0.04073f
C5790 a_61153_58263# a_61358_58354# 0.09983f
C5791 a_62181_58100# a_61929_57971# 0.27388f
C5792 VDDD a_66666_49313# 0.09155f
C5793 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP 3.55945f
C5794 c1_n1140_38418# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C5795 VCM sar10b_0.CF[3] 3.51491f
C5796 sar10b_0.SWP[5] sar10b_0.CF[9] 0.17387f
C5797 VDDA a_51603_61205# 0.01057f
C5798 VDDD a_61086_64638# 0.31749f
C5799 sar10b_0.SWP[9] sar10b_0.net15 0.01984f
C5800 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 0.26289f
C5801 sar10b_0.net38 a_63273_56639# 0.02495f
C5802 sar10b_0.net33 a_66062_57022# 0.02934f
C5803 VDDD a_66537_57971# 0.38048f
C5804 VSSR c1_n1140_28338# 0.04956f
C5805 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C5806 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VDDR 6.1813f
C5807 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y 0.32264f
C5808 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.21001f
C5809 a_61400_63620# sar10b_0.net16 0.1331f
C5810 VINN th_dif_sw_0.VCN 3.18189f
C5811 a_61419_48621# VSSD 0.28994f
C5812 m3_45124_71052# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C5813 a_65682_49313# a_66109_49318# 0.04602f
C5814 m3_45124_85612# m3_45124_84492# 0.29566f
C5815 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A 0.11547f
C5816 VSSR m3_33828_97932# 0.52359f
C5817 VDDD a_62933_58787# 0.204f
C5818 m3_33828_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.75703f
C5819 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VCM 3.62379f
C5820 m3_45124_46218# VDDR 0.0103f
C5821 a_61496_52091# sar10b_0.net1 0.01817f
C5822 VSSA tdc_0.phase_detector_0.pd_out_0.B 1.34879f
C5823 sar10b_0.SWN[5] a_20335_5779# 0.40667f
C5824 a_64238_63682# VSSD 0.16485f
C5825 VDDD a_67598_64016# 0.27393f
C5826 a_67209_59007# a_67733_58787# 0.04522f
C5827 a_62181_51440# sar10b_0.net16 0.17435f
C5828 a_66933_59067# a_67598_58688# 0.19065f
C5829 a_61358_67678# sar10b_0.net16 0.25048f
C5830 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A 0.41861f
C5831 VSSR c1_11568_97972# 0.05685f
C5832 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A 0.84106f
C5833 a_61454_50696# VSSD 0.13438f
C5834 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 1.80961f
C5835 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_4176_21578# 0.03017f
C5836 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 0.02632f
C5837 c1_1684_21618# VCM 0.01358f
C5838 c1_n1140_47378# m3_n1472_47338# 1.74381f
C5839 c1_45456_48498# m3_45124_47338# 0.01078f
C5840 c1_45456_47378# m3_45124_48458# 0.01078f
C5841 a_63804_67580# a_64238_67295# 0.17477f
C5842 VDDD a_61086_60642# 0.31562f
C5843 a_62181_58100# sar10b_0.net4 0.05003f
C5844 a_60747_63273# a_60945_63273# 0.06623f
C5845 m3_45124_86732# VDDR 0.01034f
C5846 m3_45124_83372# th_dif_sw_0.VCP 0.17339f
C5847 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR 0.38716f
C5848 VDDD a_62949_56296# 0.27318f
C5849 sar10b_0.net33 sar10b_0.net40 0.02534f
C5850 th_dif_sw_0.th_sw_1.CKB a_n8277_66083# 0.06592f
C5851 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN 0.01239f
C5852 a_60747_65937# a_61086_65970# 0.07649f
C5853 a_61395_65944# a_60945_65937# 0.03508f
C5854 tdc_0.RDY sar10b_0.CF[3] 0.14563f
C5855 a_67372_52243# sar10b_0.clk_div_0.COUNT\[0\] 0.06299f
C5856 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP 0.18415f
C5857 c1_45456_95732# VDDR 0.01153f
C5858 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A 0.04073f
C5859 c1_31336_97972# VCM 0.01358f
C5860 sar10b_0.net8 a_62313_61671# 0.23697f
C5861 sar10b_0.net3 a_68133_61624# 0.18332f
C5862 m3_n1472_68812# c1_n1140_69972# 0.01078f
C5863 m3_n1472_69932# c1_n1140_68852# 0.01078f
C5864 m3_45124_69932# c1_45456_69972# 1.74381f
C5865 a_55121_59650# tdc_0.OUTP 0.05224f
C5866 sar10b_0.clknet_0_CLK VSSD 2.12126f
C5867 VSSR c1_45456_72212# 0.0935f
C5868 m3_12648_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.31585f
C5869 c1_35572_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C5870 a_68421_68284# VSSD 0.27202f
C5871 m3_26768_97932# m3_28180_97932# 0.23959f
C5872 a_67598_58688# sar10b_0.net3 0.25973f
C5873 a_60693_51315# a_61153_51603# 0.26257f
C5874 th_dif_sw_0.VCP VDDR 0.66159f
C5875 sar10b_0.net36 a_68946_56639# 0.01509f
C5876 a_61493_67580# a_61929_67295# 0.16939f
C5877 a_60969_67295# a_61358_67678# 0.06034f
C5878 c1_14392_21618# m3_14060_21578# 1.74381f
C5879 c1_n1140_86772# c1_n1140_85652# 0.13255f
C5880 m3_n1472_47338# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C5881 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A sar10b_0.CF[1] 0.03041f
C5882 VDDD a_64831_56974# 0.1958f
C5883 sar10b_0.net16 a_62497_61303# 0.08934f
C5884 sar10b_0.net46 sar10b_0.net15 0.09997f
C5885 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VCM 1.16928f
C5886 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A a_51861_60437# 0.16495f
C5887 a_67310_60020# VSSD 0.1297f
C5888 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[3] 0.05939f
C5889 sar10b_0.net28 CLK 0.07871f
C5890 m3_16884_97932# c1_15804_97972# 0.15596f
C5891 VSSR m3_n1472_37258# 0.66371f
C5892 sar10b_0.CF[1] sar10b_0.SWP[1] 2.74424f
C5893 sar10b_0.SWP[0] sar10b_0.CF[2] 0.12314f
C5894 a_60693_67299# sar10b_0.net4 0.04972f
C5895 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VDDR 2.57696f
C5896 c1_45456_52978# VDDR 0.01151f
C5897 VSSA a_52504_60961# 0.01123f
C5898 m3_45124_56298# th_dif_sw_0.VCN 0.17719f
C5899 m3_43712_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C5900 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y VSSR 0.32296f
C5901 sar10b_0.CF[6] sar10b_0.SWN[2] 0.12251f
C5902 sar10b_0.SWN[1] sar10b_0.SWN[2] 9.06444f
C5903 VSSR c1_29924_21618# 0.05685f
C5904 a_64814_65014# sar10b_0.net16 0.27418f
C5905 sar10b_0.CF[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.12367f
C5906 a_67393_54643# a_68421_54964# 0.07826f
C5907 a_65865_57675# a_65589_57735# 0.1263f
C5908 VSSR m3_n1472_77772# 0.66316f
C5909 sar10b_0.net33 sar10b_0.net38 0.02409f
C5910 VDDD a_60843_52216# 0.22279f
C5911 a_53652_61050# tdc_0.phase_detector_0.pd_out_0.B 0.18921f
C5912 c1_45456_51858# c1_45456_50738# 0.13255f
C5913 sar10b_0.net3 a_68169_55011# 0.27649f
C5914 sar10b_0.net34 a_66197_56924# 0.01805f
C5915 a_61921_55975# a_62126_56024# 0.09983f
C5916 m3_n1472_21578# VDDR 0.02681f
C5917 w_n9655_63119# a_n4470_65264# 0.01216f
C5918 sar10b_0.SWN[8] VSSD 0.81908f
C5919 sar10b_0.net8 a_62702_61352# 0.03629f
C5920 m3_n1472_29418# VCM 0.01415f
C5921 c1_n1140_80052# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C5922 DATA[2] sar10b_0.net36 0.13468f
C5923 m3_45124_52938# m3_45124_51818# 0.29566f
C5924 a_68767_62648# VSSD 0.26814f
C5925 VDDD a_65861_51977# 0.79975f
C5926 sar10b_0.net2 a_64238_67295# 0.0126f
C5927 a_44345_5779# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A 0.01247f
C5928 sar10b_0.clk_div_0.COUNT\[2\] a_68178_51635# 0.15252f
C5929 a_61705_51992# sar10b_0.net16 0.1642f
C5930 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSSR 0.41774f
C5931 m3_n1472_62092# VDDR 0.02674f
C5932 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C5933 m3_n1472_69932# VCM 0.01412f
C5934 VDDD a_68169_65667# 0.36668f
C5935 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A 0.43651f
C5936 sar10b_0.CF[1] th_dif_sw_0.CK 0.08524f
C5937 a_63573_63303# a_63849_63299# 0.1263f
C5938 sar10b_0.net7 a_61182_52404# 0.01042f
C5939 VDDR a_24259_5788# 4.81771f
C5940 a_65857_56931# a_66885_56768# 0.07826f
C5941 sar10b_0.SWN[9] VSSD 1.25116f
C5942 a_9853_5788# VSSR 0.06033f
C5943 c1_n1140_54098# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C5944 sar10b_0.net32 sar10b_0._01_ 0.03898f
C5945 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 0.40575f
C5946 sar10b_0.CF[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP 0.17518f
C5947 VSSD a_67881_61671# 0.28968f
C5948 c1_29924_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.26825f
C5949 a_65589_69723# sar10b_0.net16 0.2698f
C5950 a_65961_68627# a_66559_68962# 0.06623f
C5951 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] th_dif_sw_0.VCN 35.0616f
C5952 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y VSSR 0.32264f
C5953 VSSR c1_n1140_44018# 0.04956f
C5954 sar10b_0.SWP[3] sar10b_0.CF[3] 2.41685f
C5955 a_67393_58639# VSSD 0.85489f
C5956 m3_45124_86732# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C5957 a_66312_50368# a_66205_50408# 0.14439f
C5958 m3_45124_93452# m3_45124_92332# 0.29566f
C5959 a_68946_49747# DATA[1] 0.14753f
C5960 sar10b_0.net34 a_67371_49579# 0.28615f
C5961 a_68178_51635# VSSD 0.16529f
C5962 m3_38064_21578# c1_38396_21618# 1.74381f
C5963 sar10b_0.clknet_1_1__leaf_CLK a_65682_51977# 0.24324f
C5964 m3_45124_23818# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C5965 a_60945_63273# VSSD 0.28732f
C5966 VDDD sar10b_0.SWP[1] 2.88437f
C5967 sar10b_0.SWP[4] a_63339_71265# 0.01261f
C5968 sar10b_0.SWN[8] sar10b_0.CF[8] 2.36938f
C5969 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP 3.71029f
C5970 a_64705_59595# sar10b_0.net11 0.01555f
C5971 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 2.74312f
C5972 a_63273_56639# a_63457_56931# 0.44532f
C5973 m3_45124_97932# c1_45456_96852# 0.01078f
C5974 m3_45124_96812# c1_45456_97972# 0.01078f
C5975 m3_n1472_96812# c1_n1140_96852# 1.74381f
C5976 VSSR m3_19708_21578# 0.40111f
C5977 a_15533_5779# sar10b_0.SWN[6] 0.32874f
C5978 a_61153_51603# VSSD 0.83916f
C5979 a_61929_67295# VSSD 0.28544f
C5980 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y 0.3196f
C5981 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.14338f
C5982 c1_n1140_55218# m3_n1472_55178# 1.74381f
C5983 c1_45456_56338# m3_45124_55178# 0.01078f
C5984 c1_45456_55218# m3_45124_56298# 0.01078f
C5985 th_dif_sw_0.VCP a_51345_60437# 0.06502f
C5986 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 1.10485p
C5987 VSSD a_64533_65967# 0.14563f
C5988 a_61677_50190# sar10b_0.net1 0.01536f
C5989 a_60945_49953# a_61609_50282# 0.16939f
C5990 sar10b_0.cyclic_flag_0.FINAL a_67209_68331# 0.22988f
C5991 sar10b_0.net28 sar10b_0.net29 0.04415f
C5992 m3_14060_97932# VCM 0.13579f
C5993 a_61395_52624# sar10b_0.net16 0.25365f
C5994 c1_44044_21618# th_dif_sw_0.VCN 0.13255f
C5995 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_35572_21618# 0.0106f
C5996 sar10b_0.net33 a_66109_49318# 0.01476f
C5997 sar10b_0.net8 a_62185_60699# 0.18642f
C5998 sar10b_0.net14 a_66021_66092# 0.01301f
C5999 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP a_24259_109594# 0.14286f
C6000 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y 0.07418f
C6001 sar10b_0.net2 sar10b_0.CF[1] 0.01023f
C6002 c1_20040_97972# th_dif_sw_0.VCP 0.13255f
C6003 VDDD a_63804_67580# 0.2086f
C6004 sar10b_0.net4 a_61065_53679# 0.25127f
C6005 sar10b_0.net2 a_61677_62178# 0.0202f
C6006 m3_39476_21578# VCM 0.15231f
C6007 m3_18296_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C6008 a_68946_53975# DATA[3] 0.1474f
C6009 sar10b_0.net1 sar10b_0.net12 0.58065f
C6010 sar10b_0.clknet_1_1__leaf_CLK sar10b_0._07_ 0.26895f
C6011 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP sar10b_0.SWP[7] 0.20251f
C6012 m3_n1472_77772# c1_n1140_76692# 0.01078f
C6013 m3_n1472_76652# c1_n1140_77812# 0.01078f
C6014 a_67564_50907# a_68035_50645# 0.01114f
C6015 m3_45124_77772# c1_45456_77812# 1.74381f
C6016 VSSR c1_45456_87892# 0.0935f
C6017 sar10b_0.CF[6] th_dif_sw_0.VCP 0.28583f
C6018 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSSR 33.417f
C6019 a_68169_64335# sar10b_0.net3 0.27548f
C6020 a_64773_60292# VSSD 0.26534f
C6021 sar10b_0.SWP[4] VCM 0.13076f
C6022 VSSD a_66885_56768# 0.26821f
C6023 VDDD sar10b_0.net5 1.73087f
C6024 m3_7000_97932# m3_8412_97932# 0.23959f
C6025 a_64949_64916# a_65385_64631# 0.16939f
C6026 c1_45456_23858# m3_45124_23818# 1.74381f
C6027 c1_n1140_23858# m3_n1472_22698# 0.01078f
C6028 c1_n1140_22738# m3_n1472_23818# 0.01078f
C6029 sar10b_0.net40 a_65865_57675# 0.05453f
C6030 sar10b_0.net21 a_68767_54656# 0.01278f
C6031 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A 0.10815f
C6032 sar10b_0.net33 sar10b_0.net14 0.52388f
C6033 a_64773_60292# a_63561_60339# 0.07766f
C6034 VDDD th_dif_sw_0.CK 0.55496f
C6035 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 1.05065f
C6036 a_61419_48621# sar10b_0.SWN[0] 0.16109f
C6037 a_61773_52237# sar10b_0.net16 0.27952f
C6038 VDDD a_65996_50650# 0.0194f
C6039 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VSSR 1.37836f
C6040 VDDD a_64197_62956# 0.26772f
C6041 VSSR m3_n1472_52938# 0.66371f
C6042 a_67209_68331# a_67393_67963# 0.44098f
C6043 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.2477f
C6044 VDDD sar10b_0._00_ 0.5815f
C6045 sar10b_0.net9 a_62985_63003# 0.20758f
C6046 c1_45456_72212# VDDR 0.01153f
C6047 a_61491_52222# sar10b_0.net6 0.01139f
C6048 m3_4176_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C6049 a_64149_64635# sar10b_0.net11 0.04964f
C6050 m3_32416_21578# m3_33828_21578# 0.23959f
C6051 a_68235_48621# VSSD 0.30699f
C6052 sar10b_0.net21 sar10b_0.net37 0.98928f
C6053 VSSR c1_3096_21618# 0.05923f
C6054 a_61833_57675# a_61557_57735# 0.1263f
C6055 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17717f
C6056 m3_n1472_62092# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24058f
C6057 a_65577_57971# a_66537_57971# 0.03432f
C6058 sar10b_0._10_ a_65188_51977# 0.02387f
C6059 VSSR m3_n1472_93452# 0.66316f
C6060 c1_45456_63252# c1_45456_62132# 0.13255f
C6061 a_65385_64631# VSSD 0.29549f
C6062 VSSR sar10b_0.SWP[0] 7.11885f
C6063 m3_n1472_37258# VDDR 0.02681f
C6064 a_65185_68919# sar10b_0.net16 0.27947f
C6065 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] sar10b_0.SWP[4] 0.2309f
C6066 m3_n1472_45098# VCM 0.01415f
C6067 sar10b_0.net17 a_64818_49979# 0.05106f
C6068 VINN a_n9133_57045# 0.01178f
C6069 a_65301_57975# VSSD 0.14241f
C6070 a_68421_58960# a_68767_58652# 0.07649f
C6071 VSSR c1_32748_97972# 0.06914f
C6072 a_61395_64612# a_62185_64695# 0.1263f
C6073 a_61400_64952# a_61609_64934# 0.24088f
C6074 sar10b_0._08_ sar10b_0._00_ 0.23008f
C6075 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] m3_21120_97932# 0.26476f
C6076 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A 0.11547f
C6077 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y VDDR 0.31995f
C6078 VDDD sar10b_0._06_ 0.66501f
C6079 sar10b_0.cyclic_flag_0.FINAL a_66921_61671# 0.22764f
C6080 sar10b_0.net23 a_68946_63299# 0.01265f
C6081 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_8412_21578# 0.0162f
C6082 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_25356_21578# 0.03017f
C6083 a_68562_49747# VSSD 0.31698f
C6084 VSSA a_n8277_66083# 22.0777f
C6085 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A 0.07418f
C6086 VDDD a_61086_49986# 0.31167f
C6087 VSSD a_61609_64934# 0.10006f
C6088 a_64910_59686# sar10b_0.net16 0.256f
C6089 m3_n1472_77772# VDDR 0.02674f
C6090 c1_20040_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 0.01078f
C6091 m3_12648_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.53746f
C6092 sar10b_0.net9 a_62185_60699# 0.03249f
C6093 m3_n1472_85612# VCM 0.01412f
C6094 a_67372_52243# sar10b_0._03_ 0.02316f
C6095 VDDD sar10b_0.net2 6.04238f
C6096 sar10b_0.net34 sar10b_0._04_ 0.0272f
C6097 c1_n1140_27218# c1_n1140_26098# 0.13255f
C6098 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.11339f
C6099 a_63369_59007# VSSD 0.283f
C6100 VDDD a_61609_66266# 0.20839f
C6101 a_67209_65667# a_67733_65447# 0.04522f
C6102 a_66933_65727# a_67598_65348# 0.19065f
C6103 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 11.9058f
C6104 m3_n1472_28298# m3_n1472_27178# 0.29566f
C6105 VSSR c1_n1140_63252# 0.04956f
C6106 a_65061_63428# sar10b_0.net12 0.01801f
C6107 sar10b_0.CF[2] sar10b_0.SWP[1] 0.12037f
C6108 VDDD sar10b_0.clk_div_0.COUNT\[3\] 0.55903f
C6109 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR 0.38377f
C6110 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A 0.41861f
C6111 m3_33828_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.75703f
C6112 a_67393_63967# a_68421_64288# 0.07826f
C6113 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A 1.37577f
C6114 sar10b_0.net47 VSSD 1.3254f
C6115 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A 0.38427f
C6116 sar10b_0.CF[9] sar10b_0.SWP[6] 0.16685f
C6117 a_61249_53311# a_61589_53459# 0.24088f
C6118 m3_45124_39498# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C6119 sar10b_0.net7 sar10b_0.CF[1] 0.18315f
C6120 m3_19708_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.09361f
C6121 VSSD a_61609_60938# 0.08276f
C6122 a_66795_71265# sar10b_0.net44 0.26209f
C6123 a_9853_5788# VDDR 2.42521f
C6124 a_60969_56639# a_61153_56931# 0.44532f
C6125 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 1.41356f
C6126 m3_26768_97932# c1_27100_97972# 1.74381f
C6127 a_65769_65963# a_66367_66298# 0.06623f
C6128 a_61065_53679# a_60789_53739# 0.1263f
C6129 VSSR m3_45124_29418# 0.63261f
C6130 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 0.01367f
C6131 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y VDDR 0.3196f
C6132 a_68479_59984# sar10b_0.net23 0.01248f
C6133 a_66933_67059# a_67393_66631# 0.26257f
C6134 a_67209_66999# a_67598_66680# 0.05462f
C6135 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VSSR 2.73845f
C6136 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.03718f
C6137 sar10b_0.net33 sar10b_0.net13 0.03442f
C6138 a_61400_60956# a_61609_60938# 0.24088f
C6139 VDDD a_61249_53311# 0.2606f
C6140 a_62187_71265# sar10b_0.net40 0.26704f
C6141 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN sar10b_0.CF[9] 0.03488f
C6142 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_8744_21618# 0.0106f
C6143 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 2.76761f
C6144 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A 0.04073f
C6145 m3_n1472_68812# m3_n1472_67692# 0.29566f
C6146 VSSR m3_45124_69932# 0.63305f
C6147 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y sar10b_0.CF[7] 0.12541f
C6148 a_21040_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A 0.01076f
C6149 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y 0.07418f
C6150 sar10b_0.clknet_1_0__leaf_CLK a_65586_50645# 0.05317f
C6151 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A 1.11894f
C6152 m3_n60_21578# VCM 0.15231f
C6153 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN 0.02638f
C6154 m3_n1472_84492# c1_n1140_85652# 0.01078f
C6155 m3_45124_85612# c1_45456_85652# 1.74381f
C6156 m3_n1472_85612# c1_n1140_84532# 0.01078f
C6157 th_dif_sw_0.CK sar10b_0.CF[2] 0.08539f
C6158 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C6159 sar10b_0.clknet_1_1__leaf_CLK a_65394_52643# 0.29811f
C6160 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.95164f
C6161 VDDD a_61035_48621# 0.25976f
C6162 sar10b_0.net19 DATA[4] 0.01539f
C6163 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 3.7115f
C6164 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A 0.41861f
C6165 c1_45456_31698# m3_45124_31658# 1.74381f
C6166 c1_n1140_31698# m3_n1472_30538# 0.01078f
C6167 c1_n1140_30578# m3_n1472_31658# 0.01078f
C6168 VSSA a_51345_58977# 0.4784f
C6169 sar10b_0.SWP[4] sar10b_0.SWP[3] 12.5824f
C6170 VDDD a_65407_63634# 0.21226f
C6171 sar10b_0.net16 a_65966_58354# 0.24295f
C6172 sar10b_0.SWP[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 0.3013f
C6173 a_68169_66999# a_68421_66952# 0.27388f
C6174 VDDD a_61249_50647# 0.25603f
C6175 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 0.12358f
C6176 a_61491_52222# VSSD 0.48779f
C6177 c1_45456_87892# VDDR 0.01153f
C6178 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A 0.28117f
C6179 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VDDR 8.23921f
C6180 m3_12648_21578# m3_14060_21578# 0.23959f
C6181 VSSD a_63045_57628# 0.25727f
C6182 VSSR c1_45456_36178# 0.09348f
C6183 CLK sar10b_0.CF[9] 0.10704f
C6184 a_61249_50647# a_61589_50795# 0.24088f
C6185 a_61065_51015# a_62025_51015# 0.03529f
C6186 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A sar10b_0.CF[3] 0.06369f
C6187 sar10b_0.net34 a_66593_50645# 0.02136f
C6188 m3_n1472_77772# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C6189 VDDD sar10b_0.net7 2.2805f
C6190 sar10b_0.net14 a_65865_57675# 0.02761f
C6191 VSSR m3_15472_97932# 0.44987f
C6192 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VDDR 0.83559f
C6193 c1_45456_71092# c1_45456_69972# 0.13255f
C6194 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.55567p
C6195 m3_15472_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.2724f
C6196 sar10b_0.SWN[2] sar10b_0.CF[7] 0.12695f
C6197 m3_n1472_52938# VDDR 0.02681f
C6198 VDDD a_65355_53949# 1.5132f
C6199 VDDA th_dif_sw_0.th_sw_1.CKB 2.79588f
C6200 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] 7.81593f
C6201 VSSR m3_40888_21578# 0.54637f
C6202 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP sar10b_0.SWN[5] 0.24476f
C6203 a_64245_59307# sar10b_0.net16 0.28698f
C6204 sar10b_0.CF[5] sar10b_0.CF[9] 0.1103f
C6205 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A sar10b_0.CF[3] 0.03041f
C6206 sar10b_0.SWP[8] VDDA 0.24929f
C6207 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.21974f
C6208 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C6209 VDDD a_68169_68331# 0.36685f
C6210 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A 0.02842f
C6211 m3_45124_23818# th_dif_sw_0.VCN 0.17339f
C6212 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VCM 2.64983f
C6213 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VCM 3.87097f
C6214 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP a_29939_5779# 0.01299f
C6215 sar10b_0.net14 a_65961_68627# 0.02371f
C6216 sar10b_0.net33 a_65586_50645# 0.0296f
C6217 m3_n1472_93452# VDDR 0.02674f
C6218 VDDD a_67105_59971# 0.27834f
C6219 VDDR sar10b_0.SWP[0] 3.85632f
C6220 VDDD a_68946_56639# 0.28035f
C6221 sar10b_0._01_ CLK 0.01823f
C6222 m3_35240_97932# VCM 0.15231f
C6223 sar10b_0.net3 sar10b_0.net17 0.3001f
C6224 sar10b_0.net43 VSSD 1.84798f
C6225 c1_n1140_35058# c1_n1140_33938# 0.13255f
C6226 m3_45124_55178# sar10b_0.CF[0] 0.01071f
C6227 sar10b_0.net3 a_67598_66680# 0.25604f
C6228 VDDD a_66837_56403# 0.33237f
C6229 a_65394_52643# a_65821_53072# 0.04602f
C6230 a_61929_51311# sar10b_0.net1 0.0614f
C6231 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] VSSR 18.4213f
C6232 c1_12980_97972# VCM 0.01358f
C6233 m3_39476_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C6234 m3_n1472_36138# m3_n1472_35018# 0.29566f
C6235 VSSR c1_n1140_78932# 0.04956f
C6236 m3_25356_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.57708f
C6237 sar10b_0.net46 a_66254_69344# 0.01964f
C6238 sar10b_0.SWN[3] sar10b_0.SWN[4] 12.5823f
C6239 c1_17216_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C6240 c1_4508_21618# m3_5588_21578# 0.15596f
C6241 a_62025_53679# sar10b_0.net16 0.26997f
C6242 m3_45124_55178# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C6243 a_65185_68919# a_65390_69010# 0.09983f
C6244 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A 0.39559f
C6245 a_61131_70891# sar10b_0.net38 0.24738f
C6246 a_64521_59303# a_65045_59588# 0.05022f
C6247 sar10b_0.CF[0] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 0.10544f
C6248 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] 1.63975f
C6249 VDDD a_68421_62956# 0.27523f
C6250 VINP w_n9655_63119# 0.08726f
C6251 m3_7000_97932# c1_7332_97972# 1.74381f
C6252 VSSR m3_45124_45098# 0.63261f
C6253 a_54372_59599# tdc_0.OUTP 0.01017f
C6254 a_68169_68331# a_68767_67976# 0.06623f
C6255 a_51603_58977# CLK 0.02753f
C6256 VSSR sar10b_0.SWP[1] 5.94102f
C6257 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A sar10b_0.CF[2] 0.02149f
C6258 a_61041_52340# a_61491_52222# 0.03432f
C6259 VDDD DATA[2] 0.44638f
C6260 m3_25356_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C6261 VSSD a_64888_67630# 0.42371f
C6262 a_63169_62635# a_63374_62684# 0.09983f
C6263 a_61929_57971# sar10b_0.net40 0.01233f
C6264 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A sar10b_0.CF[7] 0.26294f
C6265 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A 0.02842f
C6266 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A sar10b_0.SWN[0] 0.02058f
C6267 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP a_43467_106170# 0.23957f
C6268 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A 0.83994f
C6269 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 5.3129f
C6270 a_67209_55011# a_66933_55071# 0.1263f
C6271 m3_n1472_76652# m3_n1472_75532# 0.29566f
C6272 a_61153_58263# sar10b_0.net16 0.08375f
C6273 VSSR m3_45124_85612# 0.63305f
C6274 a_67105_59971# a_67445_60119# 0.24088f
C6275 a_66921_60339# a_68133_60292# 0.07766f
C6276 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A 1.34717f
C6277 m3_45124_29418# VDDR 0.0103f
C6278 a_62025_51015# sar10b_0.net16 0.27023f
C6279 a_67372_52833# sar10b_0._14_ 0.33036f
C6280 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN 4.82055f
C6281 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] sar10b_0.SWP[8] 0.22497f
C6282 VDDD sar10b_0._09_ 0.52059f
C6283 a_66785_50875# VSSD 0.5236f
C6284 m3_45124_93452# c1_45456_93492# 1.74381f
C6285 m3_n1472_92332# c1_n1140_93492# 0.01078f
C6286 m3_n1472_93452# c1_n1140_92372# 0.01078f
C6287 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.40249f
C6288 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VDDR 2.62306f
C6289 VSSR c1_45456_94612# 0.0935f
C6290 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP 0.02666f
C6291 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A sar10b_0.CF[2] 0.03041f
C6292 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_29592_21578# 0.0162f
C6293 sar10b_0.net32 a_64199_50761# 0.02376f
C6294 VINN th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 0.36273f
C6295 c1_31336_21618# VCM 0.01358f
C6296 VDDD a_61395_63280# 0.85861f
C6297 c1_45456_39538# m3_45124_39498# 1.74381f
C6298 c1_n1140_38418# m3_n1472_39498# 0.01078f
C6299 c1_n1140_39538# m3_n1472_38378# 0.01078f
C6300 a_67113_56343# a_67297_55975# 0.44098f
C6301 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] c1_20040_97972# 0.02068f
C6302 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.11339f
C6303 m3_45124_69932# VDDR 0.01034f
C6304 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y 0.07183f
C6305 m3_45124_66572# th_dif_sw_0.VCP 0.17339f
C6306 sar10b_0.net10 a_63573_63303# 0.0507f
C6307 th_dif_sw_0.VCP sar10b_0.CF[7] 0.28584f
C6308 VSSR cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 27.5187f
C6309 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VDDR 0.95338f
C6310 sar10b_0.net4 sar10b_0.net40 3.61184f
C6311 VDDD sar10b_0.net45 2.00128f
C6312 sar10b_0.CF[6] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] 0.01377f
C6313 sar10b_0.net32 sar10b_0._11_ 0.04846f
C6314 VSSR th_dif_sw_0.CK 11.5936f
C6315 th_dif_sw_0.CKB th_dif_sw_0.th_sw_1.CKB 0.07475f
C6316 VSSD a_67393_66631# 0.85332f
C6317 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VSSR 1.37482f
C6318 VDDD a_60969_51311# 0.81714f
C6319 sar10b_0.net7 sar10b_0.CF[2] 0.27698f
C6320 VDDD a_62181_67424# 0.26952f
C6321 a_64609_64923# sar10b_0.net12 0.0169f
C6322 a_66933_55071# sar10b_0.net35 0.02103f
C6323 sar10b_0._09_ sar10b_0._08_ 0.79396f
C6324 VDDD sar10b_0.net34 1.50082f
C6325 c1_11568_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.26825f
C6326 m3_n1472_57418# c1_n1140_57458# 1.74381f
C6327 VSSR c1_45456_51858# 0.09348f
C6328 sar10b_0._14_ sar10b_0.net35 0.02355f
C6329 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VDDR 2.68527f
C6330 VDDD tdc_0.OUTP 0.36938f
C6331 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A sar10b_0.CF[5] 0.26294f
C6332 VDDA sar10b_0.CF[0] 0.11532f
C6333 m3_n1472_93452# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C6334 m3_31004_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.53746f
C6335 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] sar10b_0.SWP[0] 0.2377f
C6336 c1_45456_78932# c1_45456_77812# 0.13255f
C6337 sar10b_0.net16 a_61461_56403# 0.25197f
C6338 m3_29592_21578# c1_28512_21618# 0.15596f
C6339 m3_n1472_30538# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C6340 a_60747_52617# sar10b_0.net5 0.28232f
C6341 th_dif_sw_0.VCN a_51345_58977# 0.06502f
C6342 sar10b_0.net19 sar10b_0.net22 0.76458f
C6343 a_61609_50282# VSSD 0.10006f
C6344 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] 3.0756f
C6345 tdc_0.RDY a_60690_53975# 0.19682f
C6346 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP 0.02666f
C6347 a_66049_69295# a_66825_69663# 0.3578f
C6348 m3_38064_97932# c1_36984_97972# 0.15596f
C6349 VSSR m3_1352_21578# 0.54637f
C6350 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VCM 0.12357f
C6351 sar10b_0.net46 a_65961_68627# 0.01772f
C6352 sar10b_0.SWP[9] sar10b_0.CF[9] 2.43738f
C6353 sar10b_0.net34 sar10b_0._08_ 0.0219f
C6354 VDDD a_64521_60339# 0.34849f
C6355 c1_18628_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.02523f
C6356 VDDD a_66197_56924# 0.20139f
C6357 c1_45456_36178# VDDR 0.01151f
C6358 m3_45124_39498# th_dif_sw_0.VCN 0.17339f
C6359 VSSD a_62185_66027# 0.15809f
C6360 sar10b_0.net3 a_60690_49683# 0.86891f
C6361 sar10b_0.CF[6] sar10b_0.SWP[0] 0.13213f
C6362 sar10b_0.SWN[3] VSSA 0.24827f
C6363 m3_23944_97932# th_dif_sw_0.VCP 0.01078f
C6364 sar10b_0._10_ sar10b_0.net16 0.38615f
C6365 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] a_19457_110450# 1.48701f
C6366 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP 2.92171f
C6367 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN sar10b_0.CF[3] 0.12378f
C6368 sar10b_0.net16 a_62997_56643# 0.25095f
C6369 VSSR m3_n1472_57418# 0.74361f
C6370 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 0.21577f
C6371 sar10b_0.net2 a_61677_60846# 0.01865f
C6372 c1_n1140_42898# c1_n1140_41778# 0.13255f
C6373 sar10b_0.SWN[9] sar10b_0.SWN[8] 21.3652f
C6374 sar10b_0.net38 sar10b_0.net4 0.12818f
C6375 m3_n60_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03808f
C6376 m3_21120_21578# VCM 0.6299f
C6377 sar10b_0.SWN[2] a_34741_5779# 0.64048f
C6378 c1_n1140_63252# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C6379 m3_n1472_43978# m3_n1472_42858# 0.29566f
C6380 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[4] 0.01887f
C6381 DATA[5] sar10b_0.net22 0.07431f
C6382 a_66666_51977# sar10b_0.net35 0.01391f
C6383 VDDA a_n8277_54249# 1.0219f
C6384 sar10b_0.SWN[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.45621f
C6385 sar10b_0.net3 sar10b_0.net41 0.13347f
C6386 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN 3.1317f
C6387 VDDD a_65637_64760# 0.2745f
C6388 a_n9133_63315# a_n8277_66083# 0.97211f
C6389 sar10b_0.net30 a_62187_48621# 0.25742f
C6390 sar10b_0.net39 sar10b_0.net16 2.69525f
C6391 sar10b_0.net3 sar10b_0.clk_div_0.COUNT\[0\] 0.15704f
C6392 VSSA a_53564_59480# 0.02937f
C6393 c1_14392_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.26836f
C6394 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] VDDR 2.16044f
C6395 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VCM 4.85259f
C6396 sar10b_0.net8 a_63273_56639# 0.20582f
C6397 a_61929_57971# a_62527_58306# 0.06623f
C6398 VDDD a_67371_49579# 0.27466f
C6399 c1_n1140_37298# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C6400 a_62185_63363# sar10b_0.net40 0.0117f
C6401 VSSR cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 94.3862f
C6402 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP sar10b_0.CF[7] 0.10502f
C6403 a_45050_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A 0.01076f
C6404 w_n9655_56533# VDDA 1.47643f
C6405 th_dif_sw_0.VCP th_dif_sw_0.th_sw_1.th_sw_main_0.VGS 0.09766f
C6406 sar10b_0.net3 a_67502_56024# 0.24317f
C6407 VSSD a_67077_57628# 0.27049f
C6408 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP 2.33876f
C6409 VDDD sar10b_0.net36 2.06897f
C6410 VSSR c1_n1140_27218# 0.04956f
C6411 sar10b_0.CF[4] VCM 3.51243f
C6412 a_63810_50901# a_63918_50969# 0.29821f
C6413 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y 0.07418f
C6414 a_61609_63602# sar10b_0.net16 0.20179f
C6415 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A 0.60057f
C6416 a_62187_48621# VSSD 0.34304f
C6417 m3_45124_69932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C6418 VDDA VSSA 0.63221p
C6419 a_65861_49313# a_66368_49417# 0.21226f
C6420 a_65682_49313# a_66216_49358# 0.35097f
C6421 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A 0.39629f
C6422 m3_n1472_84492# m3_n1472_83372# 0.29566f
C6423 VSSR m3_36652_97932# 0.54637f
C6424 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 2.53903f
C6425 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 1.11457f
C6426 m3_36652_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.53746f
C6427 m3_45124_45098# VDDR 0.0103f
C6428 VDDR sar10b_0.SWP[1] 3.51824f
C6429 sar10b_0.net16 a_62037_61731# 0.23934f
C6430 a_61400_52964# a_61677_52854# 0.09983f
C6431 a_60693_57975# VSSD 0.15009f
C6432 a_62409_59007# a_62527_58306# 0.01379f
C6433 sar10b_0.SWN[2] EN 0.15071f
C6434 VDDD a_63285_60399# 0.29934f
C6435 a_64609_64923# sar10b_0.net41 0.01215f
C6436 VSSR c1_14392_97972# 0.05555f
C6437 a_55121_59650# a_55282_59893# 0.19021f
C6438 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A 0.41861f
C6439 sar10b_0.net16 a_65333_66248# 0.15322f
C6440 sar10b_0.clk_div_0.COUNT\[1\] a_68276_50645# 0.0597f
C6441 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_7000_21578# 0.03017f
C6442 m3_15472_21578# th_dif_sw_0.VCN 0.01078f
C6443 th_dif_sw_0.CKB sar10b_0.CF[0] 0.17775f
C6444 c1_4508_21618# VCM 0.01358f
C6445 c1_45456_47378# m3_45124_47338# 1.74381f
C6446 c1_n1140_46258# m3_n1472_47338# 0.01078f
C6447 c1_n1140_47378# m3_n1472_46218# 0.01078f
C6448 a_64492_67433# a_64888_67630# 0.07682f
C6449 a_63804_67580# a_63663_67678# 0.35501f
C6450 sar10b_0.SWP[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 0.35053f
C6451 a_62527_58306# sar10b_0.net4 0.01139f
C6452 a_61395_63280# a_61086_63306# 0.07766f
C6453 m3_45124_85612# VDDR 0.01034f
C6454 m3_45124_82252# th_dif_sw_0.VCP 0.17339f
C6455 sar10b_0.net38 a_61557_57735# 0.02034f
C6456 sar10b_0._17_ sar10b_0._10_ 0.16138f
C6457 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A 0.74806f
C6458 a_61395_65944# a_61400_66284# 0.43707f
C6459 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP a_14655_5788# 0.09439f
C6460 VCM cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 3.63691f
C6461 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VDDR 2.59252f
C6462 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.39559f
C6463 c1_45456_94612# VDDR 0.01153f
C6464 a_67372_52833# a_67843_52961# 0.01114f
C6465 sar10b_0._14_ a_67419_52937# 0.016f
C6466 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A 0.04073f
C6467 a_62409_59007# a_62133_59067# 0.1263f
C6468 c1_34160_97972# VCM 0.01358f
C6469 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN sar10b_0.SWP[9] 0.18289f
C6470 sar10b_0.net2 a_65001_68627# 0.01132f
C6471 sar10b_0.net7 tdc_0.OUTN 0.19544f
C6472 m3_n1472_68812# c1_n1140_68852# 1.74381f
C6473 m3_45124_68812# c1_45456_69972# 0.01078f
C6474 m3_45124_69932# c1_45456_68852# 0.01078f
C6475 VSSR c1_45456_71092# 0.0935f
C6476 sar10b_0.clknet_1_1__leaf_CLK VSSD 1.64433f
C6477 a_63339_71265# VSSD 0.34625f
C6478 a_9853_5788# sar10b_0.SWN[7] 0.33169f
C6479 a_65573_52937# a_65861_51977# 0.05123f
C6480 m3_15472_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.2724f
C6481 c1_38396_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C6482 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.10847f
C6483 a_62133_59067# sar10b_0.net4 0.01335f
C6484 m3_28180_97932# m3_29592_97932# 0.23959f
C6485 a_60969_51311# a_61493_51596# 0.05022f
C6486 a_60747_69559# sar10b_0.net14 0.24795f
C6487 a_61493_67580# a_61358_67678# 0.35559f
C6488 c1_45456_86772# c1_45456_85652# 0.13255f
C6489 a_62181_67424# a_62527_67630# 0.07649f
C6490 c1_15804_21618# m3_15472_21578# 1.74381f
C6491 VDDR cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 6.76174f
C6492 m3_n1472_46218# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C6493 sar10b_0.net16 a_62837_61451# 0.14649f
C6494 VDDR th_dif_sw_0.CK 0.22777f
C6495 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VDDR 0.83958f
C6496 sar10b_0.net14 sar10b_0.net4 0.25303f
C6497 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C6498 m3_18296_97932# c1_17216_97972# 0.15596f
C6499 VSSD a_60747_56239# 0.34939f
C6500 VSSR m3_n1472_36138# 0.66371f
C6501 sar10b_0.net33 a_65577_51311# 0.06682f
C6502 c1_45456_51858# VDDR 0.01151f
C6503 m3_45124_55178# th_dif_sw_0.VCN 0.17339f
C6504 VSSA tdc_0.phase_detector_0.INP 1.12728f
C6505 a_n8277_54249# th_dif_sw_0.CKB 0.10346f
C6506 a_67297_55975# VSSD 0.8559f
C6507 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 0.24771f
C6508 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.53307f
C6509 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.38733f
C6510 VSSR c1_32748_21618# 0.06914f
C6511 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN 0.01132f
C6512 VSSR m3_n1472_76652# 0.66316f
C6513 VDDD a_61182_52404# 0.31789f
C6514 VSSA tdc_0.phase_detector_0.pd_out_0.A 2.14893f
C6515 c1_n1140_50738# c1_n1140_49618# 0.13255f
C6516 sar10b_0.net7 a_60747_52617# 0.02591f
C6517 sar10b_0.net34 a_66633_56639# 0.02327f
C6518 a_62709_63063# sar10b_0.net16 0.19785f
C6519 a_61737_56343# a_62949_56296# 0.07766f
C6520 a_62126_56024# a_62261_56123# 0.35559f
C6521 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VCM 0.12068f
C6522 m3_n1472_28298# VCM 0.01415f
C6523 VDDD a_62793_57675# 0.36014f
C6524 c1_n1140_78932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C6525 m3_n1472_51818# m3_n1472_50698# 0.29566f
C6526 sar10b_0._01_ a_65586_50645# 0.09184f
C6527 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 2.81343f
C6528 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C6529 w_n9655_56533# th_dif_sw_0.CKB 0.03685f
C6530 VDDD sar10b_0._04_ 1.71576f
C6531 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 1.75141f
C6532 a_68562_49747# sar10b_0.SWN[9] 0.14194f
C6533 sar10b_0.net16 sar10b_0.net11 1.04631f
C6534 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VSSR 3.13728f
C6535 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A 0.03041f
C6536 a_65682_51977# a_66109_51982# 0.04602f
C6537 sar10b_0.net3 sar10b_0.net37 0.35384f
C6538 a_17274_111642# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01076f
C6539 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.02632f
C6540 th_dif_sw_0.CKB VSSA 4.21414f
C6541 a_68073_56343# a_68325_56296# 0.27388f
C6542 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A 0.26364f
C6543 a_10731_5779# VSSR 1.11603f
C6544 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VCM 2.04844f
C6545 m3_n1472_57418# VDDR 0.02681f
C6546 m3_n1472_68812# VCM 0.01412f
C6547 a_64521_60339# a_65119_59984# 0.06623f
C6548 VDDD a_68767_65312# 0.21423f
C6549 a_64761_51028# VSSD 0.01332f
C6550 sar10b_0.net33 a_65673_56639# 0.01071f
C6551 VSSD DATA[7] 0.61149f
C6552 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSSR 1.11457f
C6553 a_63573_63303# a_64033_63591# 0.26257f
C6554 a_66197_56924# a_66633_56639# 0.16939f
C6555 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A 0.26364f
C6556 c1_n1140_52978# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C6557 a_65821_53072# VSSD 0.0151f
C6558 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A 0.02842f
C6559 a_62798_58688# sar10b_0.net39 0.05905f
C6560 VSSD a_68479_61316# 0.26072f
C6561 c1_32748_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.01078f
C6562 a_66049_69295# sar10b_0.net16 0.10408f
C6563 VSSR cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 18.4213f
C6564 VDDD a_68946_65963# 0.28035f
C6565 sar10b_0._04_ sar10b_0._08_ 0.37263f
C6566 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.04073f
C6567 sar10b_0.net33 a_66027_53575# 0.03168f
C6568 VSSR c1_n1140_42898# 0.04956f
C6569 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y sar10b_0.CF[7] 0.12541f
C6570 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A 1.33794f
C6571 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04073f
C6572 VDDD a_65643_71265# 0.25648f
C6573 a_67733_58787# VSSD 0.10006f
C6574 m3_45124_85612# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C6575 a_65957_50273# a_66762_50329# 0.29207f
C6576 tdc_0.RDY VSSD 0.81553f
C6577 m3_n1472_92332# m3_n1472_91212# 0.29566f
C6578 sar10b_0.CF[6] sar10b_0.SWP[1] 0.12434f
C6579 sar10b_0.CF[4] sar10b_0.SWP[3] 0.1195f
C6580 sar10b_0.CF[5] sar10b_0.SWP[2] 0.12163f
C6581 a_29061_5788# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 0.70991f
C6582 VSSR a_29061_108738# 0.06033f
C6583 sar10b_0.net32 a_64454_51311# 0.02117f
C6584 VDDA a_52417_60961# 0.37887f
C6585 m3_39476_21578# c1_39808_21618# 1.74381f
C6586 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A 0.03718f
C6587 m3_45124_22698# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.23379f
C6588 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A 0.4383f
C6589 a_61400_63620# VSSD 0.85606f
C6590 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 sar10b_0.CF[4] 0.40665f
C6591 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP a_34741_111361# 0.01488f
C6592 a_66109_51982# sar10b_0._07_ 0.01819f
C6593 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.12068f
C6594 VCM sar10b_0.CF[8] 3.50776f
C6595 a_55121_59650# tdc_0.OUTN 0.01823f
C6596 a_63273_56639# a_64485_56768# 0.07766f
C6597 a_67890_69727# VSSD 0.34173f
C6598 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.38072f
C6599 VDDR cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 12.9105f
C6600 m3_45124_96812# c1_45456_96852# 1.74381f
C6601 m3_n1472_96812# c1_n1140_95732# 0.01078f
C6602 m3_n1472_95692# c1_n1140_96852# 0.01078f
C6603 VSSR m3_22532_21578# 0.34286f
C6604 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y 0.32492f
C6605 sar10b_0._07_ a_65068_49569# 0.17376f
C6606 sar10b_0.net14 a_64725_68631# 0.09089f
C6607 a_62181_51440# VSSD 0.25195f
C6608 a_61358_67678# VSSD 0.13401f
C6609 sar10b_0.net10 sar10b_0.net4 0.0381f
C6610 sar10b_0.net3 sar10b_0.SWN[6] 0.02852f
C6611 c1_45456_55218# m3_45124_55178# 1.74381f
C6612 c1_n1140_54098# m3_n1472_55178# 0.01078f
C6613 c1_n1140_55218# m3_n1472_54058# 0.01078f
C6614 sar10b_0.net21 a_68169_59007# 0.0273f
C6615 sar10b_0.net13 sar10b_0.net4 0.02238f
C6616 VSSR a_34741_111361# 2.80455f
C6617 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A 0.60027f
C6618 sar10b_0.SWP[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A 0.01506f
C6619 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 2.60252f
C6620 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 0.40216f
C6621 a_62185_50043# sar10b_0.net1 0.2257f
C6622 a_61400_50300# a_61609_50282# 0.24088f
C6623 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.95194f
C6624 m3_16884_97932# VCM 0.13579f
C6625 a_n4470_65264# th_dif_sw_0.th_sw_1.CKB 0.01594f
C6626 a_61086_52650# sar10b_0.net16 0.18291f
C6627 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_38396_21618# 0.0106f
C6628 VDDA th_dif_sw_0.VCN 2.2775f
C6629 sar10b_0.net14 sar10b_0.net44 0.20061f
C6630 a_68421_54964# VSSD 0.27193f
C6631 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 0.02632f
C6632 VDDD a_64238_67295# 0.37774f
C6633 c1_22864_97972# th_dif_sw_0.VCP 0.13255f
C6634 tdc_0.OUTP tdc_0.OUTN 2.47168f
C6635 sar10b_0.net33 a_66101_58256# 0.01382f
C6636 VDDD sar10b_0._05_ 0.53894f
C6637 m3_42300_21578# VCM 0.15231f
C6638 m3_21120_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.45971f
C6639 sar10b_0.SWP[5] VDDA 0.24911f
C6640 a_64521_59303# sar10b_0.net1 0.06529f
C6641 m3_n1472_76652# c1_n1140_76692# 1.74381f
C6642 m3_45124_76652# c1_45456_77812# 0.01078f
C6643 m3_45124_77772# c1_45456_76692# 0.01078f
C6644 VSSR c1_45456_86772# 0.0935f
C6645 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 4.6018f
C6646 sar10b_0.net2 sar10b_0.net12 0.13451f
C6647 sar10b_0.net21 a_68946_53975# 0.24871f
C6648 sar10b_0.net18 DATA[3] 0.06978f
C6649 sar10b_0.CF[6] th_dif_sw_0.CK 0.17829f
C6650 VSSD a_67231_56974# 0.26829f
C6651 c1_n1140_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C6652 m3_8412_97932# m3_9824_97932# 0.23959f
C6653 a_64949_64916# a_64814_65014# 0.35559f
C6654 a_65637_64760# a_65983_64966# 0.07649f
C6655 c1_n1140_22738# m3_n1472_22698# 1.74381f
C6656 c1_45456_22738# m3_45124_23818# 0.01078f
C6657 c1_45456_23858# m3_45124_22698# 0.01078f
C6658 a_61677_66174# a_62185_66027# 0.19065f
C6659 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 21.8133f
C6660 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[8] 0.17717f
C6661 VDDD a_66593_50645# 0.17506f
C6662 sar10b_0.net3 sar10b_0._03_ 0.45714f
C6663 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.60057f
C6664 VSSR m3_n1472_51818# 0.66371f
C6665 VSSD a_62497_61303# 0.85871f
C6666 a_67209_68331# a_67733_68111# 0.04522f
C6667 a_66933_68391# a_67598_68012# 0.19065f
C6668 c1_45456_71092# VDDR 0.01153f
C6669 m3_7000_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C6670 a_67393_62635# sar10b_0.cyclic_flag_0.FINAL 0.02261f
C6671 m3_33828_21578# m3_35240_21578# 0.23959f
C6672 a_52417_60961# tdc_0.phase_detector_0.INP 0.10793f
C6673 a_69003_48621# VSSD 0.3314f
C6674 VSSR c1_5920_21618# 0.05923f
C6675 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.95198f
C6676 sar10b_0.cyclic_flag_0.FINAL sar10b_0.net40 0.04349f
C6677 a_63918_50969# a_64199_50761# 0.29207f
C6678 a_61833_57675# a_62017_57307# 0.44098f
C6679 sar10b_0.CF[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.26269f
C6680 a_66666_49313# sar10b_0.SWN[6] 0.02696f
C6681 sar10b_0._10_ sar10b_0._07_ 0.3122f
C6682 VSSR m3_n1472_92332# 0.66316f
C6683 sar10b_0.net4 a_62997_67299# 0.05102f
C6684 a_64814_65014# VSSD 0.14209f
C6685 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 sar10b_0.CF[8] 0.40665f
C6686 VSSD DATA[4] 0.70792f
C6687 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[0] 0.17732f
C6688 sar10b_0.SWP[0] sar10b_0.CF[7] 0.1469f
C6689 m3_n1472_36138# VDDR 0.02681f
C6690 a_66213_68756# sar10b_0.net16 0.24155f
C6691 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 1.30896f
C6692 a_65394_52643# a_66080_53027# 0.27693f
C6693 m3_n1472_43978# VCM 0.01415f
C6694 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSSR 1.11631f
C6695 VSSR c1_35572_97972# 0.05923f
C6696 sar10b_0.net28 sar10b_0.SWN[2] 0.05742f
C6697 VSSD sar10b_0.SWP[3] 0.96963f
C6698 sar10b_0._04_ sar10b_0._15_ 0.11741f
C6699 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 2.37549f
C6700 sar10b_0.net32 a_64188_51135# 0.03153f
C6701 sar10b_0.clknet_0_CLK a_66785_50875# 0.01395f
C6702 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_11236_21578# 0.0162f
C6703 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_28180_21578# 0.03017f
C6704 a_62185_63363# sar10b_0.net10 0.16858f
C6705 VDDD sar10b_0.CF[1] 0.46222f
C6706 m3_n1472_76652# VDDR 0.02674f
C6707 m3_n1472_84492# VCM 0.01412f
C6708 VDDD a_61677_62178# 0.27179f
C6709 m3_15472_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.59803f
C6710 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.43131f
C6711 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.14341f
C6712 a_61705_51992# VSSD 0.09782f
C6713 a_64725_68631# sar10b_0.net13 0.05536f
C6714 c1_45456_27218# c1_45456_26098# 0.13255f
C6715 a_62277_50968# sar10b_0.net1 0.01196f
C6716 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 2.47682f
C6717 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP a_38665_107026# 0.21556f
C6718 a_63967_58652# VSSD 0.28625f
C6719 a_67393_65299# a_67598_65348# 0.09983f
C6720 sar10b_0.net42 a_66645_61731# 0.17078f
C6721 a_61035_71265# sar10b_0.SWP[1] 0.1428f
C6722 m3_45124_28298# m3_45124_27178# 0.29566f
C6723 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VDDR 3.03843f
C6724 VSSR c1_n1140_62132# 0.08469f
C6725 a_68421_64288# VSSD 0.27173f
C6726 VDDD DATA[9] 0.33948f
C6727 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] a_20335_5779# 0.56899f
C6728 a_65589_69723# VSSD 0.15761f
C6729 sar10b_0.net38 sar10b_0.cyclic_flag_0.FINAL 0.18537f
C6730 m3_36652_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.53746f
C6731 m3_12648_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.53746f
C6732 th_dif_sw_0.CKB th_dif_sw_0.VCN 17.2595f
C6733 m3_19708_21578# c1_20040_21618# 1.74381f
C6734 m3_45124_38378# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C6735 a_65865_57675# a_65673_56639# 0.22273f
C6736 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VDDR 0.95194f
C6737 m3_22532_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.07708f
C6738 sar10b_0.cyclic_flag_0.FINAL a_66933_55071# 0.041f
C6739 a_60969_56639# a_62181_56768# 0.07766f
C6740 a_61153_56931# a_61493_56924# 0.24088f
C6741 m3_28180_97932# c1_28512_97972# 1.74381f
C6742 VSSR m3_45124_28298# 0.63261f
C6743 sar10b_0.net3 sar10b_0.net25 0.06225f
C6744 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] VDDR 2.16043f
C6745 sar10b_0.SWN[0] VCM 0.13077f
C6746 sar10b_0.SWP[3] sar10b_0.CF[8] 0.12688f
C6747 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y 0.07183f
C6748 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 sar10b_0.CF[8] 0.26243f
C6749 CLK a_51345_58977# 0.32697f
C6750 sar10b_0.CF[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 0.40665f
C6751 a_67209_63003# a_68169_63003# 0.03471f
C6752 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VDDR 0.75888f
C6753 a_67393_62635# a_67598_62684# 0.09983f
C6754 sar10b_0.net2 sar10b_0.net41 1.78956f
C6755 a_68562_71291# a_68235_71265# 0.08997f
C6756 sar10b_0.net46 sar10b_0.net44 1.15473f
C6757 sar10b_0.net4 a_61395_61948# 0.21842f
C6758 VDDR a_29061_108738# 5.61521f
C6759 VDDD a_61589_53459# 0.20895f
C6760 sar10b_0.net27 VSSD 0.51132f
C6761 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN 0.12375f
C6762 sar10b_0.net18 a_68946_52411# 0.03028f
C6763 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A VDDR 0.38427f
C6764 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_11568_21618# 0.0106f
C6765 m3_45124_68812# m3_45124_67692# 0.29566f
C6766 VSSR m3_45124_68812# 0.63305f
C6767 sar10b_0.net10 a_63273_61671# 0.0299f
C6768 VDDA a_n9133_63315# 0.48884f
C6769 a_69003_71265# sar10b_0.net46 0.29844f
C6770 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y VDDR 0.31983f
C6771 a_61395_52624# VSSD 0.48568f
C6772 sar10b_0.net2 a_61737_56343# 0.06927f
C6773 a_60690_54641# a_60690_53975# 0.01036f
C6774 m3_2764_21578# VCM 0.15231f
C6775 a_61035_71265# th_dif_sw_0.CK 0.15613f
C6776 VDDD a_66825_57675# 0.40103f
C6777 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] sar10b_0.SWP[1] 0.23548f
C6778 m3_n1472_84492# c1_n1140_84532# 1.74381f
C6779 m3_45124_84492# c1_45456_85652# 0.01078f
C6780 m3_45124_85612# c1_45456_84532# 0.01078f
C6781 a_61035_48621# sar10b_0.SWN[1] 0.15514f
C6782 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP 0.02666f
C6783 VDDD a_61803_48621# 0.22405f
C6784 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN 4.11482f
C6785 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A 0.41861f
C6786 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN sar10b_0.SWP[2] 0.23318f
C6787 sar10b_0.net4 a_61677_52854# 0.03455f
C6788 c1_45456_30578# m3_45124_31658# 0.01078f
C6789 c1_45456_31698# m3_45124_30538# 0.01078f
C6790 c1_n1140_30578# m3_n1472_30538# 1.74381f
C6791 VSSA tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A 0.57249f
C6792 m3_9824_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 0.0122f
C6793 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN 0.01239f
C6794 a_66153_48647# VSSD 2.27819f
C6795 sar10b_0.SWN[3] a_29061_5788# 0.75451f
C6796 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A 0.68875f
C6797 a_68421_66952# a_68767_66644# 0.07649f
C6798 a_61041_52340# a_61705_51992# 0.16939f
C6799 VDDD a_61589_50795# 0.20863f
C6800 sar10b_0.net10 a_63374_62684# 0.02124f
C6801 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN 0.02638f
C6802 a_61773_52237# VSSD 0.13186f
C6803 c1_45456_86772# VDDR 0.01153f
C6804 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 2.76083f
C6805 a_66921_61671# a_67310_61352# 0.05462f
C6806 a_66645_61731# a_67105_61303# 0.26257f
C6807 m3_14060_21578# m3_15472_21578# 0.23959f
C6808 sar10b_0.net38 a_61493_56924# 0.01297f
C6809 VSSR c1_45456_35058# 0.09348f
C6810 a_65397_56643# a_66062_57022# 0.19065f
C6811 VSSD a_60747_65937# 0.26067f
C6812 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A 0.68875f
C6813 VDDD sar10b_0._08_ 0.96396f
C6814 a_65385_64631# sar10b_0.net43 0.02718f
C6815 m3_n1472_76652# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C6816 VSSR m3_18296_97932# 0.39907f
C6817 c1_n1140_69972# c1_n1140_68852# 0.13255f
C6818 sar10b_0._01_ a_65577_51311# 0.06407f
C6819 sar10b_0._10_ a_65394_52643# 0.02781f
C6820 m3_18296_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.25796f
C6821 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C6822 m3_n1472_51818# VDDR 0.02681f
C6823 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 0.38722f
C6824 a_63273_61671# a_63525_61624# 0.27388f
C6825 sar10b_0.CF[0] sar10b_0.CF[3] 0.11787f
C6826 sar10b_0.CF[1] sar10b_0.CF[2] 44.0085f
C6827 VSSR m3_43712_21578# 0.54637f
C6828 a_65185_68919# VSSD 0.81827f
C6829 sar10b_0.net45 sar10b_0.SWP[7] 0.11955f
C6830 a_66933_63063# sar10b_0.net3 0.2327f
C6831 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 0.02638f
C6832 VDDD a_68767_67976# 0.21501f
C6833 m3_45124_22698# th_dif_sw_0.VCN 0.16468f
C6834 VSSA a_n4470_65264# 2.16169f
C6835 a_65957_50273# VSSD 0.53191f
C6836 VDDD DATA[6] 0.41818f
C6837 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A 0.07183f
C6838 a_64339_51661# a_64454_51311# 0.22516f
C6839 a_67209_64335# sar10b_0.cyclic_flag_0.FINAL 0.24121f
C6840 sar10b_0.net14 sar10b_0.cyclic_flag_0.FINAL 0.14652f
C6841 a_63273_67295# a_62997_67299# 0.12579f
C6842 sar10b_0.net33 a_66255_50749# 0.01101f
C6843 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A 0.05472f
C6844 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.38733f
C6845 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 2.47087f
C6846 m3_n1472_92332# VDDR 0.02674f
C6847 VDDD a_67445_60119# 0.21629f
C6848 sar10b_0.SWP[8] a_5929_113881# 0.17051f
C6849 m3_38064_97932# VCM 0.15231f
C6850 sar10b_0.net10 a_60747_61941# 0.27587f
C6851 a_64910_59686# VSSD 0.12961f
C6852 c1_45456_35058# c1_45456_33938# 0.13255f
C6853 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VDDR 0.95259f
C6854 c1_44044_97972# th_dif_sw_0.VCP 0.13255f
C6855 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.44217f
C6856 sar10b_0.net28 sar10b_0.net1 0.56463f
C6857 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 0.40665f
C6858 c1_15804_97972# VCM 0.01358f
C6859 m3_42300_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C6860 VDDA a_n9133_57045# 0.48884f
C6861 m3_45124_36138# m3_45124_35018# 0.29566f
C6862 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 1.71649f
C6863 VSSR c1_n1140_77812# 0.04956f
C6864 a_68562_71291# VSSD 0.29379f
C6865 VSSD sar10b_0.net22 0.93976f
C6866 a_64454_51311# CLK 0.01921f
C6867 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] a_10731_113461# 0.3365f
C6868 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A 1.11457f
C6869 c1_20040_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C6870 sar10b_0.clknet_0_CLK sar10b_0.clknet_1_1__leaf_CLK 0.01122f
C6871 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 0.24774f
C6872 c1_5920_21618# m3_7000_21578# 0.15596f
C6873 m3_45124_54058# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C6874 a_5051_5788# sar10b_0.SWN[8] 0.22599f
C6875 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.41861f
C6876 a_64521_59303# a_65481_59303# 0.03432f
C6877 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR 0.95166f
C6878 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN 3.31932f
C6879 m3_8412_97932# c1_8744_97972# 1.74381f
C6880 VSSR m3_45124_43978# 0.63261f
C6881 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VSSR 1.33727f
C6882 a_62025_53679# sar10b_0.net6 0.01814f
C6883 sar10b_0.SWP[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.33822f
C6884 a_61182_52404# a_61496_52091# 0.07826f
C6885 sar10b_0.SWP[1] sar10b_0.CF[7] 0.13044f
C6886 c1_1684_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26825f
C6887 sar10b_0.SWP[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A 0.01506f
C6888 m3_28180_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C6889 a_62985_63003# a_64197_62956# 0.07766f
C6890 a_63374_62684# a_63509_62783# 0.35559f
C6891 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 6.79685f
C6892 sar10b_0.net34 a_65573_52937# 0.01473f
C6893 sar10b_0.net3 sar10b_0._13_ 0.22626f
C6894 a_62793_57675# a_63391_57320# 0.06623f
C6895 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[1] 0.01887f
C6896 m3_45124_76652# m3_45124_75532# 0.29566f
C6897 a_64199_50761# a_64428_50947# 0.18757f
C6898 a_64521_60339# sar10b_0.net12 0.02517f
C6899 a_62181_58100# sar10b_0.net16 0.16986f
C6900 VSSR m3_45124_84492# 0.63305f
C6901 sar10b_0.net38 a_65397_56643# 0.06828f
C6902 VDDD a_68133_61624# 0.27603f
C6903 m3_45124_28298# VDDR 0.0103f
C6904 VDDD sar10b_0.CF[2] 0.41245f
C6905 a_65577_51311# sar10b_0.net35 0.04658f
C6906 m3_45124_92332# c1_45456_93492# 0.01078f
C6907 m3_n1472_92332# c1_n1140_92372# 1.74381f
C6908 m3_45124_93452# c1_45456_92372# 0.01078f
C6909 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP 3.13167f
C6910 sar10b_0.clk_div_0.COUNT\[3\] sar10b_0.net37 0.04961f
C6911 a_67209_63003# VSSD 0.55646f
C6912 VSSA sar10b_0.CF[3] 0.90846f
C6913 VDDD a_67598_58688# 0.27431f
C6914 a_62025_51015# sar10b_0.net6 0.01187f
C6915 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_32416_21578# 0.0162f
C6916 sar10b_0.net32 a_64356_51029# 0.0167f
C6917 VDDD sar10b_0._15_ 0.2348f
C6918 c1_34160_21618# VCM 0.01358f
C6919 c1_n1140_38418# m3_n1472_38378# 1.74381f
C6920 c1_45456_38418# m3_45124_39498# 0.01078f
C6921 VDDD a_61086_63306# 0.31749f
C6922 c1_45456_39538# m3_45124_38378# 0.01078f
C6923 a_67113_56343# a_67637_56123# 0.04522f
C6924 a_66837_56403# a_67502_56024# 0.19065f
C6925 VDDA sar10b_0.SWP[6] 0.24919f
C6926 m3_45124_68812# VDDR 0.01034f
C6927 m3_45124_65452# th_dif_sw_0.VCP 0.17339f
C6928 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_36482_8700# 0.01076f
C6929 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP 0.02666f
C6930 sar10b_0.CF[7] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 0.01386f
C6931 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C6932 VSSD a_67733_66779# 0.09755f
C6933 th_dif_sw_0.CK sar10b_0.CF[7] 0.17893f
C6934 VDDD a_61493_51596# 0.20732f
C6935 a_61929_57971# sar10b_0.net8 0.01111f
C6936 VDDD a_62527_67630# 0.20174f
C6937 sar10b_0.net40 a_61395_60616# 0.01513f
C6938 sar10b_0.net13 sar10b_0.cyclic_flag_0.FINAL 0.02792f
C6939 VSSD a_65966_58354# 0.13412f
C6940 c1_14392_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.26836f
C6941 sar10b_0.CF[6] tdc_0.OUTP 0.16093f
C6942 a_62985_63003# sar10b_0.net2 0.01879f
C6943 VDDD a_64809_65963# 0.86421f
C6944 sar10b_0.clk_div_0.COUNT\[2\] a_68331_52243# 0.03312f
C6945 a_14655_5788# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 0.3928f
C6946 a_60693_67299# sar10b_0.net16 0.22905f
C6947 m3_n1472_57418# c1_n1140_56338# 0.01078f
C6948 VSSR c1_45456_50738# 0.09348f
C6949 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y 0.07183f
C6950 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] th_dif_sw_0.VCN 4.58977f
C6951 a_61358_58354# sar10b_0.net38 0.02848f
C6952 sar10b_0._08_ sar10b_0._15_ 0.05089f
C6953 VDDD a_68169_55011# 0.36731f
C6954 m3_n1472_92332# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C6955 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] a_29939_111781# 0.80139f
C6956 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VCM 3.3783f
C6957 c1_n1140_77812# c1_n1140_76692# 0.13255f
C6958 sar10b_0.net16 a_61921_55975# 0.09742f
C6959 VINP th_dif_sw_0.th_sw_1.CKB 0.08416f
C6960 m3_31004_21578# c1_29924_21618# 0.15596f
C6961 m3_n1472_29418# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C6962 sar10b_0.SWN[8] VCM 0.13075f
C6963 a_64188_51135# CLK 0.01407f
C6964 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C6965 sar10b_0.CF[5] sar10b_0.SWN[3] 0.12071f
C6966 c1_35572_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26825f
C6967 a_66389_69443# a_66825_69663# 0.16939f
C6968 m3_39476_97932# c1_38396_97972# 0.15596f
C6969 VSSR m3_4176_21578# 0.54637f
C6970 a_62409_59007# sar10b_0.net8 0.01926f
C6971 sar10b_0.net6 a_61461_56403# 0.04357f
C6972 sar10b_0.net46 sar10b_0.cyclic_flag_0.FINAL 0.03151f
C6973 VDDD a_65119_59984# 0.19838f
C6974 sar10b_0._12_ a_67439_50041# 0.1709f
C6975 VDDD a_66633_56639# 0.37013f
C6976 c1_45456_35058# VDDR 0.01151f
C6977 sar10b_0.CF[1] tdc_0.OUTN 0.14506f
C6978 m3_45124_38378# th_dif_sw_0.VCN 0.17339f
C6979 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A 0.68875f
C6980 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C6981 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 a_10731_113461# 0.20413f
C6982 sar10b_0.net3 a_65682_49313# 0.15872f
C6983 a_64245_59307# VSSD 0.1667f
C6984 a_68331_52243# VSSD 0.30889f
C6985 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.11339f
C6986 sar10b_0.CF[5] a_60747_62899# 0.14278f
C6987 sar10b_0.SWN[2] sar10b_0.CF[9] 0.23443f
C6988 sar10b_0.net4 sar10b_0.net8 0.25575f
C6989 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] a_14655_111306# 1.18623f
C6990 m3_26768_97932# th_dif_sw_0.VCP 0.01078f
C6991 m3_23944_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 0.15657f
C6992 m3_n1472_97932# VCM 0.16643f
C6993 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 0.12357f
C6994 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_20040_21618# 0.0106f
C6995 a_60690_54641# VSSD 0.41541f
C6996 VSSR sar10b_0.CF[1] 17.4137f
C6997 a_60693_67299# a_60969_67295# 0.1263f
C6998 c1_45456_42898# c1_45456_41778# 0.13255f
C6999 sar10b_0.SWN[9] VCM 0.13075f
C7000 a_66080_53027# VSSD 0.14927f
C7001 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN sar10b_0.CF[4] 0.09303f
C7002 VDDD a_68562_48647# 0.22445f
C7003 m3_2764_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C7004 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A 0.43651f
C7005 m3_23944_21578# VCM 0.13579f
C7006 c1_n1140_62132# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C7007 m3_45124_43978# m3_45124_42858# 0.29566f
C7008 sar10b_0._10_ a_64780_52239# 0.0209f
C7009 sar10b_0.net34 sar10b_0.clk_div_0.COUNT\[0\] 0.07533f
C7010 VSSR c1_n1140_93492# 0.04956f
C7011 a_61833_57675# a_61929_56639# 0.02084f
C7012 VDDA CLK 4.80039f
C7013 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.68971f
C7014 a_67372_52243# sar10b_0.net35 0.03376f
C7015 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 2.82798f
C7016 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A sar10b_0.CF[4] 0.02149f
C7017 VDDD a_65983_64966# 0.21491f
C7018 sar10b_0.net40 a_62017_57307# 0.14471f
C7019 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.12068f
C7020 a_61400_52964# sar10b_0.net1 0.0193f
C7021 sar10b_0.net14 a_65397_56643# 0.04311f
C7022 a_64521_60339# sar10b_0.net41 0.07097f
C7023 VDDD a_65577_57971# 0.8319f
C7024 a_62025_53679# VSSD 0.28996f
C7025 a_68133_60292# sar10b_0.net3 0.18334f
C7026 a_66666_51977# a_66865_52076# 0.29821f
C7027 sar10b_0.net16 a_61833_57675# 0.21251f
C7028 sar10b_0.CF[5] VDDA 0.39815f
C7029 VDDD a_68946_49747# 0.23306f
C7030 c1_n1140_36178# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C7031 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A 0.95194f
C7032 VDDD a_61677_64842# 0.2729f
C7033 a_67881_61671# a_68479_61316# 0.06623f
C7034 sar10b_0.net38 a_63797_56924# 0.02061f
C7035 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A 0.02842f
C7036 a_24259_109594# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 0.60421f
C7037 VSSR a_39543_5779# 3.14203f
C7038 VSSR c1_n1140_26098# 0.04956f
C7039 a_62025_51015# sar10b_0.net30 0.02363f
C7040 a_63918_50969# a_64188_51135# 0.08669f
C7041 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 0.21044f
C7042 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 0.40665f
C7043 sar10b_0._01_ a_64924_52385# 0.01119f
C7044 m3_45124_68812# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C7045 a_65682_49313# a_66666_49313# 0.08669f
C7046 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 2.56917f
C7047 m3_45124_84492# m3_45124_83372# 0.29566f
C7048 VSSR m3_39476_97932# 0.54637f
C7049 sar10b_0.SWP[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 0.38458f
C7050 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 sar10b_0.SWN[8] 0.25013f
C7051 VDDD a_63621_58960# 0.27383f
C7052 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A 0.02842f
C7053 m3_39476_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.53746f
C7054 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.17717f
C7055 m3_45124_43978# VDDR 0.0103f
C7056 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VDDR 0.74952f
C7057 a_61400_52964# a_62185_52707# 0.26257f
C7058 a_61609_52946# a_61677_52854# 0.35559f
C7059 a_62409_59007# sar10b_0.net9 0.21037f
C7060 a_61153_58263# VSSD 0.85034f
C7061 VDDD a_68169_64335# 0.36668f
C7062 a_67209_59007# a_68421_58960# 0.07766f
C7063 a_67393_58639# a_67733_58787# 0.24088f
C7064 VDDD tdc_0.OUTN 0.32622f
C7065 VSSR c1_17216_97972# 0.04949f
C7066 sar10b_0.clk_div_0.COUNT\[2\] a_68276_50645# 0.01108f
C7067 VDDD a_65865_69663# 0.85773f
C7068 a_62025_51015# VSSD 0.28732f
C7069 sar10b_0.net16 a_65769_65963# 0.26571f
C7070 a_61065_53679# sar10b_0.net16 0.17797f
C7071 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.40463f
C7072 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_9824_21578# 0.03017f
C7073 m3_18296_21578# th_dif_sw_0.VCN 0.01078f
C7074 a_65068_49569# VSSD 0.15845f
C7075 a_61493_67580# sar10b_0.net39 0.02035f
C7076 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A 0.05472f
C7077 c1_7332_21618# VCM 0.01358f
C7078 a_62527_51646# sar10b_0.net6 0.01293f
C7079 c1_n1140_46258# m3_n1472_46218# 1.74381f
C7080 c1_45456_46258# m3_45124_47338# 0.01078f
C7081 c1_45456_47378# m3_45124_46218# 0.01078f
C7082 sar10b_0.net9 sar10b_0.net4 0.91592f
C7083 VDDD a_61677_60846# 0.27219f
C7084 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[9] 0.01887f
C7085 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C7086 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 a_29939_111781# 0.51724f
C7087 a_60945_63273# a_61400_63620# 0.3578f
C7088 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A 0.43773f
C7089 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C7090 m3_45124_81132# th_dif_sw_0.VCP 0.17339f
C7091 m3_45124_84492# VDDR 0.01034f
C7092 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] a_24259_5788# 1.78742f
C7093 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y sar10b_0.CF[8] 0.12541f
C7094 a_61395_65944# a_61609_66266# 0.04522f
C7095 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] a_33863_107882# 2.38822f
C7096 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A VSSR 0.43728f
C7097 CLK tdc_0.phase_detector_0.INP 0.18399f
C7098 sar10b_0.net3 sar10b_0.clknet_1_0__leaf_CLK 0.03833f
C7099 sar10b_0.net14 a_65761_58263# 0.03028f
C7100 a_10731_5779# sar10b_0.SWN[7] 0.24998f
C7101 a_62409_59007# a_62593_58639# 0.44098f
C7102 sar10b_0.net4 a_61395_64612# 0.2205f
C7103 a_53652_59132# tdc_0.phase_detector_0.pd_out_0.A 0.18921f
C7104 c1_36984_97972# VCM 0.01358f
C7105 a_68946_59303# sar10b_0.net23 0.24949f
C7106 m3_n1472_68812# c1_n1140_67732# 0.01078f
C7107 a_69003_48621# sar10b_0.SWN[8] 0.15514f
C7108 m3_45124_68812# c1_45456_68852# 1.74381f
C7109 m3_n1472_67692# c1_n1140_68852# 0.01078f
C7110 VSSR c1_45456_69972# 0.0935f
C7111 a_64705_59595# sar10b_0.net13 0.02363f
C7112 th_dif_sw_0.VCN sar10b_0.CF[3] 0.42231f
C7113 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 1.39285f
C7114 th_dif_sw_0.VCP sar10b_0.CF[9] 0.33356f
C7115 VDDA a_52417_59293# 0.37887f
C7116 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN sar10b_0.CF[8] 0.05167f
C7117 m3_18296_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.25796f
C7118 c1_41220_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C7119 a_68169_59007# sar10b_0.net3 0.27767f
C7120 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] 2.78256f
C7121 m3_29592_97932# m3_31004_97932# 0.23959f
C7122 a_60969_51311# a_61929_51311# 0.03432f
C7123 a_61153_51603# a_62181_51440# 0.07826f
C7124 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VCM 1.75387f
C7125 a_67209_64335# a_66933_64395# 0.1263f
C7126 VDDA th_dif_sw_0.th_sw_0.th_sw_main_0.VGS 0.12838f
C7127 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN 0.02638f
C7128 c1_n1140_85652# c1_n1140_84532# 0.13255f
C7129 c1_17216_21618# m3_16884_21578# 1.74381f
C7130 VDDD a_60747_52617# 0.22239f
C7131 m3_n1472_45098# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C7132 sar10b_0._07_ a_65021_50292# 0.01579f
C7133 a_67881_60339# VSSD 0.29f
C7134 VSSD a_61461_56403# 0.14658f
C7135 m3_19708_97932# c1_18628_97972# 0.15596f
C7136 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.11339f
C7137 VSSR m3_n1472_35018# 0.66371f
C7138 sar10b_0.net3 a_66933_65727# 0.23174f
C7139 sar10b_0.SWN[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.02058f
C7140 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.36778f
C7141 th_dif_sw_0.CKB CLK 0.64701f
C7142 a_63745_59971# sar10b_0.net10 0.01713f
C7143 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C7144 c1_45456_50738# VDDR 0.01151f
C7145 m3_45124_54058# th_dif_sw_0.VCN 0.17339f
C7146 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A 0.05472f
C7147 a_67637_56123# VSSD 0.09882f
C7148 sar10b_0.net3 sar10b_0.net28 0.04428f
C7149 VDDD a_65643_48621# 0.26113f
C7150 VSSR c1_35572_21618# 0.05923f
C7151 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A 0.41861f
C7152 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A 0.10815f
C7153 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45324f
C7154 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26364f
C7155 a_65589_57735# a_66049_57307# 0.26257f
C7156 a_65865_57675# a_66254_57356# 0.05462f
C7157 tdc_0.phase_detector_0.pd_out_0.B a_53564_60302# 0.47998f
C7158 VSSR m3_n1472_75532# 0.66316f
C7159 VDDD a_61496_52091# 0.22325f
C7160 sar10b_0.net33 a_65481_59303# 0.01012f
C7161 c1_45456_50738# c1_45456_49618# 0.13255f
C7162 sar10b_0._10_ VSSD 2.68867f
C7163 sar10b_0.net7 a_60945_52617# 0.017f
C7164 a_63169_62635# sar10b_0.net16 0.09427f
C7165 a_61921_55975# a_62697_56343# 0.3578f
C7166 w_n9655_63119# th_dif_sw_0.th_sw_1.CK 0.0106f
C7167 sar10b_0.SWP[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 0.44186f
C7168 VSSD a_62997_56643# 0.15488f
C7169 sar10b_0.CF[5] th_dif_sw_0.CKB 0.08579f
C7170 m3_n1472_27178# VCM 0.01415f
C7171 VDDD a_63391_57320# 0.20393f
C7172 c1_n1140_77812# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C7173 m3_45124_51818# m3_45124_50698# 0.29566f
C7174 sar10b_0.net24 VSSD 0.51858f
C7175 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 3.10203f
C7176 sar10b_0.net33 sar10b_0.net3 0.02628f
C7177 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 0.9283f
C7178 a_65861_51977# a_66368_52081# 0.21226f
C7179 a_65682_51977# a_66216_52022# 0.35097f
C7180 a_68325_56296# a_68671_55988# 0.07649f
C7181 sar10b_0.net39 a_61400_64952# 0.01673f
C7182 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y sar10b_0.CF[0] 0.12541f
C7183 VDDR sar10b_0.CF[1] 1.70782f
C7184 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A 0.10815f
C7185 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 0.20254f
C7186 c1_20040_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.01445f
C7187 sar10b_0.net10 a_60747_62899# 0.28883f
C7188 m3_n1472_67692# VCM 0.01412f
C7189 sar10b_0.net32 sar10b_0.net16 0.34427f
C7190 VDDD a_65001_68627# 0.85208f
C7191 a_63849_63299# a_64373_63584# 0.05022f
C7192 sar10b_0.clknet_0_CLK a_66153_48647# 0.4836f
C7193 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A 0.38427f
C7194 a_66885_56768# a_67231_56974# 0.07649f
C7195 sar10b_0.CF[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A 0.02149f
C7196 c1_n1140_51858# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C7197 sar10b_0.SWP[9] VDDA 0.25989f
C7198 sar10b_0.net39 VSSD 4.12029f
C7199 a_51603_58977# th_dif_sw_0.VCP 0.05272f
C7200 sar10b_0.SWN[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 0.42754f
C7201 a_66389_69443# sar10b_0.net16 0.14563f
C7202 sar10b_0._05_ a_65573_52937# 0.2767f
C7203 VSSR c1_n1140_41778# 0.04956f
C7204 VSSA VINP 8.94453f
C7205 a_60747_63273# sar10b_0.net11 0.27587f
C7206 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP sar10b_0.CF[2] 0.10522f
C7207 tdc_0.OUTN sar10b_0.CF[2] 0.17678f
C7208 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP 0.02666f
C7209 m3_45124_84492# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C7210 sar10b_0.net13 a_65761_58263# 0.0203f
C7211 m3_45124_92332# m3_45124_91212# 0.29566f
C7212 VSSR m3_n60_97932# 0.54178f
C7213 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 0.24802f
C7214 sar10b_0.net34 sar10b_0.SWN[6] 0.24707f
C7215 m3_40888_21578# c1_41220_21618# 1.74381f
C7216 VDDA a_51861_60437# 0.18641f
C7217 m3_n60_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.53633f
C7218 a_61609_63602# VSSD 0.09912f
C7219 a_66216_52022# sar10b_0._07_ 0.03801f
C7220 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 a_20335_5779# 0.36136f
C7221 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSSR 1.10672f
C7222 a_62997_56643# sar10b_0.net31 0.01513f
C7223 a_63457_56931# a_63797_56924# 0.24088f
C7224 sar10b_0.net39 a_63295_55988# 0.2715f
C7225 m3_45124_95692# c1_45456_96852# 0.01078f
C7226 m3_n1472_95692# c1_n1140_95732# 1.74381f
C7227 m3_45124_96812# c1_45456_95732# 0.01078f
C7228 VSSR m3_25356_21578# 0.44647f
C7229 VSSD a_67209_65667# 0.51418f
C7230 VSSR sar10b_0.CF[2] 18.5824f
C7231 a_51345_58977# a_51861_59345# 0.08876f
C7232 VSSD a_62037_61731# 0.13599f
C7233 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y sar10b_0.CF[9] 0.12541f
C7234 sar10b_0._04_ sar10b_0.clk_div_0.COUNT\[0\] 0.17636f
C7235 a_62527_51646# VSSD 0.25424f
C7236 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.21389f
C7237 c1_45456_54098# m3_45124_55178# 0.01078f
C7238 c1_n1140_54098# m3_n1472_54058# 1.74381f
C7239 sar10b_0.net21 a_68767_58652# 0.01441f
C7240 c1_45456_55218# m3_45124_54058# 0.01078f
C7241 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] a_34741_5779# 0.91754f
C7242 VSSD a_65333_66248# 0.10258f
C7243 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 4.10362f
C7244 a_1127_114301# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.10438f
C7245 sar10b_0.clknet_0_CLK a_65957_50273# 0.05665f
C7246 m3_45124_96812# th_dif_sw_0.VCP 0.16468f
C7247 m3_19708_97932# VCM 0.13579f
C7248 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_41220_21618# 0.0106f
C7249 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 0.94823f
C7250 th_dif_sw_0.CKB sar10b_0.net29 0.04821f
C7251 VDDD a_63663_67678# 0.27789f
C7252 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.11339f
C7253 a_66921_60339# sar10b_0.cyclic_flag_0.FINAL 0.24734f
C7254 a_61677_62178# a_62185_62031# 0.19065f
C7255 sar10b_0.net39 sar10b_0.net31 0.14337f
C7256 c1_22864_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 0.02527f
C7257 m3_45124_21578# VCM 0.15685f
C7258 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C7259 a_64491_71265# sar10b_0.net42 0.26512f
C7260 m3_23944_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C7261 m3_45124_76652# c1_45456_76692# 1.74381f
C7262 m3_n1472_75532# c1_n1140_76692# 0.01078f
C7263 sar10b_0.net34 sar10b_0._03_ 0.02569f
C7264 m3_n1472_76652# c1_n1140_75572# 0.01078f
C7265 VSSR c1_45456_85652# 0.0935f
C7266 sar10b_0.net38 a_60945_61941# 0.0238f
C7267 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A 0.28117f
C7268 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A 0.38472f
C7269 c1_1684_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C7270 m3_9824_97932# m3_11236_97932# 0.23959f
C7271 VDDD VDDR 0.29087f
C7272 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04073f
C7273 c1_n1140_93492# c1_n1140_92372# 0.13255f
C7274 c1_45456_22738# m3_45124_22698# 1.74381f
C7275 sar10b_0.net40 a_66049_57307# 0.15223f
C7276 c1_n1140_21618# m3_n1472_22698# 0.01078f
C7277 c1_n1140_22738# m3_n1472_21578# 0.01078f
C7278 tdc_0.OUTP sar10b_0.CF[7] 0.16093f
C7279 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A VDDR 0.38397f
C7280 sar10b_0.net21 sar10b_0.net18 0.01003f
C7281 th_dif_sw_0.th_sw_1.CK a_n8277_65767# 0.10085f
C7282 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A 0.39656f
C7283 m3_n60_97932# c1_n1140_97972# 0.15596f
C7284 VSSR m3_n1472_50698# 0.66371f
C7285 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A 0.04562f
C7286 VSSD a_62837_61451# 0.10385f
C7287 a_67393_67963# a_67598_68012# 0.09983f
C7288 sar10b_0.net16 a_65589_57735# 0.23596f
C7289 c1_45456_69972# VDDR 0.01153f
C7290 m3_9824_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C7291 VSSR m3_45124_57418# 0.6971f
C7292 sar10b_0.net17 a_61803_48621# 0.10448f
C7293 m3_35240_21578# m3_36652_21578# 0.23959f
C7294 VSSR c1_8744_21618# 0.054f
C7295 VDDD sar10b_0.net17 1.54571f
C7296 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 0.84046f
C7297 a_64188_51135# a_64428_50947# 0.35097f
C7298 a_63918_50969# a_64356_51029# 0.02614f
C7299 a_61557_57735# a_62222_57356# 0.19065f
C7300 a_61833_57675# a_62357_57455# 0.04522f
C7301 sar10b_0.CF[1] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.01368f
C7302 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.41774f
C7303 a_67371_49579# sar10b_0.SWN[6] 0.14195f
C7304 VDDD a_67598_66680# 0.2745f
C7305 a_63849_63299# sar10b_0.net16 0.1871f
C7306 VSSR m3_n1472_91212# 0.66316f
C7307 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A 0.02149f
C7308 VDDD sar10b_0.SWP[7] 2.63086f
C7309 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04073f
C7310 m3_n1472_35018# VDDR 0.02681f
C7311 a_66559_68962# sar10b_0.net16 0.06061f
C7312 a_65394_52643# a_66577_52883# 0.0649f
C7313 m3_n1472_42858# VCM 0.01546f
C7314 c1_n1140_93492# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C7315 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.59327f
C7316 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A sar10b_0.CF[0] 0.26303f
C7317 VSSR c1_38396_97972# 0.05923f
C7318 a_62709_63063# VSSD 0.13658f
C7319 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C7320 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN 0.74816f
C7321 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A sar10b_0.CF[7] 0.02149f
C7322 sar10b_0.cyclic_flag_0.FINAL a_67105_61303# 0.03441f
C7323 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_14060_21578# 0.0162f
C7324 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_31004_21578# 0.03017f
C7325 sar10b_0.CF[6] sar10b_0.CF[1] 0.1132f
C7326 sar10b_0._08_ sar10b_0.net17 0.12485f
C7327 sar10b_0.CF[1] sar10b_0.SWN[1] 2.74531f
C7328 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP sar10b_0.CF[8] 0.10502f
C7329 VDDD a_61677_50190# 0.27267f
C7330 VSSD sar10b_0.net11 2.28524f
C7331 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A 0.68875f
C7332 m3_n1472_75532# VDDR 0.02674f
C7333 sar10b_0.SWP[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A 0.01506f
C7334 m3_n1472_83372# VCM 0.01412f
C7335 VDDD a_62185_62031# 0.30442f
C7336 m3_18296_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.18044f
C7337 a_61929_57971# sar10b_0.net1 0.01745f
C7338 sar10b_0.clk_div_0.COUNT\[0\] a_66593_50645# 0.02636f
C7339 c1_n1140_26098# c1_n1140_24978# 0.13255f
C7340 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C7341 a_43467_106170# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 1.02702f
C7342 VDDD sar10b_0.net12 2.78966f
C7343 a_63369_59007# a_63967_58652# 0.06623f
C7344 sar10b_0.SWP[5] sar10b_0.SWP[4] 14.3376f
C7345 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 2.64269f
C7346 VSSR a_5051_113018# 0.06023f
C7347 a_67209_65667# a_68421_65620# 0.07766f
C7348 a_67598_65348# a_67733_65447# 0.35559f
C7349 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSSR 1.11457f
C7350 m3_n1472_27178# m3_n1472_26058# 0.29566f
C7351 VSSR c1_n1140_57458# 0.08618f
C7352 a_66049_69295# VSSD 0.85713f
C7353 m3_39476_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.53746f
C7354 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 sar10b_0.SWN[0] 0.48484f
C7355 m3_15472_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.59803f
C7356 sar10b_0.net16 a_66062_57022# 0.23979f
C7357 sar10b_0.net34 a_66464_50363# 0.02007f
C7358 m3_45124_22698# c1_45456_21618# 0.01078f
C7359 m3_21120_21578# c1_21452_21618# 1.74381f
C7360 m3_45124_37258# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C7361 a_61249_53311# a_62277_53632# 0.07826f
C7362 VDDD a_65573_52937# 0.84433f
C7363 m3_25356_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.57708f
C7364 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A 0.10815f
C7365 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] 17.3154f
C7366 a_61065_51015# CLK 0.01609f
C7367 a_61153_56931# a_61929_56639# 0.3578f
C7368 sar10b_0.net33 a_65861_51977# 0.02629f
C7369 sar10b_0._04_ sar10b_0.net37 0.02883f
C7370 m3_29592_97932# c1_29924_97972# 1.74381f
C7371 a_66153_48647# a_68235_48621# 0.01142f
C7372 VSSR m3_45124_27178# 0.63261f
C7373 sar10b_0.SWN[1] a_39543_5779# 0.71842f
C7374 a_61395_49960# sar10b_0.net1 0.07276f
C7375 a_60747_49953# a_60945_49953# 0.06623f
C7376 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP 5.56695f
C7377 VDDD a_63662_57022# 0.24917f
C7378 sar10b_0.net21 sar10b_0.net23 0.13134f
C7379 a_67209_66999# a_68169_66999# 0.03471f
C7380 CLK tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A 0.09504f
C7381 sar10b_0.net4 sar10b_0.net1 0.67875f
C7382 sar10b_0.SWN[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.4706f
C7383 sar10b_0.net3 a_66961_50219# 0.01933f
C7384 a_67598_62684# a_67733_62783# 0.35559f
C7385 a_66825_57675# a_67423_57320# 0.06623f
C7386 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_14392_21618# 0.0106f
C7387 sar10b_0.net16 a_61153_56931# 0.12281f
C7388 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A 0.10815f
C7389 a_67564_50907# sar10b_0._12_ 0.14435f
C7390 sar10b_0.net1 a_62126_56024# 0.01048f
C7391 m3_n1472_67692# m3_n1472_66572# 0.29566f
C7392 VSSR m3_45124_67692# 0.63305f
C7393 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VDDR 0.95741f
C7394 sar10b_0.net4 a_61400_66284# 0.01899f
C7395 VDDD DATA[0] 0.13104f
C7396 VDDR sar10b_0.CF[2] 1.70405f
C7397 a_61086_52650# VSSD 0.26848f
C7398 sar10b_0.net32 a_64233_56639# 0.02693f
C7399 sar10b_0.net16 sar10b_0.net40 0.79298f
C7400 m3_5588_21578# VCM 0.15231f
C7401 VDDD a_67423_57320# 0.23415f
C7402 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A 0.04073f
C7403 m3_n1472_83372# c1_n1140_84532# 0.01078f
C7404 m3_n1472_84492# c1_n1140_83412# 0.01078f
C7405 m3_45124_84492# c1_45456_84532# 1.74381f
C7406 sar10b_0.net47 sar10b_0.net27 0.01096f
C7407 sar10b_0.CF[6] VDDD 0.35261f
C7408 VDDD sar10b_0.SWN[1] 0.20156f
C7409 sar10b_0.net4 a_62185_52707# 0.04081f
C7410 sar10b_0.net3 a_66933_68391# 0.22293f
C7411 c1_n1140_29458# m3_n1472_30538# 0.01078f
C7412 c1_n1140_30578# m3_n1472_29418# 0.01078f
C7413 c1_45456_30578# m3_45124_30538# 1.74381f
C7414 VDDD a_60969_57971# 0.9044f
C7415 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 sar10b_0.SWP[9] 0.35379f
C7416 a_61491_52222# a_61705_51992# 0.05022f
C7417 a_249_5788# sar10b_0.SWN[9] 0.11779f
C7418 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP 1.46154f
C7419 VDDD a_60690_49683# 0.96667f
C7420 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN 0.02638f
C7421 c1_45456_85652# VDDR 0.01153f
C7422 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A 0.42509f
C7423 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.42509f
C7424 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[8] 0.05939f
C7425 sar10b_0.clk_div_0.COUNT\[1\] a_67439_50041# 0.08089f
C7426 m3_15472_21578# m3_16884_21578# 0.23959f
C7427 sar10b_0.net38 a_61929_56639# 0.05481f
C7428 a_64338_52411# sar10b_0._01_ 0.14194f
C7429 VSSR c1_45456_33938# 0.09348f
C7430 a_61249_50647# a_62277_50968# 0.07826f
C7431 a_64339_51661# sar10b_0.net16 0.06677f
C7432 sar10b_0._16_ a_67372_52833# 0.14642f
C7433 sar10b_0.CF[4] sar10b_0.SWN[4] 2.40078f
C7434 m3_n1472_75532# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C7435 sar10b_0.SWP[8] VSSD 0.74066f
C7436 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A 0.6007f
C7437 VSSR m3_21120_97932# 0.34859f
C7438 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 0.20739f
C7439 c1_45456_69972# c1_45456_68852# 0.13255f
C7440 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C7441 m3_21120_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.21656f
C7442 a_44345_5779# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 1.14986f
C7443 m3_n1472_50698# VDDR 0.02681f
C7444 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN sar10b_0.CF[0] 0.12404f
C7445 a_63525_61624# a_63871_61316# 0.07649f
C7446 VDDD a_67611_50645# 0.18977f
C7447 VSSR c1_n1140_97972# 0.07152f
C7448 VDDD sar10b_0.net41 2.35898f
C7449 sar10b_0.net38 sar10b_0.net16 4.4664f
C7450 m3_45124_57418# VDDR 0.0103f
C7451 a_66213_68756# VSSD 0.25932f
C7452 a_66312_50368# VSSD 0.11684f
C7453 sar10b_0._04_ sar10b_0._03_ 0.03466f
C7454 sar10b_0.CF[4] sar10b_0.CF[0] 0.1172f
C7455 sar10b_0.net39 a_61677_66174# 0.02955f
C7456 sar10b_0.net16 CLK 0.16473f
C7457 tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A a_52417_59293# 0.09051f
C7458 sar10b_0.net33 a_65996_50650# 0.01106f
C7459 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VDDR 0.38377f
C7460 VDDD sar10b_0.clk_div_0.COUNT\[0\] 1.43224f
C7461 sar10b_0.SWP[0] sar10b_0.CF[9] 0.88254f
C7462 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y 0.07418f
C7463 m3_n1472_91212# VDDR 0.02674f
C7464 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C7465 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN 0.01132f
C7466 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 sar10b_0.CF[7] 0.26243f
C7467 VDDD a_61737_56343# 0.85447f
C7468 m3_40888_97932# VCM 0.15231f
C7469 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VSSR 1.37694f
C7470 sar10b_0._16_ sar10b_0.net35 0.26085f
C7471 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.11339f
C7472 c1_n1140_33938# c1_n1140_32818# 0.13255f
C7473 sar10b_0.net32 sar10b_0._07_ 0.04692f
C7474 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04073f
C7475 sar10b_0.net45 sar10b_0.net15 0.10815f
C7476 sar10b_0.net3 a_68169_66999# 0.27548f
C7477 VDDD a_67502_56024# 0.27487f
C7478 c1_18628_97972# VCM 0.01358f
C7479 m3_45124_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C7480 VDDA a_51861_59345# 0.18641f
C7481 sar10b_0.net3 a_66645_61731# 0.22824f
C7482 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C7483 m3_n1472_35018# m3_n1472_33898# 0.29566f
C7484 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN 0.02638f
C7485 a_65589_69723# sar10b_0.net43 0.01686f
C7486 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A 0.10815f
C7487 VSSR c1_n1140_76692# 0.04956f
C7488 sar10b_0.SWN[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A 0.0108f
C7489 sar10b_0.net46 a_66825_69663# 0.013f
C7490 m3_n60_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.53633f
C7491 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[3] 0.01887f
C7492 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A 0.01751f
C7493 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A 0.07183f
C7494 a_67209_68331# VSSD 0.55091f
C7495 sar10b_0.clk_div_0.COUNT\[0\] sar10b_0._08_ 0.20728f
C7496 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A a_40248_111636# 0.01076f
C7497 sar10b_0.SWP[8] sar10b_0.CF[8] 2.36818f
C7498 c1_7332_21618# m3_8412_21578# 0.15596f
C7499 sar10b_0.SWN[3] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 0.23242f
C7500 m3_45124_52938# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C7501 sar10b_0.cyclic_flag_0.FINAL a_67055_68689# 0.17947f
C7502 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y 0.12541f
C7503 a_64705_59595# a_65045_59588# 0.24088f
C7504 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26364f
C7505 sar10b_0.net12 a_64809_65963# 0.25072f
C7506 CLK sar10b_0.CF[3] 0.20004f
C7507 m3_9824_97932# c1_10156_97972# 1.74381f
C7508 VSSR m3_45124_42858# 0.63261f
C7509 a_62623_53324# sar10b_0.net6 0.29288f
C7510 a_5051_113018# VDDR 1.62771f
C7511 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A 0.45324f
C7512 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VDDR 0.95194f
C7513 a_61491_52222# a_61773_52237# 0.06034f
C7514 c1_4508_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26825f
C7515 a_65586_50645# a_65765_50645# 0.53638f
C7516 m3_31004_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C7517 a_63169_62635# a_63945_63003# 0.3578f
C7518 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A sar10b_0.CF[9] 0.26294f
C7519 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP 2.62904f
C7520 a_67209_55011# a_67598_54692# 0.05462f
C7521 a_66933_55071# a_67393_54643# 0.26257f
C7522 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y sar10b_0.CF[3] 0.12541f
C7523 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.10847f
C7524 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN 1.14737f
C7525 VINP a_n9133_63315# 0.01178f
C7526 sar10b_0.CF[5] sar10b_0.CF[3] 0.11156f
C7527 sar10b_0.CF[6] sar10b_0.CF[2] 0.10536f
C7528 th_dif_sw_0.VCP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 8.84761f
C7529 m3_n1472_75532# m3_n1472_74412# 0.29566f
C7530 a_65119_59984# sar10b_0.net12 0.01665f
C7531 sar10b_0.SWN[1] sar10b_0.CF[2] 0.12048f
C7532 a_64428_50947# a_64356_51029# 0.22517f
C7533 VSSR m3_45124_83372# 0.63305f
C7534 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 0.68971f
C7535 a_64521_60339# a_64521_59303# 0.01915f
C7536 VDDD a_61035_71265# 0.26314f
C7537 a_67105_59971# a_68133_60292# 0.07826f
C7538 sar10b_0.net3 a_67209_55011# 0.18132f
C7539 VDDD a_68946_61735# 0.28108f
C7540 m3_45124_27178# VDDR 0.0103f
C7541 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C7542 sar10b_0.net3 a_67372_52833# 0.02309f
C7543 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP 6.773f
C7544 sar10b_0.clknet_0_CLK sar10b_0._10_ 0.02971f
C7545 sar10b_0.SWN[4] VSSD 4.77797f
C7546 m3_45124_92332# c1_45456_92372# 1.74381f
C7547 m3_n1472_92332# c1_n1140_91252# 0.01078f
C7548 m3_n1472_91212# c1_n1140_92372# 0.01078f
C7549 a_65301_57975# a_65966_58354# 0.19065f
C7550 a_61131_70891# sar10b_0.SWP[0] 0.14164f
C7551 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] m3_19708_21578# 0.13306f
C7552 a_62623_50660# sar10b_0.net6 0.01741f
C7553 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_35240_21578# 0.0162f
C7554 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.12367f
C7555 c1_36984_21618# VCM 0.01358f
C7556 c1_n1140_37298# m3_n1472_38378# 0.01078f
C7557 sar10b_0.CF[4] VSSA 0.41596f
C7558 c1_45456_38418# m3_45124_38378# 1.74381f
C7559 c1_n1140_38418# m3_n1472_37258# 0.01078f
C7560 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.11339f
C7561 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A 0.07183f
C7562 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A 0.03041f
C7563 m3_45124_67692# VDDR 0.01034f
C7564 m3_45124_64332# th_dif_sw_0.VCP 0.17339f
C7565 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 8.70956f
C7566 VSSR VDDR 4.8345p
C7567 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C7568 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP sar10b_0.SWN[4] 0.26593f
C7569 a_62133_59067# sar10b_0.net16 0.24959f
C7570 VDDD a_60747_65563# 0.28486f
C7571 a_63745_59971# a_63950_60020# 0.09983f
C7572 VDDD a_62313_61671# 0.85739f
C7573 sar10b_0.CF[0] VSSD 0.58092f
C7574 a_65397_56643# a_65673_56639# 0.1263f
C7575 sar10b_0.net9 a_60747_61567# 0.24888f
C7576 VDDD a_61929_51311# 0.35924f
C7577 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] m3_23944_21578# 0.15657f
C7578 sar10b_0.net14 sar10b_0.net16 1.47536f
C7579 a_67598_54692# sar10b_0.net35 0.02115f
C7580 sar10b_0._02_ a_65861_49313# 0.28227f
C7581 VSSD a_66921_61671# 0.5572f
C7582 a_68767_65312# sar10b_0.net25 0.26874f
C7583 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A 0.26364f
C7584 VDDD a_64993_66255# 0.2281f
C7585 VSSR c1_45456_49618# 0.09348f
C7586 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 0.24774f
C7587 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 3.56963f
C7588 sar10b_0.net3 sar10b_0.net35 0.91837f
C7589 sar10b_0.net34 a_66368_52081# 0.01662f
C7590 sar10b_0.net28 a_61249_50647# 0.01084f
C7591 VDDD a_68767_54656# 0.21528f
C7592 m3_n1472_91212# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C7593 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A 1.11457f
C7594 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] 1.8673f
C7595 sar10b_0.net4 a_60747_57571# 0.03063f
C7596 c1_45456_77812# c1_45456_76692# 0.13255f
C7597 sar10b_0.net34 a_65682_49313# 0.01959f
C7598 sar10b_0.net16 a_62261_56123# 0.13235f
C7599 m3_32416_21578# c1_31336_21618# 0.15596f
C7600 m3_n1472_28298# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C7601 DATA[6] a_68946_61735# 0.14493f
C7602 a_249_113874# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 0.07568f
C7603 a_65021_50292# VSSD 0.24584f
C7604 a_65185_68919# sar10b_0.net43 0.01264f
C7605 c1_38396_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26825f
C7606 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.4281f
C7607 VSSR sar10b_0.SWP[7] 3.84604f
C7608 m3_40888_97932# c1_39808_97972# 0.15596f
C7609 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 0.20006f
C7610 VSSR m3_7000_21578# 0.54637f
C7611 sar10b_0.SWN[4] sar10b_0.CF[8] 0.12496f
C7612 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 3.5696f
C7613 sar10b_0.net6 a_61921_55975# 0.08886f
C7614 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A sar10b_0.CF[0] 0.26303f
C7615 c1_24276_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.01445f
C7616 VDDD sar10b_0.net37 1.16237f
C7617 c1_45456_33938# VDDR 0.01151f
C7618 sar10b_0.net3 a_63810_50901# 0.03826f
C7619 m3_45124_37258# th_dif_sw_0.VCN 0.17339f
C7620 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.04073f
C7621 a_68767_62648# sar10b_0.net24 0.26931f
C7622 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A 0.28117f
C7623 a_60690_70625# VSSD 0.35859f
C7624 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y 0.07183f
C7625 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.02632f
C7626 sar10b_0.clk_div_0.COUNT\[0\] sar10b_0._15_ 0.04656f
C7627 a_68562_48647# DATA[0] 0.15514f
C7628 sar10b_0._16_ a_67419_52937# 0.09475f
C7629 m3_1352_97932# VCM 0.15231f
C7630 a_65733_59432# sar10b_0.net14 0.02891f
C7631 sar10b_0.net16 a_63457_56931# 0.09682f
C7632 VDDD a_62702_61352# 0.26883f
C7633 sar10b_0.net8 a_61395_60616# 0.01235f
C7634 sar10b_0.CF[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.40692f
C7635 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A 0.28117f
C7636 sar10b_0.net4 a_61153_67587# 0.10733f
C7637 sar10b_0.net41 a_64809_65963# 0.02648f
C7638 c1_n1140_41778# c1_n1140_40658# 0.13255f
C7639 sar10b_0.CF[0] sar10b_0.CF[8] 0.11652f
C7640 sar10b_0.CF[1] sar10b_0.CF[7] 0.113f
C7641 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y 0.32408f
C7642 a_60747_61941# a_61086_61974# 0.07649f
C7643 a_61395_61948# a_60945_61941# 0.03471f
C7644 a_66577_52883# VSSD 0.35974f
C7645 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 1.86731f
C7646 VDDD sar10b_0.SWN[7] 0.2088f
C7647 m3_26768_21578# VCM 0.13579f
C7648 m3_5588_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C7649 a_7670_8700# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01076f
C7650 sar10b_0.net38 a_60945_60609# 0.02222f
C7651 m3_n1472_42858# m3_n1472_41738# 0.29566f
C7652 VSSR c1_n1140_92372# 0.04956f
C7653 sar10b_0._08_ sar10b_0.net37 0.02357f
C7654 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VCM 7.03045f
C7655 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A 0.02842f
C7656 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.10847f
C7657 VDDA a_n8277_54565# 0.04963f
C7658 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A VSSR 0.39674f
C7659 a_64149_64635# a_64425_64631# 0.1263f
C7660 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP 3.19419f
C7661 sar10b_0.net40 a_62357_57455# 0.03932f
C7662 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VDDR 0.84026f
C7663 a_60945_65937# a_61086_65970# 0.27388f
C7664 a_66666_49313# sar10b_0.net35 0.0168f
C7665 sar10b_0.net33 a_65355_53949# 0.08727f
C7666 a_65119_59984# sar10b_0.net41 0.05146f
C7667 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A 0.02149f
C7668 VDDD a_62985_63003# 0.86835f
C7669 a_62623_53324# VSSD 0.27026f
C7670 a_66865_52076# a_67372_52243# 0.01842f
C7671 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.68875f
C7672 VSSA VSSD 11.9648f
C7673 VDDD sar10b_0.SWN[6] 0.57232f
C7674 c1_n1140_35058# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C7675 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 0.02632f
C7676 VDDD a_62185_64695# 0.30557f
C7677 sar10b_0.net3 a_68073_56343# 0.28303f
C7678 sar10b_0.net38 a_64233_56639# 0.06075f
C7679 th_dif_sw_0.VCP a_51345_58977# 0.1027f
C7680 VSSR c1_n1140_24978# 0.04956f
C7681 a_62623_50660# sar10b_0.net30 0.28517f
C7682 sar10b_0.net6 a_61833_57675# 0.02633f
C7683 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VCM 0.59213f
C7684 sar10b_0.net10 sar10b_0.net16 1.23061f
C7685 sar10b_0._01_ a_65861_51977# 0.06017f
C7686 sar10b_0.SWP[5] a_20335_112621# 0.40667f
C7687 m3_45124_67692# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C7688 VSSR cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.31308p
C7689 a_66368_49417# a_66216_49358# 0.22338f
C7690 a_65861_49313# a_66865_49412# 0.06302f
C7691 m3_n1472_83372# m3_n1472_82252# 0.29566f
C7692 sar10b_0.net13 sar10b_0.net16 1.1036f
C7693 VSSR m3_42300_97932# 0.54637f
C7694 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VCM 0.12074f
C7695 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.26364f
C7696 m3_42300_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.53746f
C7697 sar10b_0.SWP[1] sar10b_0.CF[9] 0.32484f
C7698 m3_45124_42858# VDDR 0.0103f
C7699 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 1.75141f
C7700 a_68946_63299# VSSD 0.33124f
C7701 a_66216_52022# VSSD 0.11778f
C7702 a_62181_58100# VSSD 0.2684f
C7703 VDDD a_68767_63980# 0.21793f
C7704 VSSR c1_20040_97972# 0.05454f
C7705 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN 0.01164f
C7706 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 sar10b_0.CF[3] 0.40665f
C7707 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] a_1127_5779# 0.10438f
C7708 a_62623_50660# VSSD 0.26816f
C7709 sar10b_0.net16 a_65198_66346# 0.24786f
C7710 a_65761_58263# a_66101_58256# 0.24088f
C7711 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_12648_21578# 0.03017f
C7712 a_65861_49313# VSSD 0.53919f
C7713 a_61929_67295# sar10b_0.net39 0.01774f
C7714 a_5929_5779# VSSR 0.77753f
C7715 sar10b_0.CF[6] VSSR 22.9171f
C7716 c1_10156_21618# VCM 0.01358f
C7717 sar10b_0.net34 a_66378_52993# 0.0215f
C7718 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.95198f
C7719 c1_n1140_46258# m3_n1472_45098# 0.01078f
C7720 c1_45456_46258# m3_45124_46218# 1.74381f
C7721 c1_n1140_45138# m3_n1472_46218# 0.01078f
C7722 VSSR sar10b_0.SWN[1] 5.99185f
C7723 VDDD a_62185_60699# 0.30727f
C7724 a_63339_71265# sar10b_0.SWP[3] 0.1431f
C7725 VDDD sar10b_0._03_ 1.13151f
C7726 a_60945_63273# a_61609_63602# 0.16939f
C7727 a_61395_63280# a_61677_63510# 0.05462f
C7728 m3_45124_80012# th_dif_sw_0.VCP 0.17339f
C7729 m3_45124_83372# VDDR 0.01034f
C7730 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSSR 2.4554f
C7731 VDDD sar10b_0.CF[7] 0.37773f
C7732 sar10b_0.net46 sar10b_0.net16 0.11838f
C7733 sar10b_0.net9 a_61395_60616# 0.05106f
C7734 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN sar10b_0.CF[9] 0.03484f
C7735 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[8] 0.17717f
C7736 sar10b_0._04_ sar10b_0._13_ 0.02397f
C7737 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A 0.03718f
C7738 VSSA sar10b_0.CF[8] 0.11513f
C7739 a_63573_63303# sar10b_0.net2 0.18388f
C7740 a_62133_59067# a_62798_58688# 0.19065f
C7741 a_62409_59007# a_62933_58787# 0.04522f
C7742 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 a_15533_5779# 0.28343f
C7743 sar10b_0.CF[2] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.01366f
C7744 c1_39808_97972# VCM 0.01358f
C7745 sar10b_0.net45 a_66933_65727# 0.18792f
C7746 m3_45124_68812# c1_45456_67732# 0.01078f
C7747 m3_45124_67692# c1_45456_68852# 0.01078f
C7748 m3_n1472_67692# c1_n1140_67732# 1.74381f
C7749 sar10b_0.net13 a_60969_67295# 0.05676f
C7750 VSSR c1_45456_68852# 0.0935f
C7751 a_68946_71059# VSSD 0.33334f
C7752 a_60747_49953# VSSD 0.25842f
C7753 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C7754 sar10b_0.CF[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.10395f
C7755 m3_21120_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.21656f
C7756 sar10b_0.net19 sar10b_0._14_ 0.33546f
C7757 c1_44044_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C7758 a_60693_67299# VSSD 0.14809f
C7759 sar10b_0._03_ sar10b_0._08_ 0.03527f
C7760 sar10b_0._07_ a_64339_51661# 0.04525f
C7761 m3_31004_97932# m3_32416_97932# 0.23959f
C7762 a_61493_51596# a_61929_51311# 0.16939f
C7763 a_67209_64335# a_67393_63967# 0.44098f
C7764 c1_45456_85652# c1_45456_84532# 0.13255f
C7765 c1_18628_21618# m3_18296_21578# 1.74381f
C7766 sar10b_0.CF[4] th_dif_sw_0.VCN 0.2926f
C7767 th_dif_sw_0.CK sar10b_0.CF[9] 4.5303f
C7768 VDDD a_60945_52617# 0.40365f
C7769 m3_n1472_43978# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C7770 sar10b_0.net5 a_60969_56639# 0.21793f
C7771 a_60693_56643# a_61153_56931# 0.26257f
C7772 sar10b_0.net16 a_63525_61624# 0.17428f
C7773 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.53307f
C7774 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A 0.03718f
C7775 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_41284_111642# 0.01076f
C7776 a_68479_59984# VSSD 0.27636f
C7777 m3_21120_97932# c1_20040_97972# 0.15596f
C7778 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 0.19508f
C7779 a_64809_65963# a_64993_66255# 0.44532f
C7780 VSSD a_61921_55975# 0.8535f
C7781 VSSR m3_n1472_33898# 0.66371f
C7782 sar10b_0.net13 a_60747_68227# 0.26298f
C7783 sar10b_0.net16 a_62997_67299# 0.25901f
C7784 sar10b_0.CF[5] sar10b_0.SWP[4] 0.1187f
C7785 a_19457_110450# VSSR 0.06033f
C7786 VCM sar10b_0.SWP[3] 0.13075f
C7787 sar10b_0.net3 a_67393_65299# 0.11277f
C7788 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VCM 0.1236f
C7789 sar10b_0._15_ sar10b_0.net37 0.15046f
C7790 sar10b_0.net18 DATA[1] 0.06811f
C7791 c1_45456_49618# VDDR 0.01151f
C7792 m3_45124_52938# th_dif_sw_0.VCN 0.17339f
C7793 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VCM 0.12068f
C7794 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP a_29939_111781# 0.01299f
C7795 sar10b_0.SWN[2] sar10b_0.SWN[3] 10.8367f
C7796 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C7797 VDDA a_53564_60302# 0.51472f
C7798 VDDD sar10b_0.SWN[5] 0.22256f
C7799 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A 1.37832f
C7800 VSSR c1_38396_21618# 0.05923f
C7801 sar10b_0.net3 sar10b_0.net44 0.13646f
C7802 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A 0.95194f
C7803 a_60747_60609# a_60945_60609# 0.06623f
C7804 a_38665_107026# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.92132f
C7805 a_68169_55011# a_68767_54656# 0.06623f
C7806 sar10b_0._07_ CLK 0.13891f
C7807 VSSR m3_n1472_74412# 0.66316f
C7808 sar10b_0.net33 sar10b_0.net34 0.68369f
C7809 c1_n1140_49618# c1_n1140_48498# 0.13255f
C7810 a_65586_50645# sar10b_0.net16 0.21093f
C7811 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38365f
C7812 VDDR sar10b_0.SWP[7] 1.55419f
C7813 sar10b_0.net14 a_65390_69010# 0.0729f
C7814 a_63509_62783# sar10b_0.net16 0.14458f
C7815 a_25137_112201# VSSR 2.12959f
C7816 a_62261_56123# a_62697_56343# 0.16939f
C7817 m3_n1472_26058# VCM 0.01415f
C7818 c1_n1140_76692# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C7819 m3_n1472_50698# m3_n1472_49578# 0.29566f
C7820 sar10b_0.CF[0] sar10b_0.SWN[0] 4.2303f
C7821 sar10b_0._01_ a_65996_50650# 0.12213f
C7822 VDDD a_61395_65944# 0.8671f
C7823 sar10b_0.net21 a_68671_55988# 0.02149f
C7824 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VSSR 1.37552f
C7825 a_68169_55011# sar10b_0.net37 0.02485f
C7826 VSSR a_43467_5788# 0.05969f
C7827 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A 0.26294f
C7828 sar10b_0._04_ a_66368_52081# 0.01997f
C7829 a_65682_51977# a_66666_51977# 0.08669f
C7830 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 3.69121f
C7831 sar10b_0.net39 a_61609_64934# 0.01413f
C7832 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 0.56487f
C7833 sar10b_0.SWP[4] a_24259_109594# 0.64881f
C7834 a_65577_51311# a_65765_50645# 0.05376f
C7835 c1_22864_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.01237f
C7836 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y 0.31995f
C7837 m3_n1472_66572# VCM 0.01412f
C7838 VDDD sar10b_0.net25 0.68585f
C7839 sar10b_0.SWN[0] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.23768f
C7840 VDDD a_65525_68912# 0.20245f
C7841 sar10b_0.net33 a_66197_56924# 0.01399f
C7842 a_67393_66631# a_67733_66779# 0.24088f
C7843 a_64033_63591# a_64373_63584# 0.24088f
C7844 a_63849_63299# a_64809_63299# 0.03432f
C7845 sar10b_0.net2 a_60969_56639# 0.03072f
C7846 VDDD a_66464_50363# 0.10435f
C7847 c1_n1140_50738# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C7848 a_63369_59007# sar10b_0.net39 0.09468f
C7849 sar10b_0._11_ a_64338_52411# 0.29092f
C7850 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.95198f
C7851 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A VDDR 0.60103f
C7852 sar10b_0.net40 a_61400_62288# 0.02425f
C7853 VSSD a_61833_57675# 0.49096f
C7854 sar10b_0._05_ a_65928_53032# 0.04234f
C7855 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN 3.3783f
C7856 VSSR c1_n1140_40658# 0.04956f
C7857 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] 2.31287f
C7858 a_68421_58960# VSSD 0.2719f
C7859 m3_45124_83372# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C7860 m3_n1472_91212# m3_n1472_90092# 0.29566f
C7861 VSSR m3_2764_97932# 0.54637f
C7862 m3_42300_21578# c1_42632_21618# 1.74381f
C7863 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y 0.07418f
C7864 sar10b_0.net16 a_61395_61948# 0.18243f
C7865 m3_2764_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.53746f
C7866 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN 0.02638f
C7867 sar10b_0.clk_div_0.COUNT\[1\] a_67564_50907# 0.14157f
C7868 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A 0.11547f
C7869 a_66666_51977# sar10b_0._07_ 0.05576f
C7870 tdc_0.phase_detector_0.INP a_53564_60302# 0.01369f
C7871 a_63457_56931# a_64233_56639# 0.3578f
C7872 a_64373_63584# sar10b_0.net42 0.0137f
C7873 m3_n1472_94572# c1_n1140_95732# 0.01078f
C7874 m3_45124_95692# c1_45456_95732# 1.74381f
C7875 m3_n1472_95692# c1_n1140_94612# 0.01078f
C7876 sar10b_0.net16 a_60945_65937# 0.29219f
C7877 VSSR m3_28180_21578# 0.46562f
C7878 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C7879 sar10b_0.CF[2] sar10b_0.CF[7] 0.10502f
C7880 a_51861_59345# tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A 0.16495f
C7881 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C7882 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 3.0756f
C7883 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.01165f
C7884 sar10b_0.net3 a_64199_50761# 0.01515f
C7885 c1_n1140_52978# m3_n1472_54058# 0.01078f
C7886 c1_45456_54098# m3_45124_54058# 1.74381f
C7887 c1_n1140_54098# m3_n1472_52938# 0.01078f
C7888 a_66795_71265# VSSD 0.33655f
C7889 a_65001_68627# sar10b_0.net41 0.0136f
C7890 VDDR cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 16.0474f
C7891 VSSD a_65769_65963# 0.29541f
C7892 a_61065_53679# VSSD 0.49348f
C7893 sar10b_0.clknet_0_CLK a_66312_50368# 0.05512f
C7894 sar10b_0.SWP[5] VSSD 0.98648f
C7895 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A 0.26364f
C7896 m3_45124_95692# th_dif_sw_0.VCP 0.17339f
C7897 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.39835f
C7898 m3_22532_97932# VCM 0.11203f
C7899 th_dif_sw_0.th_sw_1.CK th_dif_sw_0.th_sw_1.CKB 4.72448f
C7900 a_61677_52854# sar10b_0.net16 0.27974f
C7901 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_44044_21618# 0.0106f
C7902 sar10b_0.net8 a_60747_60235# 0.24795f
C7903 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45324f
C7904 c1_272_97972# VCM 0.01358f
C7905 m3_26768_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C7906 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A 0.11547f
C7907 a_64705_59595# sar10b_0.net1 0.06981f
C7908 m3_45124_75532# c1_45456_76692# 0.01078f
C7909 m3_45124_76652# c1_45456_75572# 0.01078f
C7910 m3_n1472_75532# c1_n1140_75572# 1.74381f
C7911 VSSR c1_45456_84532# 0.0935f
C7912 sar10b_0.SWN[0] VSSA 0.2658f
C7913 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.02632f
C7914 sar10b_0.CF[6] VDDR 1.74393f
C7915 sar10b_0.net23 sar10b_0.net3 0.20825f
C7916 sar10b_0.net38 a_61400_62288# 0.02065f
C7917 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN 0.02638f
C7918 VDDR sar10b_0.SWN[1] 3.45046f
C7919 sar10b_0.cyclic_flag_0.FINAL a_67209_66999# 0.24116f
C7920 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.07418f
C7921 a_61131_70891# sar10b_0.net2 0.05743f
C7922 sar10b_0.net13 a_65390_69010# 0.05809f
C7923 c1_4508_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C7924 m3_11236_97932# m3_12648_97932# 0.23959f
C7925 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VDDR 2.61522f
C7926 c1_45456_93492# c1_45456_92372# 0.13255f
C7927 c1_n1140_21618# m3_n1472_21578# 1.74381f
C7928 sar10b_0.net40 a_66389_57455# 0.0535f
C7929 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A sar10b_0.CF[7] 0.03041f
C7930 VSSR cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.16481p
C7931 VDDD a_66933_63063# 0.32502f
C7932 m3_1352_97932# c1_272_97972# 0.15596f
C7933 VSSR m3_n1472_49578# 0.66371f
C7934 c1_28512_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.26825f
C7935 a_67598_68012# a_67733_68111# 0.35559f
C7936 a_67209_68331# a_68421_68284# 0.07766f
C7937 c1_45456_68852# VDDR 0.01153f
C7938 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] m3_22532_97932# 0.59433f
C7939 th_dif_sw_0.VCN sar10b_0.CF[8] 0.28587f
C7940 m3_12648_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C7941 sar10b_0.net1 a_65397_56643# 0.17339f
C7942 m3_36652_21578# m3_38064_21578# 0.23959f
C7943 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 0.9283f
C7944 VSSR c1_11568_21618# 0.05685f
C7945 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.01165f
C7946 sar10b_0.SWP[5] sar10b_0.CF[8] 0.12388f
C7947 a_62017_57307# a_62222_57356# 0.09983f
C7948 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A 0.43728f
C7949 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A sar10b_0.SWN[6] 0.01364f
C7950 a_67372_52833# sar10b_0.clk_div_0.COUNT\[3\] 0.13721f
C7951 m3_22532_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 0.59433f
C7952 a_64033_63591# sar10b_0.net16 0.11841f
C7953 VSSR m3_n1472_90092# 0.66316f
C7954 c1_n1140_57458# c1_n1140_56338# 0.13255f
C7955 a_66921_60339# a_66645_60399# 0.1263f
C7956 sar10b_0.net7 a_60969_56639# 0.01015f
C7957 m3_n1472_33898# VDDR 0.02681f
C7958 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A 0.03718f
C7959 tdc_0.phase_detector_0.INN tdc_0.phase_detector_0.pd_out_0.B 0.03294f
C7960 a_19457_110450# VDDR 4.02021f
C7961 m3_n1472_41738# VCM 0.01415f
C7962 c1_n1140_92372# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C7963 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP a_33863_5788# 0.19132f
C7964 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A a_35446_111636# 0.01076f
C7965 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN 3.87099f
C7966 a_61677_64842# a_62185_64695# 0.19065f
C7967 VSSR c1_41220_97972# 0.05923f
C7968 a_63169_62635# VSSD 0.88416f
C7969 VSSR sar10b_0.SWN[7] 3.91401f
C7970 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A 0.83558f
C7971 sar10b_0.net4 sar10b_0.net5 1.37546f
C7972 th_dif_sw_0.CKB sar10b_0.SWN[2] 0.02596f
C7973 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_33828_21578# 0.03017f
C7974 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_16884_21578# 0.0162f
C7975 th_dif_sw_0.VCP VDDA 1.58681f
C7976 a_61358_51694# sar10b_0.net16 0.23618f
C7977 VDDD a_62185_50043# 0.30381f
C7978 VDDD sar10b_0.net15 0.57509f
C7979 a_66933_59067# sar10b_0.cyclic_flag_0.FINAL 0.05554f
C7980 m3_n1472_74412# VDDR 0.02674f
C7981 m3_n1472_82252# VCM 0.01412f
C7982 m3_21120_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.1528f
C7983 a_40248_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A 0.01076f
C7984 sar10b_0.net16 sar10b_0.net42 1.13285f
C7985 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP sar10b_0.CF[9] 0.10502f
C7986 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.01751f
C7987 c1_45456_26098# c1_45456_24978# 0.13255f
C7988 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN sar10b_0.CF[5] 0.08506f
C7989 VDDD EN 0.38815f
C7990 sar10b_0.clk_div_0.COUNT\[3\] sar10b_0.net35 0.04238f
C7991 sar10b_0.net32 VSSD 2.32308f
C7992 a_61929_57971# sar10b_0.net2 0.01246f
C7993 VDDD a_64521_59303# 0.83937f
C7994 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VDDR 0.83965f
C7995 a_67393_65299# a_68169_65667# 0.3578f
C7996 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP sar10b_0.CF[9] 0.19143f
C7997 VDDD sar10b_0._13_ 0.61845f
C7998 a_43467_5788# VDDR 8.00721f
C7999 m3_45124_27178# m3_45124_26058# 0.29566f
C8000 VSSR sar10b_0.SWN[6] 4.24189f
C8001 VSSR c1_n1140_56338# 0.04956f
C8002 a_64924_52385# a_65188_51977# 0.01136f
C8003 sar10b_0.net19 a_68946_52411# 0.01098f
C8004 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 2.69124f
C8005 a_68479_61316# sar10b_0.net22 0.27328f
C8006 a_66389_69443# VSSD 0.10029f
C8007 m3_42300_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.53746f
C8008 m3_18296_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.18044f
C8009 a_68169_64335# a_68767_63980# 0.06623f
C8010 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 0.24776f
C8011 m3_22532_21578# c1_22864_21618# 1.74381f
C8012 m3_45124_36138# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C8013 VDDD a_65928_53032# 0.14189f
C8014 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP a_29061_5788# 0.16709f
C8015 a_61153_56931# a_61358_57022# 0.09983f
C8016 sar10b_0.net33 sar10b_0._04_ 0.04275f
C8017 a_62181_56768# a_61929_56639# 0.27388f
C8018 m3_31004_97932# c1_31336_97972# 1.74381f
C8019 VSSR m3_45124_26058# 0.63261f
C8020 a_61395_49960# a_61086_49986# 0.07766f
C8021 sar10b_0.cyclic_flag_0.FINAL sar10b_0.net3 3.22052f
C8022 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A 0.05472f
C8023 sar10b_0._13_ sar10b_0._08_ 0.0226f
C8024 c1_34160_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26825f
C8025 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.05472f
C8026 sar10b_0.net43 a_65333_66248# 0.01319f
C8027 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 sar10b_0.SWN[9] 0.35379f
C8028 a_67393_62635# a_68169_63003# 0.3578f
C8029 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.40046f
C8030 a_61677_60846# a_62185_60699# 0.19065f
C8031 VDDD a_62277_53632# 0.27294f
C8032 sar10b_0.net2 sar10b_0.net4 0.09474f
C8033 a_66933_68391# sar10b_0.net45 0.02373f
C8034 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_17216_21618# 0.0106f
C8035 sar10b_0.net41 sar10b_0.net12 1.26426f
C8036 sar10b_0.net16 a_62181_56768# 0.1981f
C8037 m3_45124_67692# m3_45124_66572# 0.29566f
C8038 VSSR m3_45124_66572# 0.63305f
C8039 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 3.47757f
C8040 VSSR sar10b_0.CF[7] 24.2161f
C8041 sar10b_0.net2 a_62126_56024# 0.01526f
C8042 sar10b_0.net32 sar10b_0.net31 0.26784f
C8043 m3_8412_21578# VCM 0.15231f
C8044 sar10b_0.net6 a_61153_56931# 0.01644f
C8045 sar10b_0.CF[6] sar10b_0.SWN[1] 0.12428f
C8046 m3_45124_83372# c1_45456_84532# 0.01078f
C8047 m3_45124_84492# c1_45456_83412# 0.01078f
C8048 m3_n1472_83372# c1_n1140_83412# 1.74381f
C8049 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] th_dif_sw_0.VCP 4.58977f
C8050 sar10b_0.clknet_0_CLK a_66577_52883# 0.02701f
C8051 m3_18296_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 0.32786f
C8052 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VCM 0.12735f
C8053 a_61419_71265# sar10b_0.net16 0.26512f
C8054 sar10b_0.net3 a_67393_67963# 0.09211f
C8055 c1_n1140_29458# m3_n1472_29418# 1.74381f
C8056 c1_45456_30578# m3_45124_29418# 0.01078f
C8057 c1_45456_29458# m3_45124_30538# 0.01078f
C8058 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP 3.50689f
C8059 sar10b_0.net38 a_67113_56343# 0.01597f
C8060 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y 0.36435f
C8061 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 sar10b_0.CF[2] 0.26279f
C8062 VDDD a_66368_52081# 0.09825f
C8063 VDDD a_61493_58256# 0.20965f
C8064 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VSSR 1.3479f
C8065 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 0.24487f
C8066 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A 0.42509f
C8067 a_61773_52237# a_61705_51992# 0.35559f
C8068 VDDD a_62277_50968# 0.2588f
C8069 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45324f
C8070 a_60693_57975# a_61153_58263# 0.26257f
C8071 a_n8277_54249# th_dif_sw_0.th_sw_1.CK 0.05273f
C8072 VDDD a_65682_49313# 0.43067f
C8073 c1_45456_84532# VDDR 0.01153f
C8074 VSSR a_1127_114301# 0.4375f
C8075 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A 0.07418f
C8076 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A 0.03718f
C8077 a_66921_61671# a_67881_61671# 0.03471f
C8078 a_67105_61303# a_67310_61352# 0.09983f
C8079 a_60789_53739# sar10b_0.net5 0.19105f
C8080 m3_16884_21578# m3_18296_21578# 0.23959f
C8081 sar10b_0.SWP[2] sar10b_0.SWP[1] 9.06167f
C8082 VSSD a_65589_57735# 0.14119f
C8083 tdc_0.OUTP sar10b_0.CF[9] 0.25141f
C8084 sar10b_0._09_ sar10b_0._01_ 0.02523f
C8085 VSSR c1_45456_32818# 0.09348f
C8086 sar10b_0.net4 a_61249_53311# 0.06782f
C8087 a_65857_56931# a_66062_57022# 0.09983f
C8088 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A 0.11547f
C8089 sar10b_0.CF[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A 0.02149f
C8090 VSSR a_14655_111306# 0.06033f
C8091 m3_n1472_74412# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C8092 VSSR sar10b_0.SWN[5] 4.55583f
C8093 VSSR m3_23944_97932# 0.41298f
C8094 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A 0.28117f
C8095 c1_n1140_68852# c1_n1140_67732# 0.13255f
C8096 sar10b_0.net33 sar10b_0._05_ 0.11524f
C8097 sar10b_0.net16 sar10b_0.net8 0.8733f
C8098 VDDR cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 14.4489f
C8099 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 0.40988f
C8100 m3_23944_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26603f
C8101 m3_n1472_49578# VDDR 0.02681f
C8102 a_60747_52617# a_60945_52617# 0.06623f
C8103 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A 0.02842f
C8104 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A 0.45324f
C8105 a_63849_63299# VSSD 0.54061f
C8106 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[3] 0.05939f
C8107 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A sar10b_0.SWP[1] 0.02059f
C8108 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[5] 0.17717f
C8109 sar10b_0.net1 a_62017_57307# 0.01915f
C8110 VSSR c1_1684_97972# 0.05923f
C8111 a_65045_59588# sar10b_0.net16 0.15712f
C8112 a_66559_68962# VSSD 0.25103f
C8113 a_67598_62684# sar10b_0.net3 0.26268f
C8114 VSSA th_dif_sw_0.th_sw_1.CK 8.23354f
C8115 a_67439_50041# VSSD 0.13504f
C8116 sar10b_0.net2 a_61557_57735# 0.2575f
C8117 sar10b_0._17_ a_67084_53565# 0.09895f
C8118 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 0.88327f
C8119 sar10b_0.SWP[0] a_43467_106170# 1.0688f
C8120 a_68169_64335# sar10b_0.net25 0.01141f
C8121 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A VDDR 0.38397f
C8122 a_63273_67295# a_63804_67580# 0.04775f
C8123 a_62997_67299# a_63457_67583# 0.25898f
C8124 sar10b_0.net38 sar10b_0.net6 0.15912f
C8125 sar10b_0.clknet_0_CLK a_65861_49313# 0.0191f
C8126 m3_n1472_90092# VDDR 0.02674f
C8127 VDDD a_68133_60292# 0.27633f
C8128 m3_43712_97932# VCM 0.15231f
C8129 sar10b_0.clk_div_0.COUNT\[3\] a_67419_52937# 0.0217f
C8130 sar10b_0.net40 a_65857_56931# 0.02105f
C8131 CLK sar10b_0.net6 0.05079f
C8132 c1_45456_33938# c1_45456_32818# 0.13255f
C8133 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A 0.42509f
C8134 sar10b_0.SWN[8] VSSA 0.24847f
C8135 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.41046f
C8136 sar10b_0.net2 a_64725_68631# 0.17486f
C8137 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.20752f
C8138 VDDR sar10b_0.SWN[7] 1.48436f
C8139 c1_21452_97972# VCM 0.01311f
C8140 sar10b_0._13_ sar10b_0._15_ 0.02658f
C8141 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 0.1901f
C8142 a_63950_60020# sar10b_0.net16 0.23502f
C8143 m3_45124_35018# m3_45124_33898# 0.29566f
C8144 w_n9655_63119# a_n8277_65767# 0.05534f
C8145 sar10b_0.net16 a_65673_56639# 0.16815f
C8146 sar10b_0.net34 a_65778_49979# 0.02115f
C8147 VSSR c1_n1140_75572# 0.04956f
C8148 a_65643_48621# sar10b_0.SWN[5] 0.15514f
C8149 sar10b_0.net12 a_60747_65563# 0.28154f
C8150 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VCM 3.13306f
C8151 sar10b_0.net7 sar10b_0.net4 0.48682f
C8152 m3_2764_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.53746f
C8153 c1_25688_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C8154 m3_n1472_97932# m3_n1472_96812# 0.29566f
C8155 c1_8744_21618# m3_9824_21578# 0.15596f
C8156 m3_45124_51818# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C8157 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A 0.41861f
C8158 VDDD a_63273_56639# 0.83923f
C8159 a_64705_59595# a_65481_59303# 0.3578f
C8160 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A sar10b_0.CF[3] 0.02149f
C8161 sar10b_0.net12 a_64993_66255# 0.04659f
C8162 m3_11236_97932# c1_11568_97972# 1.74381f
C8163 VSSD a_66062_57022# 0.13048f
C8164 a_60693_51315# CLK 0.01487f
C8165 VSSR m3_45124_41738# 0.63261f
C8166 sar10b_0.SWN[9] VSSA 0.2591f
C8167 VDDR sar10b_0.SWN[6] 1.81289f
C8168 sar10b_0.clk_div_0.COUNT\[0\] a_67611_50645# 0.03884f
C8169 sar10b_0.net47 a_67209_68331# 0.06924f
C8170 c1_7332_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26825f
C8171 a_65586_50645# a_66103_50668# 0.33885f
C8172 sar10b_0.CF[4] CLK 0.10143f
C8173 a_65765_50645# a_66255_50749# 0.23951f
C8174 m3_33828_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C8175 a_63509_62783# a_63945_63003# 0.16939f
C8176 sar10b_0.SWP[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A 0.0196f
C8177 sar10b_0.SWN[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.23393f
C8178 VSSR c1_20040_21618# 0.05454f
C8179 a_64425_64631# sar10b_0.net16 0.18413f
C8180 VDDD sar10b_0.clknet_1_0__leaf_CLK 2.70388f
C8181 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] c1_21452_97972# 0.28822f
C8182 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[7] 0.05939f
C8183 m3_45124_75532# m3_45124_74412# 0.29566f
C8184 a_64199_50761# sar10b_0._00_ 0.26229f
C8185 sar10b_0.net9 sar10b_0.net16 0.9087f
C8186 VSSR m3_45124_82252# 0.63305f
C8187 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VCM 2.92973f
C8188 VDDD a_66378_52993# 0.0946f
C8189 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 17.511f
C8190 a_65119_59984# a_64521_59303# 0.0165f
C8191 sar10b_0.net38 a_65857_56931# 0.01309f
C8192 sar10b_0.net40 a_61400_64952# 0.02782f
C8193 m3_45124_26058# VDDR 0.0103f
C8194 VSSD a_61153_56931# 0.84919f
C8195 sar10b_0.CF[5] sar10b_0.CF[4] 54.1596f
C8196 VSSD sar10b_0.SWP[6] 0.9412f
C8197 sar10b_0.clknet_1_1__leaf_CLK sar10b_0._10_ 0.63131f
C8198 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VCM 0.12358f
C8199 m3_45124_92332# c1_45456_91252# 0.01078f
C8200 m3_n1472_91212# c1_n1140_91252# 1.74381f
C8201 m3_45124_91212# c1_45456_92372# 0.01078f
C8202 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A sar10b_0.CF[0] 0.06396f
C8203 a_67393_62635# VSSD 0.85606f
C8204 VDDD a_68169_59007# 0.36741f
C8205 sar10b_0.net16 a_61395_64612# 0.18967f
C8206 sar10b_0.net40 VSSD 4.61774f
C8207 a_60789_53739# a_61249_53311# 0.26257f
C8208 a_61065_53679# a_61454_53360# 0.05462f
C8209 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_38064_21578# 0.0162f
C8210 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.45324f
C8211 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_36482_111642# 0.01076f
C8212 sar10b_0.net16 a_66101_58256# 0.1647f
C8213 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A VSSR 0.43773f
C8214 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VCM 4.1148f
C8215 c1_39808_21618# VCM 0.01358f
C8216 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.12068f
C8217 c1_45456_38418# m3_45124_37258# 0.01078f
C8218 c1_45456_37298# m3_45124_38378# 0.01078f
C8219 c1_n1140_37298# m3_n1472_37258# 1.74381f
C8220 VDDD a_61677_63510# 0.26819f
C8221 a_67113_56343# a_68325_56296# 0.07766f
C8222 a_67297_55975# a_67637_56123# 0.24088f
C8223 sar10b_0._08_ sar10b_0.clknet_1_0__leaf_CLK 0.01445f
C8224 m3_45124_66572# VDDR 0.01034f
C8225 sar10b_0._04_ a_68841_51605# 0.02238f
C8226 m3_45124_63212# th_dif_sw_0.VCP 0.17719f
C8227 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 32.8146f
C8228 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 2.67074f
C8229 sar10b_0.net34 sar10b_0.net35 0.11968f
C8230 c1_17216_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.28565f
C8231 VDDR sar10b_0.CF[7] 1.75614f
C8232 a_62593_58639# sar10b_0.net16 0.09292f
C8233 a_63950_60020# a_64085_60119# 0.35559f
C8234 VDDD a_66933_65727# 0.32431f
C8235 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.08106f
C8236 sar10b_0.net28 a_61803_48621# 0.25699f
C8237 VSSD a_68421_66952# 0.27173f
C8238 DATA[8] a_68946_65963# 0.15087f
C8239 VDDD sar10b_0.net28 0.62457f
C8240 sar10b_0.net40 a_61400_60956# 0.02253f
C8241 sar10b_0.net7 a_61557_57735# 0.04908f
C8242 sar10b_0._02_ a_66109_49318# 0.11865f
C8243 VSSR a_34741_5779# 2.80455f
C8244 a_63374_62684# sar10b_0.net2 0.07566f
C8245 VDDD a_66021_66092# 0.27638f
C8246 a_65001_68627# a_65525_68912# 0.05022f
C8247 VDDD a_68946_53975# 0.27883f
C8248 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VCM 0.12734f
C8249 th_dif_sw_0.CK a_n8277_66083# 0.05224f
C8250 VSSR c1_45456_48498# 0.09348f
C8251 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 2.55256f
C8252 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A sar10b_0.CF[2] 0.26294f
C8253 sar10b_0.net28 a_61589_50795# 0.0149f
C8254 sar10b_0.CF[4] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] 0.01357f
C8255 m3_n1472_90092# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C8256 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR 0.59739f
C8257 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VDDR 0.75026f
C8258 c1_n1140_76692# c1_n1140_75572# 0.13255f
C8259 a_64339_51661# VSSD 0.2899f
C8260 m3_33828_21578# c1_32748_21618# 0.15596f
C8261 a_66027_53575# sar10b_0._17_ 0.2575f
C8262 m3_n1472_27178# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C8263 c1_41220_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26825f
C8264 a_66825_69663# a_67077_69616# 0.27388f
C8265 VCM cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 0.12068f
C8266 sar10b_0.SWP[7] sar10b_0.CF[7] 2.46901f
C8267 sar10b_0.CF[8] sar10b_0.SWP[6] 0.12317f
C8268 m3_42300_97932# c1_41220_97972# 0.15596f
C8269 VSSR m3_9824_21578# 0.4731f
C8270 a_62798_58688# sar10b_0.net8 0.02456f
C8271 sar10b_0.net6 a_62261_56123# 0.0582f
C8272 VDDD sar10b_0.net33 2.07758f
C8273 c1_27100_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 0.01078f
C8274 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A 1.12023f
C8275 c1_45456_32818# VDDR 0.01151f
C8276 m3_45124_36138# th_dif_sw_0.VCN 0.17339f
C8277 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 sar10b_0.SWN[9] 0.2346f
C8278 a_67055_68689# sar10b_0.net16 0.09867f
C8279 a_61395_63280# sar10b_0.net4 0.22034f
C8280 sar10b_0.net3 a_66368_49417# 0.04963f
C8281 sar10b_0.net7 a_60789_53739# 0.0317f
C8282 sar10b_0.net38 VSSD 2.0444f
C8283 VDDR a_14655_111306# 3.22284f
C8284 a_55121_59650# tdc_0.phase_detector_0.pd_out_0.B 0.36537f
C8285 VDDR sar10b_0.SWN[5] 2.15554f
C8286 sar10b_0.SWN[7] DATA[0] 0.10131f
C8287 m3_32416_97932# th_dif_sw_0.VCP 0.01078f
C8288 VSSR a_25137_5779# 2.12959f
C8289 m3_4176_97932# VCM 0.15231f
C8290 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 0.32628f
C8291 VSSD CLK 1.9204f
C8292 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_25688_21618# 0.0106f
C8293 sar10b_0.net16 a_64485_56768# 0.17271f
C8294 a_66933_55071# VSSD 0.13832f
C8295 sar10b_0.net4 a_62181_67424# 0.05843f
C8296 a_68946_59303# DATA[5] 0.1424f
C8297 c1_45456_41778# c1_45456_40658# 0.13255f
C8298 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 sar10b_0.CF[2] 0.26283f
C8299 c1_10156_97972# th_dif_sw_0.VCP 0.13255f
C8300 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN sar10b_0.CF[8] 0.12367f
C8301 a_60945_61941# a_61086_61974# 0.27388f
C8302 a_61395_61948# a_61400_62288# 0.44098f
C8303 sar10b_0._14_ VSSD 0.66956f
C8304 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 30.4789f
C8305 m3_29592_21578# VCM 0.13579f
C8306 m3_8412_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C8307 sar10b_0.net38 a_61400_60956# 0.01875f
C8308 m3_45124_42858# m3_45124_41738# 0.29566f
C8309 VSSR EN 11.1479f
C8310 sar10b_0.net33 sar10b_0._08_ 0.02208f
C8311 VSSR c1_n1140_91252# 0.04956f
C8312 sar10b_0.CF[7] sar10b_0.net12 0.01224f
C8313 a_66933_64395# sar10b_0.net3 0.23565f
C8314 sar10b_0.net24 a_68479_61316# 0.01569f
C8315 th_dif_sw_0.VCN th_dif_sw_0.th_sw_1.CK 0.85764f
C8316 sar10b_0.CF[5] VSSD 0.82444f
C8317 a_64149_64635# a_64609_64923# 0.26257f
C8318 tdc_0.OUTP tdc_0.phase_detector_0.pd_out_0.B 0.3649f
C8319 a_61086_65970# a_61400_66284# 0.07826f
C8320 sar10b_0.net14 a_65857_56931# 0.0395f
C8321 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.05105f
C8322 a_67372_52243# a_67696_52265# 0.23197f
C8323 sar10b_0.CF[6] sar10b_0.SWN[6] 2.43682f
C8324 a_67372_52243# sar10b_0.clk_div_0.COUNT\[1\] 0.13647f
C8325 sar10b_0.net16 a_62222_57356# 0.25176f
C8326 c1_n1140_33938# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C8327 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP 0.17513f
C8328 a_64924_52385# sar10b_0.net16 0.10679f
C8329 sar10b_0.net46 a_66933_67059# 0.17172f
C8330 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 3.25676f
C8331 sar10b_0.net42 a_63457_67583# 0.01582f
C8332 sar10b_0.net38 sar10b_0.net31 0.09934f
C8333 VSSR c1_n1140_23858# 0.04956f
C8334 VDDA sar10b_0.SWP[0] 0.26662f
C8335 sar10b_0.CF[5] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y 0.12541f
C8336 a_64491_48621# VSSD 0.36572f
C8337 sar10b_0.SWP[6] a_15533_113041# 0.32874f
C8338 VDDD a_62281_52347# 0.28909f
C8339 m3_45124_66572# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C8340 a_66368_49417# a_66666_49313# 0.02614f
C8341 CLK sar10b_0.CF[8] 0.09352f
C8342 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] sar10b_0.CF[8] 0.01331f
C8343 CLK sar10b_0.net31 0.04478f
C8344 m3_45124_83372# m3_45124_82252# 0.29566f
C8345 VSSR m3_45124_97932# 0.68166f
C8346 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 1.73977f
C8347 m3_45124_41738# VDDR 0.0103f
C8348 a_66666_51977# VSSD 0.19834f
C8349 sar10b_0.SWN[2] sar10b_0.CF[3] 0.12021f
C8350 a_62527_58306# VSSD 0.2611f
C8351 a_67393_58639# a_68421_58960# 0.07826f
C8352 a_60747_64605# a_61086_64638# 0.07649f
C8353 a_61395_64612# a_60945_64605# 0.03471f
C8354 VSSR c1_22864_97972# 0.05003f
C8355 a_63945_63003# sar10b_0.net42 0.02136f
C8356 a_65682_51977# a_65577_51311# 0.01154f
C8357 VDDD a_66254_69344# 0.27327f
C8358 a_63918_50969# VSSD 0.24952f
C8359 sar10b_0.net18 DATA[2] 0.10076f
C8360 a_65761_58263# a_66537_57971# 0.3578f
C8361 m3_23944_21578# th_dif_sw_0.VCN 0.01078f
C8362 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_15472_21578# 0.03017f
C8363 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_n1472_21578# 0.0162f
C8364 c1_12980_21618# VCM 0.01358f
C8365 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP 0.21251f
C8366 c1_45456_46258# m3_45124_45098# 0.01078f
C8367 c1_n1140_45138# m3_n1472_45098# 1.74381f
C8368 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VCM 0.9961f
C8369 c1_45456_45138# m3_45124_46218# 0.01078f
C8370 sar10b_0.CF[6] sar10b_0.CF[7] 59.0076f
C8371 sar10b_0.CF[5] sar10b_0.CF[8] 0.11478f
C8372 sar10b_0.SWN[1] sar10b_0.CF[7] 0.13032f
C8373 a_61400_63620# a_61609_63602# 0.24088f
C8374 a_61395_63280# a_62185_63363# 0.1263f
C8375 sar10b_0._06_ sar10b_0.cyclic_flag_0.FINAL 0.15186f
C8376 m3_45124_82252# VDDR 0.01034f
C8377 m3_45124_78892# th_dif_sw_0.VCP 0.17339f
C8378 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN sar10b_0.SWP[3] 0.22728f
C8379 sar10b_0.net9 a_60945_60609# 0.05622f
C8380 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y 0.07183f
C8381 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 2.33263f
C8382 a_62133_59067# VSSD 0.13087f
C8383 a_62593_58639# a_62798_58688# 0.09983f
C8384 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN 0.01136f
C8385 c1_42632_97972# VCM 0.01358f
C8386 sar10b_0.clk_div_0.COUNT\[0\] sar10b_0.SWN[6] 0.23556f
C8387 m3_45124_67692# c1_45456_67732# 1.74381f
C8388 m3_n1472_67692# c1_n1140_66612# 0.01078f
C8389 m3_n1472_66572# c1_n1140_67732# 0.01078f
C8390 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VSSR 1.33794f
C8391 VSSR c1_45456_67732# 0.0935f
C8392 a_67209_64335# VSSD 0.51583f
C8393 sar10b_0.net14 VSSD 3.10641f
C8394 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A VDDR 0.38472f
C8395 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A 0.02842f
C8396 sar10b_0.net29 VSSD 0.59651f
C8397 sar10b_0.CF[6] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A 0.06369f
C8398 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A 0.39629f
C8399 m3_23944_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26603f
C8400 m3_32416_97932# m3_33828_97932# 0.23959f
C8401 sar10b_0.net44 sar10b_0.net45 2.47089f
C8402 a_66933_64395# a_67598_64016# 0.19065f
C8403 a_67209_64335# a_67733_64115# 0.04522f
C8404 a_62181_51440# a_62527_51646# 0.07649f
C8405 VSSD DATA[3] 0.61935f
C8406 sar10b_0.net45 a_66367_66298# 0.27333f
C8407 c1_n1140_84532# c1_n1140_83412# 0.13255f
C8408 m3_n1472_42858# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C8409 VDDD a_61400_52964# 0.24411f
C8410 VSSD a_60747_60609# 0.24593f
C8411 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP sar10b_0.CF[3] 0.10517f
C8412 c1_1684_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26825f
C8413 sar10b_0.net47 a_68946_71059# 0.24802f
C8414 m3_22532_97932# c1_21452_97972# 0.15596f
C8415 a_64809_65963# a_66021_66092# 0.07766f
C8416 VSSD a_62261_56123# 0.09871f
C8417 VSSR m3_n1472_32778# 0.66371f
C8418 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A sar10b_0.CF[8] 0.01887f
C8419 sar10b_0.net3 a_67733_65447# 0.16772f
C8420 sar10b_0.net46 a_68235_71265# 0.05736f
C8421 sar10b_0._03_ a_67611_50645# 0.01375f
C8422 sar10b_0.CF[6] sar10b_0.SWN[5] 0.11864f
C8423 c1_45456_48498# VDDR 0.01151f
C8424 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 1.37832f
C8425 a_64245_59307# a_64910_59686# 0.19065f
C8426 m3_45124_51818# th_dif_sw_0.VCN 0.17339f
C8427 a_68325_56296# VSSD 0.27209f
C8428 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 3.89075f
C8429 VSSR c1_41220_21618# 0.05923f
C8430 a_61395_60616# a_61086_60642# 0.07766f
C8431 sar10b_0.clk_div_0.COUNT\[0\] sar10b_0._03_ 0.17705f
C8432 a_65865_57675# a_66825_57675# 0.03471f
C8433 a_66049_57307# a_66254_57356# 0.09983f
C8434 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 0.02632f
C8435 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_n1140_21618# 0.0106f
C8436 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSSR 2.50986f
C8437 sar10b_0.SWP[2] a_34741_111361# 0.64048f
C8438 VSSR m3_n1472_73292# 0.66316f
C8439 c1_45456_49618# c1_45456_48498# 0.13255f
C8440 a_66255_50749# sar10b_0.net16 0.03306f
C8441 sar10b_0._04_ sar10b_0.net35 0.06792f
C8442 sar10b_0.net3 sar10b_0._12_ 0.1156f
C8443 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y 0.07183f
C8444 VSSD a_63457_56931# 0.8832f
C8445 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A 0.03718f
C8446 m3_n1472_24938# VCM 0.01415f
C8447 VDDD a_65865_57675# 0.75585f
C8448 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 1.78633f
C8449 c1_n1140_75572# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C8450 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A 0.95194f
C8451 m3_45124_50698# m3_45124_49578# 0.29566f
C8452 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP 0.02666f
C8453 a_62037_61731# a_62497_61303# 0.26257f
C8454 a_62313_61671# a_62702_61352# 0.05462f
C8455 VDDD DATA[8] 0.34536f
C8456 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] 1.04257f
C8457 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.10429f
C8458 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] 2.12897f
C8459 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.41496f
C8460 a_65861_51977# a_66865_52076# 0.06302f
C8461 sar10b_0.SWP[9] VSSD 1.51924f
C8462 sar10b_0.net23 a_68421_62956# 0.01476f
C8463 sar10b_0.CF[1] sar10b_0.CF[9] 0.10934f
C8464 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.02632f
C8465 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 2.55153f
C8466 sar10b_0._09_ a_64199_50761# 0.03351f
C8467 VDDD a_63573_63303# 0.28649f
C8468 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A 1.33999f
C8469 sar10b_0.CF[1] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 0.12389f
C8470 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y 0.32264f
C8471 sar10b_0.net1 a_61929_56639# 0.05596f
C8472 c1_25688_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] 0.26825f
C8473 m3_n1472_65452# VCM 0.01412f
C8474 a_65119_59984# sar10b_0.net33 0.27246f
C8475 VDDD a_65961_68627# 0.36631f
C8476 a_63849_63299# a_64238_63682# 0.06034f
C8477 a_64033_63591# a_64809_63299# 0.3578f
C8478 th_dif_sw_0.VCP sar10b_0.CF[3] 0.29827f
C8479 VDDR EN 0.07767f
C8480 sar10b_0.net2 a_61493_56924# 0.02733f
C8481 VDDD a_66961_50219# 0.41371f
C8482 c1_n1140_49618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C8483 a_63967_58652# sar10b_0.net39 0.05073f
C8484 a_67077_69616# sar10b_0.net16 0.17594f
C8485 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP sar10b_0.SWP[5] 0.24477f
C8486 VSSR c1_n1140_39538# 0.04956f
C8487 a_61065_51015# a_60789_51075# 0.1263f
C8488 a_16238_8706# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A 0.01076f
C8489 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A 1.11457f
C8490 sar10b_0.net16 sar10b_0.net1 5.5632f
C8491 m3_45124_82252# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C8492 sar10b_0.net40 a_61677_66174# 0.01034f
C8493 m3_45124_91212# m3_45124_90092# 0.29566f
C8494 VSSR m3_5588_97932# 0.54637f
C8495 m3_43712_21578# c1_44044_21618# 1.74381f
C8496 sar10b_0.net16 a_61086_61974# 0.17419f
C8497 m3_5588_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.53746f
C8498 sar10b_0.net10 VSSD 2.06065f
C8499 a_67372_52243# sar10b_0._07_ 0.09521f
C8500 a_63457_56931# sar10b_0.net31 0.16483f
C8501 a_64485_56768# a_64233_56639# 0.27388f
C8502 sar10b_0.net13 VSSD 3.11271f
C8503 a_62497_61303# a_62837_61451# 0.24088f
C8504 m3_45124_94572# c1_45456_95732# 0.01078f
C8505 m3_n1472_94572# c1_n1140_94612# 1.74381f
C8506 m3_45124_95692# c1_45456_94612# 0.01078f
C8507 sar10b_0.net16 a_61400_66284# 0.12467f
C8508 VSSR m3_31004_21578# 0.49843f
C8509 VSSD a_67598_65348# 0.13552f
C8510 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A 0.03718f
C8511 sar10b_0.net10 a_63561_60339# 0.22325f
C8512 VDDD a_66933_68391# 0.32463f
C8513 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A 0.41861f
C8514 c1_45456_54098# m3_45124_52938# 0.01078f
C8515 c1_45456_52978# m3_45124_54058# 0.01078f
C8516 sar10b_0.net18 sar10b_0.net36 1.26518f
C8517 sar10b_0.net21 sar10b_0.net19 1.04202f
C8518 c1_n1140_52978# m3_n1472_52938# 1.74381f
C8519 VSSD a_65198_66346# 0.13937f
C8520 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.24766f
C8521 VCM cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 0.12357f
C8522 m3_45124_97932# VDDR 0.01034f
C8523 m3_45124_94572# th_dif_sw_0.VCP 0.17339f
C8524 a_61677_50190# a_62185_50043# 0.19065f
C8525 sar10b_0.CF[5] sar10b_0.SWN[0] 0.12707f
C8526 m3_25356_97932# VCM 0.13579f
C8527 a_62185_52707# sar10b_0.net16 0.44229f
C8528 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 1.71649f
C8529 a_67564_50907# VSSD 0.20153f
C8530 a_68946_52411# VSSD 0.31355f
C8531 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.02632f
C8532 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 6.04723f
C8533 sar10b_0.net46 VSSD 1.7654f
C8534 a_67105_59971# sar10b_0.cyclic_flag_0.FINAL 0.08062f
C8535 sar10b_0.CF[7] a_60747_65563# 0.14263f
C8536 sar10b_0.clk_div_0.COUNT\[0\] a_66464_50363# 0.04617f
C8537 c1_3096_97972# VCM 0.01358f
C8538 m3_29592_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C8539 m3_45124_75532# c1_45456_75572# 1.74381f
C8540 m3_n1472_74412# c1_n1140_75572# 0.01078f
C8541 m3_n1472_75532# c1_n1140_74452# 0.01078f
C8542 VSSR c1_45456_83412# 0.0935f
C8543 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A 0.28117f
C8544 a_63391_57320# a_63273_56639# 0.01379f
C8545 sar10b_0.net38 a_61609_62270# 0.0226f
C8546 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[1] 0.05939f
C8547 VDDD sar10b_0.CF[9] 0.59626f
C8548 sar10b_0.cyclic_flag_0.FINAL a_66837_56403# 0.06527f
C8549 c1_7332_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C8550 sar10b_0.SWP[8] VCM 0.13076f
C8551 m3_12648_97932# m3_14060_97932# 0.23959f
C8552 sar10b_0.clknet_1_0__leaf_CLK a_65643_48621# 0.06254f
C8553 a_62497_61303# sar10b_0.net11 0.01613f
C8554 c1_n1140_92372# c1_n1140_91252# 0.13255f
C8555 c1_272_21618# m3_n60_21578# 1.74381f
C8556 sar10b_0.SWN[6] sar10b_0.SWN[7] 17.8422f
C8557 a_64521_59303# sar10b_0.net12 0.0147f
C8558 VDDD a_60969_56639# 0.87274f
C8559 VDDA sar10b_0.SWP[1] 0.2491f
C8560 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN 5.24097f
C8561 tdc_0.phase_detector_0.INN a_53564_59480# 0.01369f
C8562 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 0.80358f
C8563 sar10b_0.SWP[1] a_38665_107026# 0.96592f
C8564 m3_2764_97932# c1_1684_97972# 0.15596f
C8565 sar10b_0.net13 sar10b_0.CF[8] 0.03777f
C8566 VSSR m3_n1472_48458# 0.66371f
C8567 c1_31336_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.26825f
C8568 VSSD a_63525_61624# 0.27801f
C8569 a_67393_67963# a_68169_68331# 0.3578f
C8570 VDDD a_62187_71265# 0.29255f
C8571 sar10b_0.net16 a_66254_57356# 0.24882f
C8572 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VDDR 0.75888f
C8573 c1_45456_67732# VDDR 0.01153f
C8574 sar10b_0.net20 a_68946_52411# 0.25709f
C8575 m3_15472_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C8576 VSSD a_62997_67299# 0.15849f
C8577 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 0.21974f
C8578 m3_38064_21578# m3_39476_21578# 0.23959f
C8579 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A 0.60027f
C8580 VSSR c1_14392_21618# 0.05555f
C8581 a_64188_51135# sar10b_0._00_ 0.06207f
C8582 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VSSR 4.77284f
C8583 a_61833_57675# a_63045_57628# 0.07766f
C8584 a_62222_57356# a_62357_57455# 0.35559f
C8585 VDDA tdc_0.phase_detector_0.INN 0.49684f
C8586 VDDD a_68169_66999# 0.36668f
C8587 a_68946_68627# DATA[9] 0.1424f
C8588 a_65061_63428# sar10b_0.net16 0.17454f
C8589 VSSR m3_n1472_88972# 0.66316f
C8590 c1_45456_57458# c1_45456_56338# 0.13255f
C8591 VDDD sar10b_0._01_ 1.11894f
C8592 VDDD a_66645_61731# 0.33536f
C8593 m3_n1472_32778# VDDR 0.02681f
C8594 a_60789_51075# sar10b_0.net16 0.23192f
C8595 a_65573_52937# a_65928_53032# 0.18757f
C8596 m3_n1472_40618# VCM 0.01415f
C8597 c1_n1140_91252# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.15596f
C8598 a_65586_50645# VSSD 1.18439f
C8599 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.83558f
C8600 VSSR c1_44044_97972# 0.07152f
C8601 a_63509_62783# VSSD 0.10689f
C8602 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 0.21577f
C8603 sar10b_0.SWN[7] sar10b_0.CF[7] 2.47018f
C8604 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_36652_21578# 0.03017f
C8605 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_19708_21578# 0.0162f
C8606 a_64428_50947# VSSD 0.13902f
C8607 c1_21452_21618# VCM 0.01311f
C8608 sar10b_0.net24 sar10b_0.net22 0.03739f
C8609 sar10b_0.net29 sar10b_0.SWN[0] 0.26385f
C8610 VDDD a_65778_49979# 0.43295f
C8611 VDDA th_dif_sw_0.CK 4.44457f
C8612 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VDDR 3.26494f
C8613 m3_n1472_73292# VDDR 0.02674f
C8614 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 0.02638f
C8615 m3_n1472_81132# VCM 0.01412f
C8616 m3_23944_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] 0.18853f
C8617 sar10b_0._01_ sar10b_0._08_ 0.02438f
C8618 sar10b_0.SWN[1] EN 0.1386f
C8619 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y sar10b_0.CF[5] 0.12541f
C8620 a_64149_64635# sar10b_0.net2 0.23439f
C8621 c1_n1140_24978# c1_n1140_23858# 0.13255f
C8622 sar10b_0.net9 a_61400_62288# 0.05162f
C8623 VDDD a_61131_70891# 0.30376f
C8624 sar10b_0.net33 a_65643_48621# 0.24997f
C8625 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 4.61507f
C8626 a_67733_65447# a_68169_65667# 0.16939f
C8627 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VCM 0.13025f
C8628 m3_n1472_26058# m3_n1472_24938# 0.29566f
C8629 sar10b_0.cyclic_flag_0.FINAL sar10b_0.net45 0.42233f
C8630 sar10b_0.net18 sar10b_0._04_ 0.01348f
C8631 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38716f
C8632 VSSR c1_n1140_55218# 0.04956f
C8633 sar10b_0.SWN[6] sar10b_0.CF[7] 0.12122f
C8634 a_51345_60437# tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A 0.14814f
C8635 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C8636 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 a_5929_113881# 0.12755f
C8637 VDDD a_67209_55011# 0.92305f
C8638 sar10b_0.net34 sar10b_0.cyclic_flag_0.FINAL 0.09027f
C8639 a_60690_49683# EN 0.44045f
C8640 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 3.8907f
C8641 m3_21120_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] 0.1528f
C8642 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A 0.75806f
C8643 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y 0.3196f
C8644 m3_23944_21578# c1_24276_21618# 1.74381f
C8645 VDDD a_67372_52833# 0.25671f
C8646 m3_45124_35018# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C8647 VDDD a_68946_68627# 0.28022f
C8648 sar10b_0.CF[0] a_60747_56239# 0.14263f
C8649 a_61454_50696# CLK 0.01211f
C8650 a_61929_56639# a_62527_56974# 0.06623f
C8651 a_65589_69723# a_66049_69295# 0.26257f
C8652 a_65865_69663# a_66254_69344# 0.05462f
C8653 sar10b_0.SWN[4] VCM 0.13075f
C8654 m3_32416_97932# c1_32748_97972# 1.74381f
C8655 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.41436f
C8656 VSSR m3_45124_24938# 0.63261f
C8657 VSSD a_61395_61948# 0.50861f
C8658 a_60693_51315# a_61358_51694# 0.19065f
C8659 tdc_0.phase_detector_0.INN tdc_0.phase_detector_0.INP 1.21226f
C8660 c1_36984_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26825f
C8661 sar10b_0.SWP[5] sar10b_0.net43 0.06335f
C8662 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A 0.07183f
C8663 VSSD a_60945_65937# 0.28817f
C8664 a_67733_62783# a_68169_63003# 0.16939f
C8665 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A 0.95194f
C8666 sar10b_0.net4 sar10b_0.CF[1] 0.03914f
C8667 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.74815f
C8668 sar10b_0.net16 a_62527_56974# 0.04026f
C8669 tdc_0.phase_detector_0.INN tdc_0.phase_detector_0.pd_out_0.A 0.06563f
C8670 m3_n1472_66572# m3_n1472_65452# 0.29566f
C8671 a_34741_111361# cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 0.01247f
C8672 VSSR m3_45124_65452# 0.63305f
C8673 sar10b_0.CF[0] VCM 38.3953f
C8674 sar10b_0.net2 a_61395_60616# 0.01319f
C8675 sar10b_0.CF[2] sar10b_0.CF[9] 0.10127f
C8676 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN sar10b_0.SWN[8] 0.19451f
C8677 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A 0.28117f
C8678 a_61677_52854# VSSD 0.13077f
C8679 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN sar10b_0.CF[2] 0.10485f
C8680 sar10b_0.SWN[6] sar10b_0.SWN[5] 16.1081f
C8681 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSSR 0.36438f
C8682 m3_11236_21578# VCM 0.13579f
C8683 VDDD sar10b_0.net35 2.58704f
C8684 m3_n1472_83372# c1_n1140_82292# 0.01078f
C8685 m3_45124_83372# c1_45456_83412# 1.74381f
C8686 m3_n1472_82252# c1_n1140_83412# 0.01078f
C8687 VDDD a_63339_48621# 0.25196f
C8688 sar10b_0.clk_div_0.COUNT\[0\] sar10b_0._13_ 0.19185f
C8689 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 0.68971f
C8690 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] 7.81593f
C8691 VCM cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 6.31441f
C8692 sar10b_0.net3 a_67733_68111# 0.15088f
C8693 c1_n1140_29458# m3_n1472_28298# 0.01078f
C8694 c1_45456_29458# m3_45124_29418# 1.74381f
C8695 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 0.2477f
C8696 c1_n1140_28338# m3_n1472_29418# 0.01078f
C8697 VDDD a_61929_57971# 0.36004f
C8698 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 3.50557f
C8699 sar10b_0.SWP[8] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 0.37026f
C8700 a_66645_60399# sar10b_0.net3 0.21939f
C8701 VDDD a_63810_50901# 0.3855f
C8702 a_61496_52091# a_62281_52347# 0.26257f
C8703 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A 1.37577f
C8704 a_60969_57971# a_61493_58256# 0.05022f
C8705 a_64338_52411# sar10b_0.net16 0.03949f
C8706 sar10b_0._08_ sar10b_0.net35 0.01974f
C8707 c1_45456_83412# VDDR 0.01153f
C8708 m3_18296_21578# m3_19708_21578# 0.23959f
C8709 a_67310_61352# a_67445_61451# 0.35559f
C8710 VSSR c1_45456_31698# 0.09348f
C8711 sar10b_0.net4 a_61589_53459# 0.0549f
C8712 a_64667_51628# sar10b_0.net16 0.01055f
C8713 tdc_0.RDY sar10b_0.CF[0] 0.14969f
C8714 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 0.40988f
C8715 m3_n1472_73292# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C8716 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 3.70208f
C8717 a_61929_67295# sar10b_0.net40 0.02168f
C8718 sar10b_0.CF[4] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] 0.01357f
C8719 a_n8277_54249# VCM 0.06006f
C8720 sar10b_0.SWN[5] sar10b_0.CF[7] 0.12305f
C8721 VSSR m3_26768_97932# 0.44047f
C8722 c1_45456_68852# c1_45456_67732# 0.13255f
C8723 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VDDR 2.96384f
C8724 sar10b_0.cyclic_flag_0.FINAL sar10b_0.net36 0.04488f
C8725 VDDD a_62409_59007# 0.86457f
C8726 m3_26768_21578# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.26806f
C8727 m3_n1472_48458# VDDR 0.02681f
C8728 sar10b_0.net29 a_61419_48621# 0.02906f
C8729 m3_n1472_56298# VCM 0.01415f
C8730 a_61395_52624# a_61086_52650# 0.07766f
C8731 sar10b_0.net28 sar10b_0.net17 0.10739f
C8732 a_64033_63591# VSSD 0.91403f
C8733 sar10b_0._09_ a_64454_51311# 0.10808f
C8734 a_67209_59007# a_66933_59067# 0.1263f
C8735 VDDD a_60747_64231# 0.28486f
C8736 VDDD a_60747_69559# 0.28829f
C8737 th_dif_sw_0.VCP VINP 3.18189f
C8738 a_61153_67587# sar10b_0.net16 0.09786f
C8739 VDDD a_61395_49960# 0.77801f
C8740 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 0.24774f
C8741 VSSR c1_4508_97972# 0.05923f
C8742 w_n9655_63119# th_dif_sw_0.th_sw_1.CKB 0.23172f
C8743 a_65481_59303# sar10b_0.net16 0.326f
C8744 sar10b_0.clknet_0_CLK a_66666_51977# 0.02018f
C8745 VDDD sar10b_0.net4 2.78913f
C8746 sar10b_0.net2 a_62017_57307# 0.02903f
C8747 sar10b_0._17_ sar10b_0._16_ 0.01353f
C8748 a_68767_63980# sar10b_0.net25 0.02266f
C8749 a_63273_56639# a_63662_57022# 0.06034f
C8750 VSSR cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 41.7127f
C8751 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VDDR 5.56064f
C8752 a_63273_67295# a_64238_67295# 0.03279f
C8753 a_65865_69663# a_65961_68627# 0.02084f
C8754 m3_n1472_88972# VDDR 0.02674f
C8755 VDDD a_62126_56024# 0.26891f
C8756 m3_n1472_96812# VCM 0.01942f
C8757 sar10b_0.net40 a_66885_56768# 0.01088f
C8758 sar10b_0.net3 sar10b_0.net16 0.02081f
C8759 a_61358_51694# VSSD 0.12906f
C8760 a_68946_59303# VSSD 0.33361f
C8761 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A 0.42509f
C8762 c1_n1140_32818# c1_n1140_31698# 0.13255f
C8763 VSSA VCM 0.51555f
C8764 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN sar10b_0.SWP[7] 0.20154f
C8765 VDDD a_68073_56343# 0.36728f
C8766 a_65573_52937# a_66378_52993# 0.29207f
C8767 sar10b_0.net42 VSSD 2.71416f
C8768 sar10b_0.net28 a_61677_50190# 0.02841f
C8769 sar10b_0._03_ a_66464_50363# 0.0233f
C8770 c1_24276_97972# VCM 0.01358f
C8771 a_60945_63273# sar10b_0.net38 0.0131f
C8772 m3_n1472_33898# m3_n1472_32778# 0.29566f
C8773 sar10b_0.net3 a_67310_61352# 0.24012f
C8774 VSSR c1_n1140_74452# 0.04956f
C8775 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_2868_111642# 0.01076f
C8776 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A 1.11457f
C8777 m3_5588_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.53746f
C8778 c1_28512_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.0106f
C8779 a_67598_68012# VSSD 0.13567f
C8780 a_67209_59007# sar10b_0.net3 0.18208f
C8781 a_60969_67295# a_61153_67587# 0.44532f
C8782 c1_10156_21618# m3_11236_21578# 0.15596f
C8783 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A 0.41861f
C8784 m3_45124_50698# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.22792f
C8785 sar10b_0._14_ a_68178_51635# 0.10544f
C8786 a_65733_59432# a_65481_59303# 0.27388f
C8787 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A 0.03718f
C8788 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A 0.02842f
C8789 a_66921_60339# VSSD 0.51575f
C8790 m3_12648_97932# c1_12980_97972# 1.74381f
C8791 a_61153_51603# CLK 0.04116f
C8792 VSSR m3_45124_40618# 0.63261f
C8793 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP a_9853_5788# 0.07015f
C8794 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y sar10b_0.CF[4] 0.17717f
C8795 sar10b_0._10_ a_65068_49569# 0.09553f
C8796 c1_10156_21618# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.01541f
C8797 a_65765_50645# a_65996_50650# 0.08144f
C8798 a_66255_50749# a_66103_50668# 0.2328f
C8799 m3_36652_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] 0.0162f
C8800 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS th_dif_sw_0.th_sw_1.CK 0.22609f
C8801 VSSR c1_22864_21618# 0.05003f
C8802 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A sar10b_0.CF[2] 0.06369f
C8803 a_64609_64923# sar10b_0.net16 0.12678f
C8804 a_67084_53565# VSSD 0.15662f
C8805 a_67209_55011# a_68169_55011# 0.03529f
C8806 a_67393_54643# a_67598_54692# 0.09983f
C8807 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN 0.01175f
C8808 tdc_0.RDY VSSA 0.34723f
C8809 m3_n1472_74412# m3_n1472_73292# 0.29566f
C8810 sar10b_0.net33 sar10b_0.net12 0.0218f
C8811 VSSR m3_45124_81132# 0.63305f
C8812 VDDD a_67419_52937# 0.19467f
C8813 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 0.84046f
C8814 sar10b_0.net3 a_67393_54643# 0.11049f
C8815 sar10b_0.net38 a_66885_56768# 0.03017f
C8816 a_68946_63299# DATA[7] 0.14522f
C8817 sar10b_0._13_ sar10b_0.net37 0.88482f
C8818 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VCM 3.21926f
C8819 VDDR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.38864f
C8820 m3_45124_24938# VDDR 0.0103f
C8821 VSSD a_62181_56768# 0.26639f
C8822 VDDD a_61557_57735# 0.28784f
C8823 sar10b_0.SWP[0] sar10b_0.CF[3] 0.12401f
C8824 m3_n1472_91212# c1_n1140_90132# 0.01078f
C8825 m3_n1472_90092# c1_n1140_91252# 0.01078f
C8826 m3_45124_91212# c1_45456_91252# 1.74381f
C8827 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A 0.10815f
C8828 a_67733_62783# VSSD 0.10006f
C8829 VDDD a_68767_58652# 0.2137f
C8830 sar10b_0.net16 a_61086_64638# 0.18334f
C8831 m3_45124_57418# m3_45124_56298# 0.29566f
C8832 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_40888_21578# 0.0162f
C8833 sar10b_0.net16 a_66537_57971# 0.27846f
C8834 sar10b_0.net33 a_65573_52937# 0.0254f
C8835 c1_42632_21618# VCM 0.01358f
C8836 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 2.7512f
C8837 sar10b_0.CF[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN 0.07717f
C8838 c1_45456_37298# m3_45124_37258# 1.74381f
C8839 c1_n1140_37298# m3_n1472_36138# 0.01078f
C8840 c1_n1140_36178# m3_n1472_37258# 0.01078f
C8841 sar10b_0._09_ a_64188_51135# 0.01872f
C8842 VDDD a_62185_63363# 0.29064f
C8843 sar10b_0.SWN[7] EN 0.38739f
C8844 VSSR sar10b_0.CF[9] 25.4939f
C8845 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y a_31680_8700# 0.01076f
C8846 m3_45124_65452# VDDR 0.01034f
C8847 m3_45124_62092# th_dif_sw_0.VCP 0.34926f
C8848 VDDD a_64725_68631# 0.28578f
C8849 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 7.63271f
C8850 a_61419_71265# VSSD 0.34238f
C8851 a_62933_58787# sar10b_0.net16 0.13986f
C8852 a_63745_59971# a_64521_60339# 0.3578f
C8853 VDDD a_67393_65299# 0.25553f
C8854 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A sar10b_0.CF[1] 0.06369f
C8855 VSSD CKO 0.90878f
C8856 th_dif_sw_0.th_sw_1.CKB a_n8277_65767# 0.0331f
C8857 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VDDR 0.59881f
C8858 a_65673_56639# a_65857_56931# 0.44532f
C8859 th_dif_sw_0.CKB a_61035_48621# 0.12004f
C8860 a_67696_52265# a_67747_51991# 0.01442f
C8861 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A 0.42509f
C8862 sar10b_0.net7 a_62017_57307# 0.01713f
C8863 VSSD a_67105_61303# 0.85524f
C8864 VDDD sar10b_0.net44 1.4571f
C8865 a_65185_68919# a_66213_68756# 0.07826f
C8866 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VCM 0.12735f
C8867 VDDD a_66367_66298# 0.22141f
C8868 VDDD a_60789_53739# 0.33151f
C8869 m3_n1472_21578# m3_n60_21578# 0.23959f
C8870 a_65001_68627# a_65961_68627# 0.03432f
C8871 VSSR c1_45456_47378# 0.09348f
C8872 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A 0.42509f
C8873 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] 14.1554f
C8874 sar10b_0.net16 a_61086_60642# 0.17376f
C8875 VDDD sar10b_0.net18 1.20288f
C8876 m3_n1472_88972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.24158f
C8877 sar10b_0.SWN[6] EN 0.25349f
C8878 a_65957_50273# a_66312_50368# 0.18757f
C8879 sar10b_0.net28 a_60690_49683# 0.01515f
C8880 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A 0.11547f
C8881 sar10b_0.clk_div_0.COUNT\[0\] sar10b_0.clknet_1_0__leaf_CLK 0.15275f
C8882 c1_45456_76692# c1_45456_75572# 0.13255f
C8883 a_65577_51311# VSSD 2.2036f
C8884 sar10b_0.net16 a_62949_56296# 0.17491f
C8885 VDDD a_69003_71265# 0.26713f
C8886 sar10b_0.net34 a_66368_49417# 0.01335f
C8887 m3_35240_21578# c1_34160_21618# 0.15596f
C8888 m3_n1472_26058# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C8889 sar10b_0.net3 a_67696_52265# 0.0214f
C8890 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VDDR 0.83994f
C8891 a_1127_5779# VSSR 0.4375f
C8892 sar10b_0.net38 a_61609_64934# 0.0226f
C8893 a_64245_59307# sar10b_0.net11 0.03948f
C8894 a_67077_69616# a_67423_69308# 0.07649f
C8895 c1_44044_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.01078f
C8896 sar10b_0.net3 sar10b_0.clk_div_0.COUNT\[1\] 0.13628f
C8897 sar10b_0.net34 a_65761_58263# 0.02743f
C8898 m3_43712_97932# c1_42632_97972# 0.15596f
C8899 VSSD sar10b_0.net8 1.95974f
C8900 VSSR m3_12648_21578# 0.49843f
C8901 a_55121_59650# VDDA 0.22342f
C8902 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP sar10b_0.CF[5] 0.10502f
C8903 c1_45456_31698# VDDR 0.01151f
C8904 m3_45124_35018# th_dif_sw_0.VCN 0.17339f
C8905 a_65045_59588# VSSD 0.10257f
C8906 a_55282_59893# tdc_0.phase_detector_0.pd_out_0.B 0.01666f
C8907 sar10b_0.net18 sar10b_0._08_ 0.01869f
C8908 sar10b_0.net14 a_61929_67295# 0.01289f
C8909 m3_7000_97932# VCM 0.15231f
C8910 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] c1_28512_21618# 0.0106f
C8911 VDDD a_63273_61671# 0.35949f
C8912 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 0.01239f
C8913 sar10b_0.net4 a_62527_67630# 0.05787f
C8914 a_60693_67299# a_61358_67678# 0.19065f
C8915 c1_n1140_40658# c1_n1140_39538# 0.13255f
C8916 VDDD sar10b_0.SWP[2] 1.61241f
C8917 VDDD a_63273_67295# 0.87242f
C8918 a_61395_61948# a_61609_62270# 0.04522f
C8919 a_61086_61974# a_61400_62288# 0.07826f
C8920 sar10b_0.net39 a_62997_56643# 0.01689f
C8921 a_67142_68689# VSSD 0.01178f
C8922 m3_32416_21578# VCM 0.13579f
C8923 m3_11236_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 0.03017f
C8924 m3_n1472_41738# m3_n1472_40618# 0.29566f
C8925 sar10b_0.net38 a_61609_60938# 0.02142f
C8926 VSSR c1_n1140_90132# 0.04956f
C8927 sar10b_0._13_ sar10b_0._03_ 0.02837f
C8928 tdc_0.OUTP VDDA 0.42203f
C8929 a_24259_5788# cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 0.60421f
C8930 VDDR cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] 9.88107f
C8931 a_67393_63967# sar10b_0.net3 0.1307f
C8932 VSSR cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A 1.10847f
C8933 a_63950_60020# VSSD 0.18203f
C8934 VSSD a_65673_56639# 0.49715f
C8935 a_64425_64631# a_64949_64916# 0.05022f
C8936 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A 0.26364f
C8937 sar10b_0.net40 a_63045_57628# 0.04523f
C8938 a_67696_52265# a_67798_52206# 0.15528f
C8939 a_63745_59971# a_63285_60399# 0.26257f
C8940 a_63950_60020# a_63561_60339# 0.05462f
C8941 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 2.76344f
C8942 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] 14.1554f
C8943 sar10b_0.net33 sar10b_0.net41 0.14461f
C8944 a_67372_52243# sar10b_0.clk_div_0.COUNT\[2\] 0.0428f
C8945 a_66027_53575# VSSD 0.33245f
C8946 VDDD a_63374_62684# 0.26028f
C8947 VSSR m3_45124_56298# 0.6325f
C8948 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A 0.04073f
C8949 VCM th_dif_sw_0.VCN 2.83149f
C8950 c1_n1140_32818# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.15596f
C8951 VDDD a_64199_50761# 0.85101f
C8952 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 0.02632f
C8953 sar10b_0.net33 sar10b_0.clk_div_0.COUNT\[0\] 0.02515f
C8954 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A 0.95194f
C8955 sar10b_0.net42 a_64492_67433# 0.02184f
C8956 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A 0.28117f
C8957 VSSR c1_n1140_22738# 0.04956f
C8958 sar10b_0.SWP[5] VCM 0.13076f
C8959 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSSR 4.4718f
C8960 VDDD sar10b_0._11_ 0.20552f
C8961 sar10b_0.CF[6] cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A 0.01887f
C8962 m3_45124_65452# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.22792f
C8963 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP a_25137_112201# 0.01111f
C8964 VSSA w_n9655_63119# 4.20223f
C8965 m3_n1472_82252# m3_n1472_81132# 0.29566f
C8966 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A sar10b_0.CF[0] 0.03041f
C8967 VSSR m3_45124_96812# 0.63305f
C8968 a_64425_64631# VSSD 0.58328f
C8969 a_64780_52239# a_64924_52385# 0.2119f
C8970 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VSSR 1.37482f
C8971 m3_45124_40618# VDDR 0.0103f
C8972 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A sar10b_0.CF[2] 0.05939f
C8973 sar10b_0.SWN[5] EN 0.19974f
C8974 sar10b_0.net9 VSSD 2.39929f
C8975 a_67372_52243# VSSD 0.43309f
C8976 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y 0.07183f
C8977 VDDD sar10b_0.net23 0.91724f
C8978 a_65385_64631# sar10b_0.net14 0.01658f
C8979 a_61395_64612# a_61400_64952# 0.44098f
C8980 a_60945_64605# a_61086_64638# 0.27388f
C8981 VSSR c1_25688_97972# 0.05451f
C8982 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 0.01239f
C8983 a_64543_62648# sar10b_0.net42 0.29032f
C8984 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A 1.29717f
C8985 sar10b_0.SWN[4] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN 0.22176f
C8986 a_66789_58100# a_66537_57971# 0.27388f
C8987 sar10b_0.CF[4] sar10b_0.SWN[2] 0.12162f
C8988 m3_26768_21578# th_dif_sw_0.VCN 0.01078f
C8989 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] m3_18296_21578# 0.03017f
C8990 a_65301_57975# sar10b_0.net14 0.01941f
C8991 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] m3_1352_21578# 0.0162f
C8992 a_55121_59650# tdc_0.phase_detector_0.pd_out_0.A 0.09615f
C8993 a_66216_49358# VSSD 0.11861f
C8994 c1_15804_21618# VCM 0.01358f
C8995 c1_n1140_44018# m3_n1472_45098# 0.01078f
C8996 c1_n1140_45138# m3_n1472_43978# 0.01078f
C8997 c1_45456_45138# m3_45124_45098# 1.74381f
C8998 VSSD a_61395_64612# 0.51698f
C8999 sar10b_0.net12 a_65865_57675# 0.22361f
C9000 m3_45124_81132# VDDR 0.01034f
C9001 m3_45124_77772# th_dif_sw_0.VCP 0.17339f
C9002 VSSD a_66101_58256# 0.09962f
C9003 VSSR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A 1.12023f
C9004 VDDD a_60747_61941# 0.22504f
C9005 sar10b_0.net9 a_61400_60956# 0.19593f
C9006 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A 0.68875f
C9007 a_62593_58639# VSSD 0.85157f
C9008 a_62798_58688# a_62933_58787# 0.35559f
C9009 a_62409_59007# a_63621_58960# 0.07766f
C9010 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSSR 33.417f
C9011 c1_45456_97972# VCM 0.02046f
C9012 m3_45124_66572# c1_45456_67732# 0.01078f
C9013 m3_45124_67692# c1_45456_66612# 0.01078f
C9014 m3_n1472_66572# c1_n1140_66612# 1.74381f
C9015 th_dif_sw_0.CK a_n4470_65264# 0.69236f
C9016 VSSR c1_45456_66612# 0.0935f
C9017 sar10b_0.net32 sar10b_0.clknet_1_1__leaf_CLK 0.09495f
C9018 tdc_0.OUTP tdc_0.phase_detector_0.pd_out_0.A 0.25963f
C9019 VDDR sar10b_0.CF[9] 1.96206f
C9020 m3_26768_97932# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26806f
C9021 m3_33828_97932# m3_35240_97932# 0.23959f
C9022 a_67393_63967# a_67598_64016# 0.09983f
C9023 a_61929_51311# sar10b_0.net28 0.03748f
C9024 VDDR cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN 4.58095f
C9025 c1_45456_84532# c1_45456_83412# 0.13255f
C9026 c1_45456_22738# m3_45124_21578# 0.01078f
C9027 VDDD a_61609_52946# 0.20857f
C9028 m3_n1472_41738# cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] 0.24158f
C9029 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN 2.12902f
C9030 sar10b_0.net4 tdc_0.OUTN 0.27011f
C9031 c1_4508_97972# cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] 0.26825f
C9032 sar10b_0.net21 VSSD 0.9203f
C9033 m3_23944_97932# c1_22864_97972# 0.15596f
C9034 a_64993_66255# a_66021_66092# 0.07826f
C9035 a_64533_65967# a_65198_66346# 0.19065f
C9036 DATA[0] VSUBS 0.32243f
C9037 DATA[1] VSUBS 0.24591f
C9038 EN VSUBS 52.1026f
C9039 DATA[2] VSUBS 0.24591f
C9040 DATA[3] VSUBS 0.24606f
C9041 DATA[4] VSUBS 0.25018f
C9042 DATA[5] VSUBS 0.28478f
C9043 VINN VSUBS 6.40269f
C9044 DATA[6] VSUBS 0.26478f
C9045 CLK VSUBS 14.2148f
C9046 DATA[7] VSUBS 0.26596f
C9047 VINP VSUBS 6.40267f
C9048 DATA[8] VSUBS 0.27426f
C9049 DATA[9] VSUBS 0.27818f
C9050 CKO VSUBS 0.30123f
C9051 VCM VSUBS 40.4602f
C9052 VSSD VSUBS 66.43021f
C9053 VSSA VSUBS 0.10406p
C9054 VSSR VSUBS 0.10351p
C9055 VDDD VSUBS 1.09863p
C9056 VDDR VSUBS 18.2562p
C9057 VDDA VSUBS 0.75978p
C9058 c1_45456_21618# VSUBS 0.10766f $ **FLOATING
C9059 c1_44044_21618# VSUBS 0.05383f $ **FLOATING
C9060 c1_42632_21618# VSUBS 0.05383f $ **FLOATING
C9061 c1_41220_21618# VSUBS 0.05383f $ **FLOATING
C9062 c1_39808_21618# VSUBS 0.05383f $ **FLOATING
C9063 c1_38396_21618# VSUBS 0.05383f $ **FLOATING
C9064 c1_36984_21618# VSUBS 0.05383f $ **FLOATING
C9065 c1_35572_21618# VSUBS 0.05383f $ **FLOATING
C9066 c1_34160_21618# VSUBS 0.05383f $ **FLOATING
C9067 c1_32748_21618# VSUBS 0.05383f $ **FLOATING
C9068 c1_31336_21618# VSUBS 0.05383f $ **FLOATING
C9069 c1_29924_21618# VSUBS 0.05383f $ **FLOATING
C9070 c1_28512_21618# VSUBS 0.05383f $ **FLOATING
C9071 c1_27100_21618# VSUBS 0.05383f $ **FLOATING
C9072 c1_25688_21618# VSUBS 0.05383f $ **FLOATING
C9073 c1_24276_21618# VSUBS 0.05383f $ **FLOATING
C9074 c1_22864_21618# VSUBS 0.05383f $ **FLOATING
C9075 c1_21452_21618# VSUBS 0.05383f $ **FLOATING
C9076 c1_20040_21618# VSUBS 0.05383f $ **FLOATING
C9077 c1_18628_21618# VSUBS 0.05383f $ **FLOATING
C9078 c1_17216_21618# VSUBS 0.05383f $ **FLOATING
C9079 c1_15804_21618# VSUBS 0.05383f $ **FLOATING
C9080 c1_14392_21618# VSUBS 0.05383f $ **FLOATING
C9081 c1_12980_21618# VSUBS 0.05383f $ **FLOATING
C9082 c1_11568_21618# VSUBS 0.05383f $ **FLOATING
C9083 c1_10156_21618# VSUBS 0.05383f $ **FLOATING
C9084 c1_8744_21618# VSUBS 0.05383f $ **FLOATING
C9085 c1_7332_21618# VSUBS 0.05383f $ **FLOATING
C9086 c1_5920_21618# VSUBS 0.05383f $ **FLOATING
C9087 c1_4508_21618# VSUBS 0.05383f $ **FLOATING
C9088 c1_3096_21618# VSUBS 0.05383f $ **FLOATING
C9089 c1_1684_21618# VSUBS 0.05383f $ **FLOATING
C9090 c1_272_21618# VSUBS 0.05383f $ **FLOATING
C9091 c1_n1140_21618# VSUBS 0.05383f $ **FLOATING
C9092 c1_45456_22738# VSUBS 0.05383f $ **FLOATING
C9093 c1_45456_23858# VSUBS 0.05383f $ **FLOATING
C9094 c1_45456_24978# VSUBS 0.05383f $ **FLOATING
C9095 c1_45456_26098# VSUBS 0.05383f $ **FLOATING
C9096 c1_45456_27218# VSUBS 0.05383f $ **FLOATING
C9097 c1_45456_28338# VSUBS 0.05383f $ **FLOATING
C9098 c1_45456_29458# VSUBS 0.05383f $ **FLOATING
C9099 c1_45456_30578# VSUBS 0.05383f $ **FLOATING
C9100 c1_45456_31698# VSUBS 0.05383f $ **FLOATING
C9101 c1_45456_32818# VSUBS 0.05383f $ **FLOATING
C9102 c1_45456_33938# VSUBS 0.05383f $ **FLOATING
C9103 c1_45456_35058# VSUBS 0.05383f $ **FLOATING
C9104 c1_45456_36178# VSUBS 0.05383f $ **FLOATING
C9105 c1_45456_37298# VSUBS 0.05383f $ **FLOATING
C9106 c1_45456_38418# VSUBS 0.05383f $ **FLOATING
C9107 c1_45456_39538# VSUBS 0.05383f $ **FLOATING
C9108 c1_45456_40658# VSUBS 0.05383f $ **FLOATING
C9109 c1_45456_41778# VSUBS 0.05383f $ **FLOATING
C9110 c1_45456_42898# VSUBS 0.05383f $ **FLOATING
C9111 c1_45456_44018# VSUBS 0.05383f $ **FLOATING
C9112 c1_45456_45138# VSUBS 0.05383f $ **FLOATING
C9113 c1_45456_46258# VSUBS 0.05383f $ **FLOATING
C9114 c1_45456_47378# VSUBS 0.05383f $ **FLOATING
C9115 c1_45456_48498# VSUBS 0.05383f $ **FLOATING
C9116 c1_45456_49618# VSUBS 0.05383f $ **FLOATING
C9117 c1_45456_50738# VSUBS 0.05383f $ **FLOATING
C9118 c1_45456_51858# VSUBS 0.05383f $ **FLOATING
C9119 c1_45456_52978# VSUBS 0.05383f $ **FLOATING
C9120 c1_45456_54098# VSUBS 0.05383f $ **FLOATING
C9121 c1_45456_55218# VSUBS 0.05383f $ **FLOATING
C9122 c1_45456_56338# VSUBS 0.05383f $ **FLOATING
C9123 c1_45456_57458# VSUBS 0.10766f $ **FLOATING
C9124 c1_n1140_57458# VSUBS 0.05383f $ **FLOATING
C9125 c1_45456_62132# VSUBS 0.10766f $ **FLOATING
C9126 c1_n1140_62132# VSUBS 0.05383f $ **FLOATING
C9127 c1_45456_63252# VSUBS 0.05383f $ **FLOATING
C9128 c1_45456_64372# VSUBS 0.05383f $ **FLOATING
C9129 c1_45456_65492# VSUBS 0.05383f $ **FLOATING
C9130 c1_45456_66612# VSUBS 0.05383f $ **FLOATING
C9131 c1_45456_67732# VSUBS 0.05383f $ **FLOATING
C9132 c1_45456_68852# VSUBS 0.05383f $ **FLOATING
C9133 c1_45456_69972# VSUBS 0.05383f $ **FLOATING
C9134 c1_45456_71092# VSUBS 0.05383f $ **FLOATING
C9135 c1_45456_72212# VSUBS 0.05383f $ **FLOATING
C9136 c1_45456_73332# VSUBS 0.05383f $ **FLOATING
C9137 c1_45456_74452# VSUBS 0.05383f $ **FLOATING
C9138 c1_45456_75572# VSUBS 0.05383f $ **FLOATING
C9139 c1_45456_76692# VSUBS 0.05383f $ **FLOATING
C9140 c1_45456_77812# VSUBS 0.05383f $ **FLOATING
C9141 c1_45456_78932# VSUBS 0.05383f $ **FLOATING
C9142 c1_45456_80052# VSUBS 0.05383f $ **FLOATING
C9143 c1_45456_81172# VSUBS 0.05383f $ **FLOATING
C9144 c1_45456_82292# VSUBS 0.05383f $ **FLOATING
C9145 c1_45456_83412# VSUBS 0.05383f $ **FLOATING
C9146 c1_45456_84532# VSUBS 0.05383f $ **FLOATING
C9147 c1_45456_85652# VSUBS 0.05383f $ **FLOATING
C9148 c1_45456_86772# VSUBS 0.05383f $ **FLOATING
C9149 c1_45456_87892# VSUBS 0.05383f $ **FLOATING
C9150 c1_45456_89012# VSUBS 0.05383f $ **FLOATING
C9151 c1_45456_90132# VSUBS 0.05383f $ **FLOATING
C9152 c1_45456_91252# VSUBS 0.05383f $ **FLOATING
C9153 c1_45456_92372# VSUBS 0.05383f $ **FLOATING
C9154 c1_45456_93492# VSUBS 0.05383f $ **FLOATING
C9155 c1_45456_94612# VSUBS 0.05383f $ **FLOATING
C9156 c1_45456_95732# VSUBS 0.05383f $ **FLOATING
C9157 c1_45456_96852# VSUBS 0.05383f $ **FLOATING
C9158 c1_45456_97972# VSUBS 0.10766f $ **FLOATING
C9159 c1_44044_97972# VSUBS 0.05383f $ **FLOATING
C9160 c1_42632_97972# VSUBS 0.05383f $ **FLOATING
C9161 c1_41220_97972# VSUBS 0.05383f $ **FLOATING
C9162 c1_39808_97972# VSUBS 0.05383f $ **FLOATING
C9163 c1_38396_97972# VSUBS 0.05383f $ **FLOATING
C9164 c1_36984_97972# VSUBS 0.05383f $ **FLOATING
C9165 c1_35572_97972# VSUBS 0.05383f $ **FLOATING
C9166 c1_34160_97972# VSUBS 0.05383f $ **FLOATING
C9167 c1_32748_97972# VSUBS 0.05383f $ **FLOATING
C9168 c1_31336_97972# VSUBS 0.05383f $ **FLOATING
C9169 c1_29924_97972# VSUBS 0.05383f $ **FLOATING
C9170 c1_28512_97972# VSUBS 0.05383f $ **FLOATING
C9171 c1_27100_97972# VSUBS 0.05383f $ **FLOATING
C9172 c1_25688_97972# VSUBS 0.05383f $ **FLOATING
C9173 c1_24276_97972# VSUBS 0.05383f $ **FLOATING
C9174 c1_22864_97972# VSUBS 0.05383f $ **FLOATING
C9175 c1_21452_97972# VSUBS 0.05383f $ **FLOATING
C9176 c1_20040_97972# VSUBS 0.05383f $ **FLOATING
C9177 c1_18628_97972# VSUBS 0.05383f $ **FLOATING
C9178 c1_17216_97972# VSUBS 0.05383f $ **FLOATING
C9179 c1_15804_97972# VSUBS 0.05383f $ **FLOATING
C9180 c1_14392_97972# VSUBS 0.05383f $ **FLOATING
C9181 c1_12980_97972# VSUBS 0.05383f $ **FLOATING
C9182 c1_11568_97972# VSUBS 0.05383f $ **FLOATING
C9183 c1_10156_97972# VSUBS 0.05383f $ **FLOATING
C9184 c1_8744_97972# VSUBS 0.05383f $ **FLOATING
C9185 c1_7332_97972# VSUBS 0.05383f $ **FLOATING
C9186 c1_5920_97972# VSUBS 0.05383f $ **FLOATING
C9187 c1_4508_97972# VSUBS 0.05383f $ **FLOATING
C9188 c1_3096_97972# VSUBS 0.05383f $ **FLOATING
C9189 c1_1684_97972# VSUBS 0.05383f $ **FLOATING
C9190 c1_272_97972# VSUBS 0.05383f $ **FLOATING
C9191 c1_n1140_97972# VSUBS 0.05383f $ **FLOATING
C9192 m3_45124_21578# VSUBS 0.14242f $ **FLOATING
C9193 m3_43712_21578# VSUBS 0.0787f $ **FLOATING
C9194 m3_42300_21578# VSUBS 0.0787f $ **FLOATING
C9195 m3_40888_21578# VSUBS 0.0787f $ **FLOATING
C9196 m3_39476_21578# VSUBS 0.0787f $ **FLOATING
C9197 m3_38064_21578# VSUBS 0.0787f $ **FLOATING
C9198 m3_36652_21578# VSUBS 0.0787f $ **FLOATING
C9199 m3_35240_21578# VSUBS 0.0787f $ **FLOATING
C9200 m3_33828_21578# VSUBS 0.0787f $ **FLOATING
C9201 m3_32416_21578# VSUBS 0.0787f $ **FLOATING
C9202 m3_31004_21578# VSUBS 0.0787f $ **FLOATING
C9203 m3_29592_21578# VSUBS 0.0787f $ **FLOATING
C9204 m3_28180_21578# VSUBS 0.0787f $ **FLOATING
C9205 m3_26768_21578# VSUBS 0.0787f $ **FLOATING
C9206 m3_25356_21578# VSUBS 0.0787f $ **FLOATING
C9207 m3_23944_21578# VSUBS 0.0787f $ **FLOATING
C9208 m3_22532_21578# VSUBS 0.0787f $ **FLOATING
C9209 m3_21120_21578# VSUBS 0.0787f $ **FLOATING
C9210 m3_19708_21578# VSUBS 0.0787f $ **FLOATING
C9211 m3_18296_21578# VSUBS 0.0787f $ **FLOATING
C9212 m3_16884_21578# VSUBS 0.0787f $ **FLOATING
C9213 m3_15472_21578# VSUBS 0.0787f $ **FLOATING
C9214 m3_14060_21578# VSUBS 0.0787f $ **FLOATING
C9215 m3_12648_21578# VSUBS 0.0787f $ **FLOATING
C9216 m3_11236_21578# VSUBS 0.0787f $ **FLOATING
C9217 m3_9824_21578# VSUBS 0.0787f $ **FLOATING
C9218 m3_8412_21578# VSUBS 0.0787f $ **FLOATING
C9219 m3_7000_21578# VSUBS 0.0787f $ **FLOATING
C9220 m3_5588_21578# VSUBS 0.0787f $ **FLOATING
C9221 m3_4176_21578# VSUBS 0.0787f $ **FLOATING
C9222 m3_2764_21578# VSUBS 0.0787f $ **FLOATING
C9223 m3_1352_21578# VSUBS 0.0787f $ **FLOATING
C9224 m3_n60_21578# VSUBS 0.0787f $ **FLOATING
C9225 m3_n1472_21578# VSUBS 0.25459f $ **FLOATING
C9226 m3_45124_22698# VSUBS 0.06371f $ **FLOATING
C9227 m3_n1472_22698# VSUBS 0.17588f $ **FLOATING
C9228 m3_45124_23818# VSUBS 0.06371f $ **FLOATING
C9229 m3_n1472_23818# VSUBS 0.17588f $ **FLOATING
C9230 m3_45124_24938# VSUBS 0.06371f $ **FLOATING
C9231 m3_n1472_24938# VSUBS 0.17588f $ **FLOATING
C9232 m3_45124_26058# VSUBS 0.06371f $ **FLOATING
C9233 m3_n1472_26058# VSUBS 0.17588f $ **FLOATING
C9234 m3_45124_27178# VSUBS 0.06371f $ **FLOATING
C9235 m3_n1472_27178# VSUBS 0.17588f $ **FLOATING
C9236 m3_45124_28298# VSUBS 0.06371f $ **FLOATING
C9237 m3_n1472_28298# VSUBS 0.17588f $ **FLOATING
C9238 m3_45124_29418# VSUBS 0.06371f $ **FLOATING
C9239 m3_n1472_29418# VSUBS 0.17588f $ **FLOATING
C9240 m3_45124_30538# VSUBS 0.06371f $ **FLOATING
C9241 m3_n1472_30538# VSUBS 0.17588f $ **FLOATING
C9242 m3_45124_31658# VSUBS 0.06371f $ **FLOATING
C9243 m3_n1472_31658# VSUBS 0.17588f $ **FLOATING
C9244 m3_45124_32778# VSUBS 0.06371f $ **FLOATING
C9245 m3_n1472_32778# VSUBS 0.17588f $ **FLOATING
C9246 m3_45124_33898# VSUBS 0.06371f $ **FLOATING
C9247 m3_n1472_33898# VSUBS 0.17588f $ **FLOATING
C9248 m3_45124_35018# VSUBS 0.06371f $ **FLOATING
C9249 m3_n1472_35018# VSUBS 0.17588f $ **FLOATING
C9250 m3_45124_36138# VSUBS 0.06371f $ **FLOATING
C9251 m3_n1472_36138# VSUBS 0.17588f $ **FLOATING
C9252 m3_45124_37258# VSUBS 0.06371f $ **FLOATING
C9253 m3_n1472_37258# VSUBS 0.17588f $ **FLOATING
C9254 m3_45124_38378# VSUBS 0.06371f $ **FLOATING
C9255 m3_n1472_38378# VSUBS 0.17588f $ **FLOATING
C9256 m3_45124_39498# VSUBS 0.06371f $ **FLOATING
C9257 m3_n1472_39498# VSUBS 0.17588f $ **FLOATING
C9258 m3_45124_40618# VSUBS 0.06371f $ **FLOATING
C9259 m3_n1472_40618# VSUBS 0.17588f $ **FLOATING
C9260 m3_45124_41738# VSUBS 0.06371f $ **FLOATING
C9261 m3_n1472_41738# VSUBS 0.17588f $ **FLOATING
C9262 m3_45124_42858# VSUBS 0.06371f $ **FLOATING
C9263 m3_n1472_42858# VSUBS 0.17473f $ **FLOATING
C9264 m3_45124_43978# VSUBS 0.06371f $ **FLOATING
C9265 m3_n1472_43978# VSUBS 0.17588f $ **FLOATING
C9266 m3_45124_45098# VSUBS 0.06371f $ **FLOATING
C9267 m3_n1472_45098# VSUBS 0.17588f $ **FLOATING
C9268 m3_45124_46218# VSUBS 0.06371f $ **FLOATING
C9269 m3_n1472_46218# VSUBS 0.17588f $ **FLOATING
C9270 m3_45124_47338# VSUBS 0.06371f $ **FLOATING
C9271 m3_n1472_47338# VSUBS 0.17588f $ **FLOATING
C9272 m3_45124_48458# VSUBS 0.06371f $ **FLOATING
C9273 m3_n1472_48458# VSUBS 0.17588f $ **FLOATING
C9274 m3_45124_49578# VSUBS 0.06371f $ **FLOATING
C9275 m3_n1472_49578# VSUBS 0.17588f $ **FLOATING
C9276 m3_45124_50698# VSUBS 0.06371f $ **FLOATING
C9277 m3_n1472_50698# VSUBS 0.17588f $ **FLOATING
C9278 m3_45124_51818# VSUBS 0.06371f $ **FLOATING
C9279 m3_n1472_51818# VSUBS 0.17588f $ **FLOATING
C9280 m3_45124_52938# VSUBS 0.06371f $ **FLOATING
C9281 m3_n1472_52938# VSUBS 0.17588f $ **FLOATING
C9282 m3_45124_54058# VSUBS 0.06371f $ **FLOATING
C9283 m3_n1472_54058# VSUBS 0.17588f $ **FLOATING
C9284 m3_45124_55178# VSUBS 0.05578f $ **FLOATING
C9285 m3_n1472_55178# VSUBS 0.17588f $ **FLOATING
C9286 m3_45124_56298# VSUBS 0.06298f $ **FLOATING
C9287 m3_n1472_56298# VSUBS 0.17588f $ **FLOATING
C9288 m3_45124_57418# VSUBS 0.12654f $ **FLOATING
C9289 m3_n1472_57418# VSUBS 0.25459f $ **FLOATING
C9290 m3_45124_62092# VSUBS 0.14242f $ **FLOATING
C9291 m3_n1472_62092# VSUBS 0.25459f $ **FLOATING
C9292 m3_45124_63212# VSUBS 0.06371f $ **FLOATING
C9293 m3_n1472_63212# VSUBS 0.17588f $ **FLOATING
C9294 m3_45124_64332# VSUBS 0.06371f $ **FLOATING
C9295 m3_n1472_64332# VSUBS 0.17588f $ **FLOATING
C9296 m3_45124_65452# VSUBS 0.06371f $ **FLOATING
C9297 m3_n1472_65452# VSUBS 0.17588f $ **FLOATING
C9298 m3_45124_66572# VSUBS 0.06371f $ **FLOATING
C9299 m3_n1472_66572# VSUBS 0.17588f $ **FLOATING
C9300 m3_45124_67692# VSUBS 0.06371f $ **FLOATING
C9301 m3_n1472_67692# VSUBS 0.17588f $ **FLOATING
C9302 m3_45124_68812# VSUBS 0.06371f $ **FLOATING
C9303 m3_n1472_68812# VSUBS 0.17588f $ **FLOATING
C9304 m3_45124_69932# VSUBS 0.06371f $ **FLOATING
C9305 m3_n1472_69932# VSUBS 0.17588f $ **FLOATING
C9306 m3_45124_71052# VSUBS 0.06371f $ **FLOATING
C9307 m3_n1472_71052# VSUBS 0.17588f $ **FLOATING
C9308 m3_45124_72172# VSUBS 0.06371f $ **FLOATING
C9309 m3_n1472_72172# VSUBS 0.17588f $ **FLOATING
C9310 m3_45124_73292# VSUBS 0.06371f $ **FLOATING
C9311 m3_n1472_73292# VSUBS 0.17588f $ **FLOATING
C9312 m3_45124_74412# VSUBS 0.06371f $ **FLOATING
C9313 m3_n1472_74412# VSUBS 0.17588f $ **FLOATING
C9314 m3_45124_75532# VSUBS 0.06371f $ **FLOATING
C9315 m3_n1472_75532# VSUBS 0.17588f $ **FLOATING
C9316 m3_45124_76652# VSUBS 0.06371f $ **FLOATING
C9317 m3_n1472_76652# VSUBS 0.17588f $ **FLOATING
C9318 m3_45124_77772# VSUBS 0.06371f $ **FLOATING
C9319 m3_n1472_77772# VSUBS 0.17588f $ **FLOATING
C9320 m3_45124_78892# VSUBS 0.06371f $ **FLOATING
C9321 m3_n1472_78892# VSUBS 0.17588f $ **FLOATING
C9322 m3_45124_80012# VSUBS 0.06371f $ **FLOATING
C9323 m3_n1472_80012# VSUBS 0.17588f $ **FLOATING
C9324 m3_45124_81132# VSUBS 0.06371f $ **FLOATING
C9325 m3_n1472_81132# VSUBS 0.17588f $ **FLOATING
C9326 m3_45124_82252# VSUBS 0.06371f $ **FLOATING
C9327 m3_n1472_82252# VSUBS 0.17588f $ **FLOATING
C9328 m3_45124_83372# VSUBS 0.06371f $ **FLOATING
C9329 m3_n1472_83372# VSUBS 0.17588f $ **FLOATING
C9330 m3_45124_84492# VSUBS 0.06371f $ **FLOATING
C9331 m3_n1472_84492# VSUBS 0.17588f $ **FLOATING
C9332 m3_45124_85612# VSUBS 0.06371f $ **FLOATING
C9333 m3_n1472_85612# VSUBS 0.17588f $ **FLOATING
C9334 m3_45124_86732# VSUBS 0.06371f $ **FLOATING
C9335 m3_n1472_86732# VSUBS 0.17588f $ **FLOATING
C9336 m3_45124_87852# VSUBS 0.06371f $ **FLOATING
C9337 m3_n1472_87852# VSUBS 0.17588f $ **FLOATING
C9338 m3_45124_88972# VSUBS 0.06371f $ **FLOATING
C9339 m3_n1472_88972# VSUBS 0.17588f $ **FLOATING
C9340 m3_45124_90092# VSUBS 0.06371f $ **FLOATING
C9341 m3_n1472_90092# VSUBS 0.17588f $ **FLOATING
C9342 m3_45124_91212# VSUBS 0.06371f $ **FLOATING
C9343 m3_n1472_91212# VSUBS 0.17588f $ **FLOATING
C9344 m3_45124_92332# VSUBS 0.06371f $ **FLOATING
C9345 m3_n1472_92332# VSUBS 0.17588f $ **FLOATING
C9346 m3_45124_93452# VSUBS 0.06371f $ **FLOATING
C9347 m3_n1472_93452# VSUBS 0.17588f $ **FLOATING
C9348 m3_45124_94572# VSUBS 0.06371f $ **FLOATING
C9349 m3_n1472_94572# VSUBS 0.17588f $ **FLOATING
C9350 m3_45124_95692# VSUBS 0.06371f $ **FLOATING
C9351 m3_n1472_95692# VSUBS 0.17588f $ **FLOATING
C9352 m3_45124_96812# VSUBS 0.06371f $ **FLOATING
C9353 m3_n1472_96812# VSUBS 0.17588f $ **FLOATING
C9354 m3_45124_97932# VSUBS 0.14242f $ **FLOATING
C9355 m3_43712_97932# VSUBS 0.0787f $ **FLOATING
C9356 m3_42300_97932# VSUBS 0.0787f $ **FLOATING
C9357 m3_40888_97932# VSUBS 0.0787f $ **FLOATING
C9358 m3_39476_97932# VSUBS 0.0787f $ **FLOATING
C9359 m3_38064_97932# VSUBS 0.0787f $ **FLOATING
C9360 m3_36652_97932# VSUBS 0.0787f $ **FLOATING
C9361 m3_35240_97932# VSUBS 0.0787f $ **FLOATING
C9362 m3_33828_97932# VSUBS 0.0787f $ **FLOATING
C9363 m3_32416_97932# VSUBS 0.0787f $ **FLOATING
C9364 m3_31004_97932# VSUBS 0.0787f $ **FLOATING
C9365 m3_29592_97932# VSUBS 0.0787f $ **FLOATING
C9366 m3_28180_97932# VSUBS 0.0787f $ **FLOATING
C9367 m3_26768_97932# VSUBS 0.0787f $ **FLOATING
C9368 m3_25356_97932# VSUBS 0.0787f $ **FLOATING
C9369 m3_23944_97932# VSUBS 0.0787f $ **FLOATING
C9370 m3_22532_97932# VSUBS 0.0787f $ **FLOATING
C9371 m3_21120_97932# VSUBS 0.0787f $ **FLOATING
C9372 m3_19708_97932# VSUBS 0.0787f $ **FLOATING
C9373 m3_18296_97932# VSUBS 0.0787f $ **FLOATING
C9374 m3_16884_97932# VSUBS 0.0787f $ **FLOATING
C9375 m3_15472_97932# VSUBS 0.0787f $ **FLOATING
C9376 m3_14060_97932# VSUBS 0.0787f $ **FLOATING
C9377 m3_12648_97932# VSUBS 0.0787f $ **FLOATING
C9378 m3_11236_97932# VSUBS 0.0787f $ **FLOATING
C9379 m3_9824_97932# VSUBS 0.0787f $ **FLOATING
C9380 m3_8412_97932# VSUBS 0.0787f $ **FLOATING
C9381 m3_7000_97932# VSUBS 0.0787f $ **FLOATING
C9382 m3_5588_97932# VSUBS 0.0787f $ **FLOATING
C9383 m3_4176_97932# VSUBS 0.0787f $ **FLOATING
C9384 m3_2764_97932# VSUBS 0.0787f $ **FLOATING
C9385 m3_1352_97932# VSUBS 0.0787f $ **FLOATING
C9386 m3_n60_97932# VSUBS 0.0787f $ **FLOATING
C9387 m3_n1472_97932# VSUBS 0.25459f $ **FLOATING
C9388 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27932f $ **FLOATING
C9389 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VSUBS 0.27476f $ **FLOATING
C9390 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03496f $ **FLOATING
C9391 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A VSUBS 0.034f $ **FLOATING
C9392 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VSUBS 0.21343f $ **FLOATING
C9393 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A VSUBS 0.22255f $ **FLOATING
C9394 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A VSUBS 0.05619f $ **FLOATING
C9395 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06692f $ **FLOATING
C9396 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y VSUBS 0.035f $ **FLOATING
C9397 a_44345_5779# VSUBS 0.22209f $ **FLOATING
C9398 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VSUBS 1.32788f $ **FLOATING
C9399 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSUBS 1.7619f $ **FLOATING
C9400 a_43467_5788# VSUBS 0.76225f $ **FLOATING
C9401 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSUBS 4.42803f $ **FLOATING
C9402 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27474f $ **FLOATING
C9403 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VSUBS 0.27476f $ **FLOATING
C9404 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03399f $ **FLOATING
C9405 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A VSUBS 0.034f $ **FLOATING
C9406 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VSUBS 0.21745f $ **FLOATING
C9407 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A VSUBS 0.25929f $ **FLOATING
C9408 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A VSUBS 0.05619f $ **FLOATING
C9409 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06826f $ **FLOATING
C9410 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y VSUBS 0.035f $ **FLOATING
C9411 a_39543_5779# VSUBS 0.20157f $ **FLOATING
C9412 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VSUBS 1.20219f $ **FLOATING
C9413 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[0] VSUBS 6.81604f $ **FLOATING
C9414 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VSUBS 5.81794f $ **FLOATING
C9415 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSUBS 1.61954f $ **FLOATING
C9416 a_38665_5788# VSUBS 0.68771f $ **FLOATING
C9417 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSUBS 4.0344f $ **FLOATING
C9418 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27473f $ **FLOATING
C9419 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VSUBS 0.27476f $ **FLOATING
C9420 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03399f $ **FLOATING
C9421 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VSUBS 0.034f $ **FLOATING
C9422 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VSUBS 0.21745f $ **FLOATING
C9423 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VSUBS 0.25929f $ **FLOATING
C9424 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VSUBS 0.05619f $ **FLOATING
C9425 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06825f $ **FLOATING
C9426 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VSUBS 0.035f $ **FLOATING
C9427 a_34741_5779# VSUBS 0.18104f $ **FLOATING
C9428 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VSUBS 1.07669f $ **FLOATING
C9429 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[1] VSUBS 3.66021f $ **FLOATING
C9430 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VSUBS 5.31109f $ **FLOATING
C9431 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSUBS 1.47906f $ **FLOATING
C9432 a_33863_5788# VSUBS 0.61316f $ **FLOATING
C9433 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSUBS 3.64064f $ **FLOATING
C9434 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27473f $ **FLOATING
C9435 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VSUBS 0.27476f $ **FLOATING
C9436 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03399f $ **FLOATING
C9437 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A VSUBS 0.034f $ **FLOATING
C9438 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A VSUBS 0.21745f $ **FLOATING
C9439 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A VSUBS 0.25929f $ **FLOATING
C9440 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A VSUBS 0.05619f $ **FLOATING
C9441 a_29939_5779# VSUBS 0.16052f $ **FLOATING
C9442 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VSUBS 0.95119f $ **FLOATING
C9443 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06825f $ **FLOATING
C9444 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y VSUBS 0.03532f $ **FLOATING
C9445 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[2] VSUBS 2.98506f $ **FLOATING
C9446 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VSUBS 4.74711f $ **FLOATING
C9447 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSUBS 1.33814f $ **FLOATING
C9448 a_29061_5788# VSUBS 0.53862f $ **FLOATING
C9449 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSUBS 3.2299f $ **FLOATING
C9450 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27473f $ **FLOATING
C9451 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSUBS 0.27476f $ **FLOATING
C9452 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03399f $ **FLOATING
C9453 a_25137_5779# VSUBS 0.13999f $ **FLOATING
C9454 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VSUBS 0.8257f $ **FLOATING
C9455 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A VSUBS 0.034f $ **FLOATING
C9456 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VSUBS 0.21745f $ **FLOATING
C9457 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VSUBS 0.25984f $ **FLOATING
C9458 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A VSUBS 0.05733f $ **FLOATING
C9459 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06825f $ **FLOATING
C9460 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[3] VSUBS 2.52477f $ **FLOATING
C9461 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VSUBS 4.16406f $ **FLOATING
C9462 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y VSUBS 0.03532f $ **FLOATING
C9463 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSUBS 1.19734f $ **FLOATING
C9464 a_24259_5788# VSUBS 0.46408f $ **FLOATING
C9465 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSUBS 2.83779f $ **FLOATING
C9466 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27473f $ **FLOATING
C9467 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSUBS 0.27476f $ **FLOATING
C9468 a_20335_5779# VSUBS 0.11946f $ **FLOATING
C9469 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VSUBS 0.7002f $ **FLOATING
C9470 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03399f $ **FLOATING
C9471 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A VSUBS 0.03496f $ **FLOATING
C9472 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[4] VSUBS 2.90183f $ **FLOATING
C9473 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VSUBS 3.59994f $ **FLOATING
C9474 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VSUBS 0.21778f $ **FLOATING
C9475 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VSUBS 0.25984f $ **FLOATING
C9476 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A VSUBS 0.05733f $ **FLOATING
C9477 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06906f $ **FLOATING
C9478 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y VSUBS 0.03532f $ **FLOATING
C9479 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSUBS 1.05711f $ **FLOATING
C9480 a_19457_5788# VSUBS 0.38954f $ **FLOATING
C9481 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSUBS 2.44511f $ **FLOATING
C9482 a_15533_5779# VSUBS 0.09894f $ **FLOATING
C9483 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VSUBS 0.5747f $ **FLOATING
C9484 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27473f $ **FLOATING
C9485 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSUBS 0.27476f $ **FLOATING
C9486 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[5] VSUBS 3.19494f $ **FLOATING
C9487 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VSUBS 3.03543f $ **FLOATING
C9488 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03426f $ **FLOATING
C9489 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A VSUBS 0.03496f $ **FLOATING
C9490 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VSUBS 0.21915f $ **FLOATING
C9491 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VSUBS 0.25984f $ **FLOATING
C9492 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A VSUBS 0.05733f $ **FLOATING
C9493 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06883f $ **FLOATING
C9494 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y VSUBS 0.03532f $ **FLOATING
C9495 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSUBS 0.91675f $ **FLOATING
C9496 a_14655_5788# VSUBS 0.315f $ **FLOATING
C9497 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSUBS 2.05302f $ **FLOATING
C9498 a_10731_5779# VSUBS 0.07841f $ **FLOATING
C9499 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VSUBS 0.44921f $ **FLOATING
C9500 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[6] VSUBS 3.14107f $ **FLOATING
C9501 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VSUBS 2.47087f $ **FLOATING
C9502 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27473f $ **FLOATING
C9503 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSUBS 0.27589f $ **FLOATING
C9504 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03402f $ **FLOATING
C9505 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A VSUBS 0.03496f $ **FLOATING
C9506 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSUBS 0.77702f $ **FLOATING
C9507 a_9853_5788# VSUBS 0.24046f $ **FLOATING
C9508 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VSUBS 0.21907f $ **FLOATING
C9509 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VSUBS 0.26082f $ **FLOATING
C9510 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A VSUBS 0.05733f $ **FLOATING
C9511 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06891f $ **FLOATING
C9512 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y VSUBS 0.03563f $ **FLOATING
C9513 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSUBS 1.66106f $ **FLOATING
C9514 a_5929_5779# VSUBS 0.05789f $ **FLOATING
C9515 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VSUBS 0.32373f $ **FLOATING
C9516 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[7] VSUBS 1.97347f $ **FLOATING
C9517 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VSUBS 1.90639f $ **FLOATING
C9518 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSUBS 0.63619f $ **FLOATING
C9519 a_5051_5788# VSUBS 0.16592f $ **FLOATING
C9520 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27588f $ **FLOATING
C9521 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSUBS 0.27719f $ **FLOATING
C9522 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.0341f $ **FLOATING
C9523 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A VSUBS 0.03496f $ **FLOATING
C9524 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSUBS 1.26925f $ **FLOATING
C9525 a_1127_5779# VSUBS 0.03736f $ **FLOATING
C9526 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VSUBS 0.19828f $ **FLOATING
C9527 a_249_5788# VSUBS 0.09138f $ **FLOATING
C9528 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VSUBS 0.2195f $ **FLOATING
C9529 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VSUBS 0.2605f $ **FLOATING
C9530 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[8] VSUBS 1.84658f $ **FLOATING
C9531 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VSUBS 1.36596f $ **FLOATING
C9532 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSUBS 0.49731f $ **FLOATING
C9533 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSUBS 0.88064f $ **FLOATING
C9534 cdac_0.single_10b_cdac_0.x10b_cap_array_0.SW[9] VSUBS 1.7415f $ **FLOATING
C9535 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VSUBS 0.98503f $ **FLOATING
C9536 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27603f $ **FLOATING
C9537 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VSUBS 0.27884f $ **FLOATING
C9538 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03402f $ **FLOATING
C9539 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A VSUBS 0.03496f $ **FLOATING
C9540 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VSUBS 0.21886f $ **FLOATING
C9541 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A VSUBS 0.05733f $ **FLOATING
C9542 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06899f $ **FLOATING
C9543 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A VSUBS 0.21523f $ **FLOATING
C9544 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A VSUBS 0.05733f $ **FLOATING
C9545 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06854f $ **FLOATING
C9546 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y VSUBS 0.03563f $ **FLOATING
C9547 cdac_0.single_10b_cdac_0.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y VSUBS 0.03563f $ **FLOATING
C9548 sar10b_0.SWN[8] VSUBS 24.4587f $ **FLOATING
C9549 sar10b_0.SWN[7] VSUBS 23.6179f $ **FLOATING
C9550 a_69003_48621# VSUBS 0.03406f $ **FLOATING
C9551 a_68562_48647# VSUBS 0.03406f $ **FLOATING
C9552 a_68235_48621# VSUBS 0.03496f $ **FLOATING
C9553 sar10b_0.SWN[5] VSUBS 22.2287f $ **FLOATING
C9554 a_66153_48647# VSUBS 0.53978f $ **FLOATING
C9555 a_65643_48621# VSUBS 0.03451f $ **FLOATING
C9556 sar10b_0.SWN[4] VSUBS 21.5234f $ **FLOATING
C9557 sar10b_0.SWN[3] VSUBS 20.7636f $ **FLOATING
C9558 a_64491_48621# VSUBS 0.03488f $ **FLOATING
C9559 a_63339_48621# VSUBS 0.03496f $ **FLOATING
C9560 sar10b_0.SWN[2] VSUBS 19.9498f $ **FLOATING
C9561 sar10b_0.SWN[0] VSUBS 22.256f $ **FLOATING
C9562 sar10b_0.SWN[1] VSUBS 19.0511f $ **FLOATING
C9563 a_62187_48621# VSUBS 0.03406f $ **FLOATING
C9564 a_61803_48621# VSUBS 0.03414f $ **FLOATING
C9565 a_61419_48621# VSUBS 0.03406f $ **FLOATING
C9566 a_61035_48621# VSUBS 0.03418f $ **FLOATING
C9567 sar10b_0.SWN[9] VSUBS 30.9711f $ **FLOATING
C9568 sar10b_0.SWN[6] VSUBS 22.8996f $ **FLOATING
C9569 a_68946_49747# VSUBS 0.03339f $ **FLOATING
C9570 a_68562_49747# VSUBS 0.03316f $ **FLOATING
C9571 a_67371_49579# VSUBS 0.03324f $ **FLOATING
C9572 a_66865_49412# VSUBS 0.07182f $ **FLOATING
C9573 a_66666_49313# VSUBS 0.03633f $ **FLOATING
C9574 a_66216_49358# VSUBS 0.03353f $ **FLOATING
C9575 a_66368_49417# VSUBS 0.03539f $ **FLOATING
C9576 a_65861_49313# VSUBS 0.07145f $ **FLOATING
C9577 a_65682_49313# VSUBS 0.10132f $ **FLOATING
C9578 a_65068_49569# VSUBS 0.03544f $ **FLOATING
C9579 a_60690_49683# VSUBS 0.27723f $ **FLOATING
C9580 a_66762_50329# VSUBS 0.03599f $ **FLOATING
C9581 a_67439_50041# VSUBS 0.03364f $ **FLOATING
C9582 a_66961_50219# VSUBS 0.07124f $ **FLOATING
C9583 a_66312_50368# VSUBS 0.03334f $ **FLOATING
C9584 a_66464_50363# VSUBS 0.03518f $ **FLOATING
C9585 a_65957_50273# VSUBS 0.07118f $ **FLOATING
C9586 sar10b_0._02_ VSUBS 0.05751f $ **FLOATING
C9587 a_65778_49979# VSUBS 0.10136f $ **FLOATING
C9588 a_65021_50292# VSUBS 0.03623f $ **FLOATING
C9589 a_61677_50190# VSUBS 0.0363f $ **FLOATING
C9590 a_61609_50282# VSUBS 0.03316f $ **FLOATING
C9591 a_61400_50300# VSUBS 0.06971f $ **FLOATING
C9592 a_61086_49986# VSUBS 0.03316f $ **FLOATING
C9593 a_60945_49953# VSUBS 0.06951f $ **FLOATING
C9594 sar10b_0.net29 VSUBS 0.10507f $ **FLOATING
C9595 a_61395_49960# VSUBS 0.10306f $ **FLOATING
C9596 a_60747_49953# VSUBS 0.03657f $ **FLOATING
C9597 sar10b_0._12_ VSUBS 0.05275f $ **FLOATING
C9598 a_67564_50907# VSUBS 0.03316f $ **FLOATING
C9599 a_66785_50875# VSUBS 0.17026f $ **FLOATING
C9600 a_66593_50645# VSUBS 0.0526f $ **FLOATING
C9601 a_66103_50668# VSUBS 0.03394f $ **FLOATING
C9602 a_66255_50749# VSUBS 0.03664f $ **FLOATING
C9603 a_65765_50645# VSUBS 0.06946f $ **FLOATING
C9604 a_65586_50645# VSUBS 0.09961f $ **FLOATING
C9605 sar10b_0.clknet_1_0__leaf_CLK VSUBS 0.15537f $ **FLOATING
C9606 sar10b_0._00_ VSUBS 0.0557f $ **FLOATING
C9607 a_64356_51029# VSUBS 0.03576f $ **FLOATING
C9608 a_64428_50947# VSUBS 0.03476f $ **FLOATING
C9609 a_64199_50761# VSUBS 0.07267f $ **FLOATING
C9610 sar10b_0.net17 VSUBS 0.1112f $ **FLOATING
C9611 sar10b_0.net30 VSUBS 0.0674f $ **FLOATING
C9612 a_64188_51135# VSUBS 0.10447f $ **FLOATING
C9613 a_63918_50969# VSUBS 0.03655f $ **FLOATING
C9614 a_63810_50901# VSUBS 0.07251f $ **FLOATING
C9615 a_62623_50660# VSUBS 0.0379f $ **FLOATING
C9616 a_62277_50968# VSUBS 0.03316f $ **FLOATING
C9617 a_62025_51015# VSUBS 0.06924f $ **FLOATING
C9618 a_61589_50795# VSUBS 0.03316f $ **FLOATING
C9619 a_61454_50696# VSUBS 0.03547f $ **FLOATING
C9620 a_61249_50647# VSUBS 0.06885f $ **FLOATING
C9621 a_61065_51015# VSUBS 0.10173f $ **FLOATING
C9622 sar10b_0._15_ VSUBS 0.05492f $ **FLOATING
C9623 a_68178_51635# VSUBS 0.03413f $ **FLOATING
C9624 a_65577_51311# VSUBS 0.52669f $ **FLOATING
C9625 a_64454_51311# VSUBS 0.03366f $ **FLOATING
C9626 a_64339_51661# VSUBS 0.03406f $ **FLOATING
C9627 sar10b_0._08_ VSUBS 0.12597f $ **FLOATING
C9628 a_61358_51694# VSUBS 0.03547f $ **FLOATING
C9629 sar10b_0.net28 VSUBS 0.0655f $ **FLOATING
C9630 a_62527_51646# VSUBS 0.03633f $ **FLOATING
C9631 a_61929_51311# VSUBS 0.07013f $ **FLOATING
C9632 a_62181_51440# VSUBS 0.03316f $ **FLOATING
C9633 a_61493_51596# VSUBS 0.03316f $ **FLOATING
C9634 a_61153_51603# VSUBS 0.06885f $ **FLOATING
C9635 a_60969_51311# VSUBS 0.10223f $ **FLOATING
C9636 sar10b_0._03_ VSUBS 0.05066f $ **FLOATING
C9637 sar10b_0._07_ VSUBS 0.14335f $ **FLOATING
C9638 a_68946_52411# VSUBS 0.03387f $ **FLOATING
C9639 sar10b_0._13_ VSUBS 0.06311f $ **FLOATING
C9640 a_68331_52243# VSUBS 0.03454f $ **FLOATING
C9641 sar10b_0.clk_div_0.COUNT\[2\] VSUBS 0.13557f $ **FLOATING
C9642 a_67798_52206# VSUBS 0.03527f $ **FLOATING
C9643 a_67696_52265# VSUBS 0.03332f $ **FLOATING
C9644 sar10b_0.clk_div_0.COUNT\[0\] VSUBS 0.28492f $ **FLOATING
C9645 sar10b_0.clk_div_0.COUNT\[1\] VSUBS 0.2112f $ **FLOATING
C9646 a_67372_52243# VSUBS 0.03594f $ **FLOATING
C9647 a_66865_52076# VSUBS 0.07181f $ **FLOATING
C9648 a_66666_51977# VSUBS 0.03627f $ **FLOATING
C9649 a_66216_52022# VSUBS 0.03316f $ **FLOATING
C9650 a_66368_52081# VSUBS 0.03513f $ **FLOATING
C9651 sar10b_0._04_ VSUBS 0.05021f $ **FLOATING
C9652 a_65861_51977# VSUBS 0.07095f $ **FLOATING
C9653 a_65682_51977# VSUBS 0.10156f $ **FLOATING
C9654 a_64924_52385# VSUBS 0.03582f $ **FLOATING
C9655 sar10b_0._01_ VSUBS 0.0568f $ **FLOATING
C9656 sar10b_0._09_ VSUBS 0.08976f $ **FLOATING
C9657 a_64780_52239# VSUBS 0.04275f $ **FLOATING
C9658 a_64338_52411# VSUBS 0.03406f $ **FLOATING
C9659 sar10b_0._11_ VSUBS 0.0379f $ **FLOATING
C9660 a_61705_51992# VSUBS 0.03316f $ **FLOATING
C9661 a_61773_52237# VSUBS 0.03547f $ **FLOATING
C9662 a_61496_52091# VSUBS 0.06885f $ **FLOATING
C9663 a_61491_52222# VSUBS 0.10226f $ **FLOATING
C9664 a_61182_52404# VSUBS 0.03316f $ **FLOATING
C9665 a_61041_52340# VSUBS 0.06926f $ **FLOATING
C9666 a_60843_52216# VSUBS 0.03633f $ **FLOATING
C9667 a_66378_52993# VSUBS 0.03657f $ **FLOATING
C9668 sar10b_0.clk_div_0.COUNT\[3\] VSUBS 0.12893f $ **FLOATING
C9669 sar10b_0._14_ VSUBS 0.12052f $ **FLOATING
C9670 a_67372_52833# VSUBS 0.03316f $ **FLOATING
C9671 a_66577_52883# VSUBS 0.07144f $ **FLOATING
C9672 a_65928_53032# VSUBS 0.03334f $ **FLOATING
C9673 a_66080_53027# VSUBS 0.03518f $ **FLOATING
C9674 a_65573_52937# VSUBS 0.07173f $ **FLOATING
C9675 a_65394_52643# VSUBS 0.11047f $ **FLOATING
C9676 a_61677_52854# VSUBS 0.03547f $ **FLOATING
C9677 a_61609_52946# VSUBS 0.03316f $ **FLOATING
C9678 a_61400_52964# VSUBS 0.06885f $ **FLOATING
C9679 a_61086_52650# VSUBS 0.03316f $ **FLOATING
C9680 a_60945_52617# VSUBS 0.06867f $ **FLOATING
C9681 a_61395_52624# VSUBS 0.10236f $ **FLOATING
C9682 a_60747_52617# VSUBS 0.03683f $ **FLOATING
C9683 sar10b_0._16_ VSUBS 0.05717f $ **FLOATING
C9684 a_67084_53565# VSUBS 0.03957f $ **FLOATING
C9685 sar10b_0._10_ VSUBS 0.13857f $ **FLOATING
C9686 sar10b_0._05_ VSUBS 0.06019f $ **FLOATING
C9687 sar10b_0._17_ VSUBS 0.03878f $ **FLOATING
C9688 a_66027_53575# VSUBS 0.03328f $ **FLOATING
C9689 a_62623_53324# VSUBS 0.04067f $ **FLOATING
C9690 a_62277_53632# VSUBS 0.03334f $ **FLOATING
C9691 a_62025_53679# VSUBS 0.0719f $ **FLOATING
C9692 a_61589_53459# VSUBS 0.03393f $ **FLOATING
C9693 a_61454_53360# VSUBS 0.03682f $ **FLOATING
C9694 a_61249_53311# VSUBS 0.07163f $ **FLOATING
C9695 th_dif_sw_0.CKB VSUBS 8.54518f $ **FLOATING
C9696 a_61065_53679# VSUBS 0.10639f $ **FLOATING
C9697 a_68946_53975# VSUBS 0.03602f $ **FLOATING
C9698 sar10b_0.clknet_1_1__leaf_CLK VSUBS 0.16854f $ **FLOATING
C9699 sar10b_0.clknet_0_CLK VSUBS 0.31015f $ **FLOATING
C9700 a_65355_53949# VSUBS 0.54399f $ **FLOATING
C9701 a_60690_53975# VSUBS 0.13669f $ **FLOATING
C9702 sar10b_0.net18 VSUBS 0.09033f $ **FLOATING
C9703 a_68767_54656# VSUBS 0.03836f $ **FLOATING
C9704 a_68421_54964# VSUBS 0.03395f $ **FLOATING
C9705 a_68169_55011# VSUBS 0.07098f $ **FLOATING
C9706 a_67733_54791# VSUBS 0.03316f $ **FLOATING
C9707 a_67598_54692# VSUBS 0.03547f $ **FLOATING
C9708 a_67393_54643# VSUBS 0.06991f $ **FLOATING
C9709 a_n8277_54565# VSUBS 0.44235f $ **FLOATING
C9710 a_67209_55011# VSUBS 0.11026f $ **FLOATING
C9711 a_n8277_54249# VSUBS 5.11409f $ **FLOATING
C9712 a_n4470_53722# VSUBS 0.6386f $ **FLOATING
C9713 a_60690_54641# VSUBS 0.07927f $ **FLOATING
C9714 sar10b_0.net20 VSUBS 0.05523f $ **FLOATING
C9715 a_68671_55988# VSUBS 0.03838f $ **FLOATING
C9716 a_68325_56296# VSUBS 0.03397f $ **FLOATING
C9717 a_68073_56343# VSUBS 0.07133f $ **FLOATING
C9718 a_67637_56123# VSUBS 0.03316f $ **FLOATING
C9719 a_67502_56024# VSUBS 0.03682f $ **FLOATING
C9720 a_67297_55975# VSUBS 0.07059f $ **FLOATING
C9721 a_67113_56343# VSUBS 0.10389f $ **FLOATING
C9722 a_63295_55988# VSUBS 0.04048f $ **FLOATING
C9723 a_62949_56296# VSUBS 0.03393f $ **FLOATING
C9724 a_62697_56343# VSUBS 0.07186f $ **FLOATING
C9725 a_62261_56123# VSUBS 0.03316f $ **FLOATING
C9726 a_62126_56024# VSUBS 0.03547f $ **FLOATING
C9727 a_61921_55975# VSUBS 0.06966f $ **FLOATING
C9728 a_61737_56343# VSUBS 0.10971f $ **FLOATING
C9729 a_60747_56239# VSUBS 0.03365f $ **FLOATING
C9730 a_68946_56639# VSUBS 0.03338f $ **FLOATING
C9731 a_66062_57022# VSUBS 0.03547f $ **FLOATING
C9732 sar10b_0.net37 VSUBS 0.06445f $ **FLOATING
C9733 a_67231_56974# VSUBS 0.03633f $ **FLOATING
C9734 a_66633_56639# VSUBS 0.06974f $ **FLOATING
C9735 a_66885_56768# VSUBS 0.03344f $ **FLOATING
C9736 a_66197_56924# VSUBS 0.03393f $ **FLOATING
C9737 a_65857_56931# VSUBS 0.07143f $ **FLOATING
C9738 a_65673_56639# VSUBS 0.10563f $ **FLOATING
C9739 a_63662_57022# VSUBS 0.03682f $ **FLOATING
C9740 sar10b_0.net31 VSUBS 0.06923f $ **FLOATING
C9741 a_64831_56974# VSUBS 0.04017f $ **FLOATING
C9742 a_64233_56639# VSUBS 0.07213f $ **FLOATING
C9743 a_64485_56768# VSUBS 0.03453f $ **FLOATING
C9744 a_63797_56924# VSUBS 0.03393f $ **FLOATING
C9745 a_63457_56931# VSUBS 0.07243f $ **FLOATING
C9746 a_63273_56639# VSUBS 0.11013f $ **FLOATING
C9747 a_61358_57022# VSUBS 0.03613f $ **FLOATING
C9748 a_62527_56974# VSUBS 0.03633f $ **FLOATING
C9749 a_61929_56639# VSUBS 0.06746f $ **FLOATING
C9750 a_62181_56768# VSUBS 0.03316f $ **FLOATING
C9751 a_61493_56924# VSUBS 0.03336f $ **FLOATING
C9752 a_61153_56931# VSUBS 0.06984f $ **FLOATING
C9753 a_60969_56639# VSUBS 0.10266f $ **FLOATING
C9754 sar10b_0.net5 VSUBS 0.29241f $ **FLOATING
C9755 sar10b_0.net35 VSUBS 0.1031f $ **FLOATING
C9756 a_67423_57320# VSUBS 0.03853f $ **FLOATING
C9757 a_67077_57628# VSUBS 0.03316f $ **FLOATING
C9758 a_66825_57675# VSUBS 0.06954f $ **FLOATING
C9759 a_66389_57455# VSUBS 0.03316f $ **FLOATING
C9760 a_66254_57356# VSUBS 0.03553f $ **FLOATING
C9761 a_66049_57307# VSUBS 0.06929f $ **FLOATING
C9762 a_65865_57675# VSUBS 0.1022f $ **FLOATING
C9763 a_63391_57320# VSUBS 0.03882f $ **FLOATING
C9764 a_63045_57628# VSUBS 0.03327f $ **FLOATING
C9765 a_62793_57675# VSUBS 0.06954f $ **FLOATING
C9766 a_62357_57455# VSUBS 0.03316f $ **FLOATING
C9767 a_62222_57356# VSUBS 0.03547f $ **FLOATING
C9768 a_62017_57307# VSUBS 0.06935f $ **FLOATING
C9769 a_61833_57675# VSUBS 0.10195f $ **FLOATING
C9770 sar10b_0.net6 VSUBS 0.23018f $ **FLOATING
C9771 a_60747_57571# VSUBS 0.03328f $ **FLOATING
C9772 a_65966_58354# VSUBS 0.03547f $ **FLOATING
C9773 sar10b_0.net36 VSUBS 0.4561f $ **FLOATING
C9774 a_67135_58306# VSUBS 0.03739f $ **FLOATING
C9775 a_66537_57971# VSUBS 0.06971f $ **FLOATING
C9776 a_66789_58100# VSUBS 0.03351f $ **FLOATING
C9777 a_66101_58256# VSUBS 0.03316f $ **FLOATING
C9778 a_65761_58263# VSUBS 0.06932f $ **FLOATING
C9779 a_65577_57971# VSUBS 0.10356f $ **FLOATING
C9780 a_61358_58354# VSUBS 0.03547f $ **FLOATING
C9781 a_62527_58306# VSUBS 0.03838f $ **FLOATING
C9782 a_61929_57971# VSUBS 0.06997f $ **FLOATING
C9783 a_62181_58100# VSUBS 0.03344f $ **FLOATING
C9784 a_61493_58256# VSUBS 0.03316f $ **FLOATING
C9785 a_61153_58263# VSUBS 0.06966f $ **FLOATING
C9786 a_60969_57971# VSUBS 0.11151f $ **FLOATING
C9787 sar10b_0.net19 VSUBS 0.056f $ **FLOATING
C9788 a_68767_58652# VSUBS 0.03895f $ **FLOATING
C9789 a_68421_58960# VSUBS 0.03385f $ **FLOATING
C9790 a_68169_59007# VSUBS 0.07191f $ **FLOATING
C9791 a_67733_58787# VSUBS 0.03316f $ **FLOATING
C9792 a_67598_58688# VSUBS 0.03553f $ **FLOATING
C9793 a_67393_58639# VSUBS 0.07008f $ **FLOATING
C9794 a_67209_59007# VSUBS 0.10732f $ **FLOATING
C9795 sar10b_0.net32 VSUBS 0.07347f $ **FLOATING
C9796 a_63967_58652# VSUBS 0.03812f $ **FLOATING
C9797 a_63621_58960# VSUBS 0.03364f $ **FLOATING
C9798 a_63369_59007# VSUBS 0.07029f $ **FLOATING
C9799 a_62933_58787# VSUBS 0.03393f $ **FLOATING
C9800 a_62798_58688# VSUBS 0.03682f $ **FLOATING
C9801 a_62593_58639# VSUBS 0.06977f $ **FLOATING
C9802 a_62409_59007# VSUBS 0.10471f $ **FLOATING
C9803 sar10b_0.net7 VSUBS 0.45796f $ **FLOATING
C9804 a_60747_58903# VSUBS 0.03328f $ **FLOATING
C9805 a_68946_59303# VSUBS 0.03607f $ **FLOATING
C9806 a_64910_59686# VSUBS 0.03569f $ **FLOATING
C9807 sar10b_0.net34 VSUBS 0.06415f $ **FLOATING
C9808 a_66079_59638# VSUBS 0.04048f $ **FLOATING
C9809 a_65481_59303# VSUBS 0.07185f $ **FLOATING
C9810 a_65733_59432# VSUBS 0.03385f $ **FLOATING
C9811 a_65045_59588# VSUBS 0.03393f $ **FLOATING
C9812 a_64705_59595# VSUBS 0.07156f $ **FLOATING
C9813 a_51603_58977# VSUBS 0.02403f $ **FLOATING
C9814 a_64521_59303# VSUBS 0.1087f $ **FLOATING
C9815 sar10b_0.net21 VSUBS 0.06493f $ **FLOATING
C9816 a_68479_59984# VSUBS 0.03662f $ **FLOATING
C9817 a_68133_60292# VSUBS 0.03317f $ **FLOATING
C9818 a_67881_60339# VSUBS 0.0693f $ **FLOATING
C9819 a_67445_60119# VSUBS 0.03316f $ **FLOATING
C9820 a_67310_60020# VSUBS 0.03547f $ **FLOATING
C9821 a_67105_59971# VSUBS 0.06885f $ **FLOATING
C9822 a_66921_60339# VSUBS 0.10312f $ **FLOATING
C9823 sar10b_0.net33 VSUBS 0.06641f $ **FLOATING
C9824 a_65119_59984# VSUBS 0.03738f $ **FLOATING
C9825 a_64773_60292# VSUBS 0.03385f $ **FLOATING
C9826 a_64521_60339# VSUBS 0.06988f $ **FLOATING
C9827 a_64085_60119# VSUBS 0.03345f $ **FLOATING
C9828 a_63950_60020# VSUBS 0.03682f $ **FLOATING
C9829 a_63745_59971# VSUBS 0.07084f $ **FLOATING
C9830 tdc_0.RDY VSUBS 3.15025f $ **FLOATING
C9831 a_55121_59650# VSUBS 0.04037f $ **FLOATING
C9832 a_53564_59480# VSUBS 0.02133f $ **FLOATING
C9833 a_52417_59293# VSUBS 0.03521f $ **FLOATING
C9834 tdc_0.delay_gate_ori_1.sky130_fd_sc_hs__and2_1_0.A VSUBS 0.10957f $ **FLOATING
C9835 a_51861_59345# VSUBS 0.07865f $ **FLOATING
C9836 a_51345_58977# VSUBS 0.36323f $ **FLOATING
C9837 a_n9133_57045# VSUBS 0.6686f $ **FLOATING
C9838 th_dif_sw_0.th_sw_0.th_sw_main_0.VGS VSUBS 1.31272f $ **FLOATING
C9839 tdc_0.OUTN VSUBS 1.81995f $ **FLOATING
C9840 a_63561_60339# VSUBS 0.10571f $ **FLOATING
C9841 sar10b_0.net1 VSUBS 0.54298f $ **FLOATING
C9842 a_60747_60235# VSUBS 0.03922f $ **FLOATING
C9843 a_61677_60846# VSUBS 0.03682f $ **FLOATING
C9844 a_61609_60938# VSUBS 0.03393f $ **FLOATING
C9845 a_61400_60956# VSUBS 0.07163f $ **FLOATING
C9846 a_61086_60642# VSUBS 0.03385f $ **FLOATING
C9847 a_60945_60609# VSUBS 0.07029f $ **FLOATING
C9848 a_53564_60302# VSUBS 0.02133f $ **FLOATING
C9849 a_61395_60616# VSUBS 0.10483f $ **FLOATING
C9850 a_60747_60609# VSUBS 0.03683f $ **FLOATING
C9851 sar10b_0.net22 VSUBS 0.17039f $ **FLOATING
C9852 tdc_0.phase_detector_0.pd_out_0.B VSUBS 0.35505f $ **FLOATING
C9853 tdc_0.phase_detector_0.INP VSUBS 0.11803f $ **FLOATING
C9854 a_51861_60437# VSUBS 0.07865f $ **FLOATING
C9855 a_52417_60961# VSUBS 0.03527f $ **FLOATING
C9856 a_68946_61735# VSUBS 0.03333f $ **FLOATING
C9857 a_68479_61316# VSUBS 0.03662f $ **FLOATING
C9858 a_68133_61624# VSUBS 0.03316f $ **FLOATING
C9859 a_67881_61671# VSUBS 0.06926f $ **FLOATING
C9860 a_67445_61451# VSUBS 0.03316f $ **FLOATING
C9861 a_67310_61352# VSUBS 0.03547f $ **FLOATING
C9862 a_67105_61303# VSUBS 0.06915f $ **FLOATING
C9863 a_66921_61671# VSUBS 0.10289f $ **FLOATING
C9864 tdc_0.phase_detector_0.pd_out_0.A VSUBS 0.30959f $ **FLOATING
C9865 tdc_0.phase_detector_0.INN VSUBS 0.10813f $ **FLOATING
C9866 a_63871_61316# VSUBS 0.03647f $ **FLOATING
C9867 a_63525_61624# VSUBS 0.03385f $ **FLOATING
C9868 a_63273_61671# VSUBS 0.06874f $ **FLOATING
C9869 a_62837_61451# VSUBS 0.03323f $ **FLOATING
C9870 a_62702_61352# VSUBS 0.03574f $ **FLOATING
C9871 a_62497_61303# VSUBS 0.06906f $ **FLOATING
C9872 tdc_0.delay_gate_ori_0.sky130_fd_sc_hs__and2_1_0.A VSUBS 0.10957f $ **FLOATING
C9873 a_51603_61205# VSUBS 0.02403f $ **FLOATING
C9874 a_51345_60437# VSUBS 0.36323f $ **FLOATING
C9875 th_dif_sw_0.VCN VSUBS 23.1467f $ **FLOATING
C9876 a_62313_61671# VSUBS 0.10889f $ **FLOATING
C9877 sar10b_0.net8 VSUBS 0.24783f $ **FLOATING
C9878 a_60747_61567# VSUBS 0.03328f $ **FLOATING
C9879 a_61677_62178# VSUBS 0.03547f $ **FLOATING
C9880 a_61609_62270# VSUBS 0.03316f $ **FLOATING
C9881 a_61400_62288# VSUBS 0.06885f $ **FLOATING
C9882 a_61086_61974# VSUBS 0.03316f $ **FLOATING
C9883 a_60945_61941# VSUBS 0.06867f $ **FLOATING
C9884 a_61395_61948# VSUBS 0.10173f $ **FLOATING
C9885 a_60747_61941# VSUBS 0.03633f $ **FLOATING
C9886 sar10b_0.net24 VSUBS 0.11092f $ **FLOATING
C9887 a_68767_62648# VSUBS 0.03763f $ **FLOATING
C9888 a_68421_62956# VSUBS 0.03316f $ **FLOATING
C9889 a_68169_63003# VSUBS 0.06955f $ **FLOATING
C9890 a_67733_62783# VSUBS 0.03316f $ **FLOATING
C9891 a_67598_62684# VSUBS 0.03547f $ **FLOATING
C9892 a_67393_62635# VSUBS 0.06903f $ **FLOATING
C9893 a_67209_63003# VSUBS 0.10262f $ **FLOATING
C9894 a_64543_62648# VSUBS 0.03843f $ **FLOATING
C9895 a_64197_62956# VSUBS 0.03385f $ **FLOATING
C9896 a_63945_63003# VSUBS 0.07098f $ **FLOATING
C9897 a_63509_62783# VSUBS 0.03393f $ **FLOATING
C9898 a_63374_62684# VSUBS 0.03615f $ **FLOATING
C9899 a_63169_62635# VSUBS 0.07052f $ **FLOATING
C9900 a_62985_63003# VSUBS 0.10487f $ **FLOATING
C9901 sar10b_0.net9 VSUBS 0.20916f $ **FLOATING
C9902 a_60747_62899# VSUBS 0.0426f $ **FLOATING
C9903 a_68946_63299# VSUBS 0.03602f $ **FLOATING
C9904 a_64238_63682# VSUBS 0.03547f $ **FLOATING
C9905 a_65407_63634# VSUBS 0.04087f $ **FLOATING
C9906 a_64809_63299# VSUBS 0.07202f $ **FLOATING
C9907 a_65061_63428# VSUBS 0.03316f $ **FLOATING
C9908 a_64373_63584# VSUBS 0.0332f $ **FLOATING
C9909 a_64033_63591# VSUBS 0.07064f $ **FLOATING
C9910 a_63849_63299# VSUBS 0.1058f $ **FLOATING
C9911 sar10b_0.net10 VSUBS 0.23927f $ **FLOATING
C9912 a_61677_63510# VSUBS 0.03547f $ **FLOATING
C9913 a_61609_63602# VSUBS 0.03316f $ **FLOATING
C9914 a_61400_63620# VSUBS 0.06885f $ **FLOATING
C9915 a_61086_63306# VSUBS 0.03316f $ **FLOATING
C9916 a_60945_63273# VSUBS 0.06867f $ **FLOATING
C9917 a_61395_63280# VSUBS 0.10173f $ **FLOATING
C9918 a_60747_63273# VSUBS 0.03633f $ **FLOATING
C9919 sar10b_0.net23 VSUBS 0.10684f $ **FLOATING
C9920 a_68767_63980# VSUBS 0.03633f $ **FLOATING
C9921 a_68421_64288# VSUBS 0.03316f $ **FLOATING
C9922 a_68169_64335# VSUBS 0.06867f $ **FLOATING
C9923 a_67733_64115# VSUBS 0.03316f $ **FLOATING
C9924 a_67598_64016# VSUBS 0.03547f $ **FLOATING
C9925 a_67393_63967# VSUBS 0.06885f $ **FLOATING
C9926 a_67209_64335# VSUBS 0.10173f $ **FLOATING
C9927 a_60747_64231# VSUBS 0.0426f $ **FLOATING
C9928 th_dif_sw_0.VCP VSUBS 23.1328f $ **FLOATING
C9929 a_64814_65014# VSUBS 0.03576f $ **FLOATING
C9930 a_65983_64966# VSUBS 0.04092f $ **FLOATING
C9931 a_65385_64631# VSUBS 0.07234f $ **FLOATING
C9932 a_65637_64760# VSUBS 0.0336f $ **FLOATING
C9933 a_64949_64916# VSUBS 0.03316f $ **FLOATING
C9934 a_64609_64923# VSUBS 0.06885f $ **FLOATING
C9935 a_64425_64631# VSUBS 0.10434f $ **FLOATING
C9936 sar10b_0.net11 VSUBS 0.25793f $ **FLOATING
C9937 a_61677_64842# VSUBS 0.03547f $ **FLOATING
C9938 a_61609_64934# VSUBS 0.03316f $ **FLOATING
C9939 a_61400_64952# VSUBS 0.06885f $ **FLOATING
C9940 a_61086_64638# VSUBS 0.03316f $ **FLOATING
C9941 a_60945_64605# VSUBS 0.06867f $ **FLOATING
C9942 a_61395_64612# VSUBS 0.10173f $ **FLOATING
C9943 a_60747_64605# VSUBS 0.03633f $ **FLOATING
C9944 sar10b_0.net25 VSUBS 0.14852f $ **FLOATING
C9945 a_68767_65312# VSUBS 0.03633f $ **FLOATING
C9946 a_68421_65620# VSUBS 0.03316f $ **FLOATING
C9947 a_68169_65667# VSUBS 0.06867f $ **FLOATING
C9948 a_67733_65447# VSUBS 0.03316f $ **FLOATING
C9949 a_67598_65348# VSUBS 0.03547f $ **FLOATING
C9950 a_67393_65299# VSUBS 0.06885f $ **FLOATING
C9951 a_67209_65667# VSUBS 0.10173f $ **FLOATING
C9952 a_60747_65563# VSUBS 0.0426f $ **FLOATING
C9953 th_dif_sw_0.th_sw_1.th_sw_main_0.VGS VSUBS 1.31272f $ **FLOATING
C9954 a_n8277_65767# VSUBS 0.44237f $ **FLOATING
C9955 a_68946_65963# VSUBS 0.03338f $ **FLOATING
C9956 a_65198_66346# VSUBS 0.03591f $ **FLOATING
C9957 a_66367_66298# VSUBS 0.03643f $ **FLOATING
C9958 a_65769_65963# VSUBS 0.07254f $ **FLOATING
C9959 a_66021_66092# VSUBS 0.03385f $ **FLOATING
C9960 a_65333_66248# VSUBS 0.03316f $ **FLOATING
C9961 a_64993_66255# VSUBS 0.06995f $ **FLOATING
C9962 a_64809_65963# VSUBS 0.10976f $ **FLOATING
C9963 sar10b_0.net12 VSUBS 0.32746f $ **FLOATING
C9964 a_61677_66174# VSUBS 0.03547f $ **FLOATING
C9965 a_61609_66266# VSUBS 0.03316f $ **FLOATING
C9966 a_61400_66284# VSUBS 0.06885f $ **FLOATING
C9967 a_61086_65970# VSUBS 0.03316f $ **FLOATING
C9968 a_60945_65937# VSUBS 0.06975f $ **FLOATING
C9969 a_n8277_66083# VSUBS 4.76062f $ **FLOATING
C9970 a_n9133_63315# VSUBS 0.6686f $ **FLOATING
C9971 th_dif_sw_0.th_sw_1.CKB VSUBS 2.53243f $ **FLOATING
C9972 a_61395_65944# VSUBS 0.10289f $ **FLOATING
C9973 a_60747_65937# VSUBS 0.03707f $ **FLOATING
C9974 sar10b_0.net26 VSUBS 0.09967f $ **FLOATING
C9975 a_68767_66644# VSUBS 0.03633f $ **FLOATING
C9976 a_68421_66952# VSUBS 0.03316f $ **FLOATING
C9977 a_68169_66999# VSUBS 0.06867f $ **FLOATING
C9978 a_67733_66779# VSUBS 0.03316f $ **FLOATING
C9979 a_67598_66680# VSUBS 0.03547f $ **FLOATING
C9980 a_67393_66631# VSUBS 0.06885f $ **FLOATING
C9981 th_dif_sw_0.th_sw_1.CK VSUBS 0.84578f $ **FLOATING
C9982 a_67209_66999# VSUBS 0.10173f $ **FLOATING
C9983 a_n4470_65264# VSUBS 0.64281f $ **FLOATING
C9984 a_63663_67678# VSUBS 0.03464f $ **FLOATING
C9985 a_64888_67630# VSUBS 0.06856f $ **FLOATING
C9986 a_64238_67295# VSUBS 0.07155f $ **FLOATING
C9987 a_64492_67433# VSUBS 0.03442f $ **FLOATING
C9988 a_63804_67580# VSUBS 0.03442f $ **FLOATING
C9989 a_63457_67583# VSUBS 0.07201f $ **FLOATING
C9990 a_63273_67295# VSUBS 0.11573f $ **FLOATING
C9991 a_61358_67678# VSUBS 0.03547f $ **FLOATING
C9992 a_62527_67630# VSUBS 0.03912f $ **FLOATING
C9993 a_61929_67295# VSUBS 0.06952f $ **FLOATING
C9994 a_62181_67424# VSUBS 0.03385f $ **FLOATING
C9995 a_61493_67580# VSUBS 0.03316f $ **FLOATING
C9996 a_61153_67587# VSUBS 0.06982f $ **FLOATING
C9997 a_60969_67295# VSUBS 0.11222f $ **FLOATING
C9998 sar10b_0.net4 VSUBS 0.59847f $ **FLOATING
C9999 a_68767_67976# VSUBS 0.03758f $ **FLOATING
C10000 a_68421_68284# VSUBS 0.03385f $ **FLOATING
C10001 a_68169_68331# VSUBS 0.07103f $ **FLOATING
C10002 a_67733_68111# VSUBS 0.03327f $ **FLOATING
C10003 a_67598_68012# VSUBS 0.03597f $ **FLOATING
C10004 a_67393_67963# VSUBS 0.07034f $ **FLOATING
C10005 a_67209_68331# VSUBS 0.10301f $ **FLOATING
C10006 sar10b_0.net3 VSUBS 1.45805f $ **FLOATING
C10007 a_60747_68227# VSUBS 0.0431f $ **FLOATING
C10008 a_68946_68627# VSUBS 0.03338f $ **FLOATING
C10009 sar10b_0.net27 VSUBS 0.08896f $ **FLOATING
C10010 a_65390_69010# VSUBS 0.03682f $ **FLOATING
C10011 a_67055_68689# VSUBS 0.03365f $ **FLOATING
C10012 sar10b_0.cyclic_flag_0.FINAL VSUBS 0.5844f $ **FLOATING
C10013 a_66559_68962# VSUBS 0.03837f $ **FLOATING
C10014 a_65961_68627# VSUBS 0.0685f $ **FLOATING
C10015 a_66213_68756# VSUBS 0.03385f $ **FLOATING
C10016 a_65525_68912# VSUBS 0.03393f $ **FLOATING
C10017 a_65185_68919# VSUBS 0.07163f $ **FLOATING
C10018 a_65001_68627# VSUBS 0.11207f $ **FLOATING
C10019 sar10b_0.net13 VSUBS 0.29111f $ **FLOATING
C10020 a_67890_69727# VSUBS 0.03424f $ **FLOATING
C10021 sar10b_0._06_ VSUBS 0.10382f $ **FLOATING
C10022 a_67423_69308# VSUBS 0.03811f $ **FLOATING
C10023 a_67077_69616# VSUBS 0.03385f $ **FLOATING
C10024 a_66825_69663# VSUBS 0.07141f $ **FLOATING
C10025 a_66389_69443# VSUBS 0.03393f $ **FLOATING
C10026 a_66254_69344# VSUBS 0.03682f $ **FLOATING
C10027 a_66049_69295# VSUBS 0.07131f $ **FLOATING
C10028 a_65865_69663# VSUBS 0.10839f $ **FLOATING
C10029 sar10b_0.net14 VSUBS 0.32658f $ **FLOATING
C10030 a_60747_69559# VSUBS 0.04298f $ **FLOATING
C10031 a_68946_71059# VSUBS 0.04272f $ **FLOATING
C10032 sar10b_0.net47 VSUBS 0.13679f $ **FLOATING
C10033 sar10b_0.net2 VSUBS 0.58012f $ **FLOATING
C10034 sar10b_0.net38 VSUBS 0.28999f $ **FLOATING
C10035 a_61131_70891# VSUBS 0.04379f $ **FLOATING
C10036 a_60690_70625# VSUBS 0.07107f $ **FLOATING
C10037 tdc_0.OUTP VSUBS 4.28464f $ **FLOATING
C10038 sar10b_0.net46 VSUBS 0.11908f $ **FLOATING
C10039 a_69003_71265# VSUBS 0.03406f $ **FLOATING
C10040 a_68562_71291# VSUBS 0.03496f $ **FLOATING
C10041 sar10b_0.net15 VSUBS 0.13372f $ **FLOATING
C10042 sar10b_0.net45 VSUBS 0.1018f $ **FLOATING
C10043 a_68235_71265# VSUBS 0.03496f $ **FLOATING
C10044 sar10b_0.net44 VSUBS 0.11796f $ **FLOATING
C10045 a_66795_71265# VSUBS 0.03465f $ **FLOATING
C10046 sar10b_0.net43 VSUBS 0.11815f $ **FLOATING
C10047 a_65643_71265# VSUBS 0.03456f $ **FLOATING
C10048 sar10b_0.net42 VSUBS 0.32039f $ **FLOATING
C10049 a_64491_71265# VSUBS 0.03496f $ **FLOATING
C10050 sar10b_0.net41 VSUBS 0.13925f $ **FLOATING
C10051 a_63339_71265# VSUBS 0.03496f $ **FLOATING
C10052 th_dif_sw_0.CK VSUBS 9.30918f $ **FLOATING
C10053 sar10b_0.net40 VSUBS 0.22391f $ **FLOATING
C10054 a_62187_71265# VSUBS 0.03496f $ **FLOATING
C10055 sar10b_0.net16 VSUBS 3.84761f $ **FLOATING
C10056 a_61419_71265# VSUBS 0.03496f $ **FLOATING
C10057 sar10b_0.net39 VSUBS 0.14593f $ **FLOATING
C10058 a_61035_71265# VSUBS 0.03508f $ **FLOATING
C10059 sar10b_0.CF[0] VSUBS 5.33124f $ **FLOATING
C10060 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x3.Y VSUBS 0.035f $ **FLOATING
C10061 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06692f $ **FLOATING
C10062 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x4.A VSUBS 0.05619f $ **FLOATING
C10063 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03496f $ **FLOATING
C10064 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x6.A VSUBS 0.034f $ **FLOATING
C10065 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x1.A VSUBS 0.22255f $ **FLOATING
C10066 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x8.A VSUBS 0.21343f $ **FLOATING
C10067 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27932f $ **FLOATING
C10068 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.x10.A VSUBS 0.27476f $ **FLOATING
C10069 a_44345_110521# VSUBS 0.22209f $ **FLOATING
C10070 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLK0 VSUBS 1.32788f $ **FLOATING
C10071 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.nooverlap_clk_0.CLKB0 VSUBS 1.76172f $ **FLOATING
C10072 a_43467_106170# VSUBS 0.76225f $ **FLOATING
C10073 sar10b_0.SWP[0] VSUBS 22.2183f $ **FLOATING
C10074 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[0] VSUBS 6.81604f $ **FLOATING
C10075 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWP VSUBS 5.81794f $ **FLOATING
C10076 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_1_0.tg_sw_1_2.SWN VSUBS 4.42867f $ **FLOATING
C10077 sar10b_0.CF[1] VSUBS 3.42286f $ **FLOATING
C10078 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x3.Y VSUBS 0.035f $ **FLOATING
C10079 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06826f $ **FLOATING
C10080 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x4.A VSUBS 0.05619f $ **FLOATING
C10081 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03399f $ **FLOATING
C10082 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x6.A VSUBS 0.034f $ **FLOATING
C10083 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x1.A VSUBS 0.25929f $ **FLOATING
C10084 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x8.A VSUBS 0.21745f $ **FLOATING
C10085 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27474f $ **FLOATING
C10086 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.x10.A VSUBS 0.27476f $ **FLOATING
C10087 a_39543_110941# VSUBS 0.20157f $ **FLOATING
C10088 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLK0 VSUBS 1.20219f $ **FLOATING
C10089 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.nooverlap_clk_0.CLKB0 VSUBS 1.61928f $ **FLOATING
C10090 a_38665_107026# VSUBS 0.68771f $ **FLOATING
C10091 sar10b_0.SWP[1] VSUBS 18.9244f $ **FLOATING
C10092 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[1] VSUBS 3.66021f $ **FLOATING
C10093 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWP VSUBS 5.31078f $ **FLOATING
C10094 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_2_0.tg_sw_2_2.SWN VSUBS 4.03497f $ **FLOATING
C10095 sar10b_0.CF[2] VSUBS 2.70866f $ **FLOATING
C10096 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x3.Y VSUBS 0.035f $ **FLOATING
C10097 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06825f $ **FLOATING
C10098 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x4.A VSUBS 0.05619f $ **FLOATING
C10099 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03399f $ **FLOATING
C10100 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x6.A VSUBS 0.034f $ **FLOATING
C10101 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x1.A VSUBS 0.25929f $ **FLOATING
C10102 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x8.A VSUBS 0.21745f $ **FLOATING
C10103 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27473f $ **FLOATING
C10104 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.x10.A VSUBS 0.27476f $ **FLOATING
C10105 a_34741_111361# VSUBS 0.18104f $ **FLOATING
C10106 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLK0 VSUBS 1.07669f $ **FLOATING
C10107 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.nooverlap_clk_0.CLKB0 VSUBS 1.47858f $ **FLOATING
C10108 a_33863_107882# VSUBS 0.61316f $ **FLOATING
C10109 sar10b_0.SWP[2] VSUBS 19.8581f $ **FLOATING
C10110 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[2] VSUBS 2.98506f $ **FLOATING
C10111 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWP VSUBS 4.7468f $ **FLOATING
C10112 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_3_0.tg_sw_3_3.SWN VSUBS 3.641f $ **FLOATING
C10113 sar10b_0.CF[3] VSUBS 3.59461f $ **FLOATING
C10114 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x3.Y VSUBS 0.03532f $ **FLOATING
C10115 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06825f $ **FLOATING
C10116 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x4.A VSUBS 0.05619f $ **FLOATING
C10117 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03399f $ **FLOATING
C10118 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x6.A VSUBS 0.034f $ **FLOATING
C10119 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x1.A VSUBS 0.25929f $ **FLOATING
C10120 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x8.A VSUBS 0.21745f $ **FLOATING
C10121 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27473f $ **FLOATING
C10122 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.x10.A VSUBS 0.27476f $ **FLOATING
C10123 a_29939_111781# VSUBS 0.16052f $ **FLOATING
C10124 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLK0 VSUBS 0.95119f $ **FLOATING
C10125 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.nooverlap_clk_0.CLKB0 VSUBS 1.33767f $ **FLOATING
C10126 a_29061_108738# VSUBS 0.53862f $ **FLOATING
C10127 sar10b_0.SWP[3] VSUBS 20.6716f $ **FLOATING
C10128 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[3] VSUBS 2.52477f $ **FLOATING
C10129 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWP VSUBS 4.16372f $ **FLOATING
C10130 sar10b_0.CF[4] VSUBS 4.05359f $ **FLOATING
C10131 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_4_0.tg_sw_4_4.SWN VSUBS 3.22955f $ **FLOATING
C10132 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x3.Y VSUBS 0.03532f $ **FLOATING
C10133 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06825f $ **FLOATING
C10134 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x4.A VSUBS 0.05733f $ **FLOATING
C10135 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03399f $ **FLOATING
C10136 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x6.A VSUBS 0.034f $ **FLOATING
C10137 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x1.A VSUBS 0.25984f $ **FLOATING
C10138 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x8.A VSUBS 0.21745f $ **FLOATING
C10139 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27473f $ **FLOATING
C10140 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.x10.A VSUBS 0.27476f $ **FLOATING
C10141 a_25137_112201# VSUBS 0.13999f $ **FLOATING
C10142 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLK0 VSUBS 0.8257f $ **FLOATING
C10143 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.nooverlap_clk_0.CLKB0 VSUBS 1.19685f $ **FLOATING
C10144 a_24259_109594# VSUBS 0.46408f $ **FLOATING
C10145 sar10b_0.SWP[4] VSUBS 21.4186f $ **FLOATING
C10146 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[4] VSUBS 2.90183f $ **FLOATING
C10147 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWP VSUBS 3.59961f $ **FLOATING
C10148 sar10b_0.CF[5] VSUBS 3.5484f $ **FLOATING
C10149 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x3.Y VSUBS 0.03532f $ **FLOATING
C10150 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06923f $ **FLOATING
C10151 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x4.A VSUBS 0.05733f $ **FLOATING
C10152 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_5_0.tg_sw_5_5.SWN VSUBS 2.83745f $ **FLOATING
C10153 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03399f $ **FLOATING
C10154 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x6.A VSUBS 0.03496f $ **FLOATING
C10155 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x1.A VSUBS 0.25984f $ **FLOATING
C10156 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x8.A VSUBS 0.21778f $ **FLOATING
C10157 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27473f $ **FLOATING
C10158 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.x10.A VSUBS 0.27476f $ **FLOATING
C10159 a_20335_112621# VSUBS 0.11946f $ **FLOATING
C10160 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLK0 VSUBS 0.7002f $ **FLOATING
C10161 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.nooverlap_clk_0.CLKB0 VSUBS 1.05653f $ **FLOATING
C10162 a_19457_110450# VSUBS 0.38954f $ **FLOATING
C10163 sar10b_0.SWP[5] VSUBS 22.1328f $ **FLOATING
C10164 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[5] VSUBS 3.19494f $ **FLOATING
C10165 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWP VSUBS 3.03512f $ **FLOATING
C10166 sar10b_0.CF[6] VSUBS 4.19596f $ **FLOATING
C10167 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x3.Y VSUBS 0.03532f $ **FLOATING
C10168 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06883f $ **FLOATING
C10169 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x4.A VSUBS 0.05733f $ **FLOATING
C10170 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03445f $ **FLOATING
C10171 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x6.A VSUBS 0.03496f $ **FLOATING
C10172 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_6_0.tg_sw_6_6.SWN VSUBS 2.44487f $ **FLOATING
C10173 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x1.A VSUBS 0.25984f $ **FLOATING
C10174 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x8.A VSUBS 0.21915f $ **FLOATING
C10175 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27473f $ **FLOATING
C10176 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.x10.A VSUBS 0.27476f $ **FLOATING
C10177 a_15533_113041# VSUBS 0.09894f $ **FLOATING
C10178 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLK0 VSUBS 0.5747f $ **FLOATING
C10179 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.nooverlap_clk_0.CLKB0 VSUBS 0.91609f $ **FLOATING
C10180 a_14655_111306# VSUBS 0.315f $ **FLOATING
C10181 sar10b_0.SWP[6] VSUBS 22.8133f $ **FLOATING
C10182 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[6] VSUBS 3.14107f $ **FLOATING
C10183 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWP VSUBS 2.47031f $ **FLOATING
C10184 sar10b_0.CF[7] VSUBS 4.24451f $ **FLOATING
C10185 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x3.Y VSUBS 0.03563f $ **FLOATING
C10186 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06891f $ **FLOATING
C10187 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x4.A VSUBS 0.05733f $ **FLOATING
C10188 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03402f $ **FLOATING
C10189 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x6.A VSUBS 0.03496f $ **FLOATING
C10190 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x1.A VSUBS 0.26095f $ **FLOATING
C10191 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x8.A VSUBS 0.21907f $ **FLOATING
C10192 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_7_0.tg_sw_7_7.SWN VSUBS 2.05286f $ **FLOATING
C10193 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27473f $ **FLOATING
C10194 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.x10.A VSUBS 0.27589f $ **FLOATING
C10195 a_10731_113461# VSUBS 0.07841f $ **FLOATING
C10196 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLK0 VSUBS 0.44921f $ **FLOATING
C10197 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.nooverlap_clk_0.CLKB0 VSUBS 0.77702f $ **FLOATING
C10198 a_9853_112162# VSUBS 0.24046f $ **FLOATING
C10199 sar10b_0.SWP[7] VSUBS 23.5031f $ **FLOATING
C10200 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[7] VSUBS 1.97347f $ **FLOATING
C10201 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWP VSUBS 1.90627f $ **FLOATING
C10202 sar10b_0.CF[8] VSUBS 4.63235f $ **FLOATING
C10203 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x3.Y VSUBS 0.03563f $ **FLOATING
C10204 sar10b_0.CF[9] VSUBS 28.9156f $ **FLOATING
C10205 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06899f $ **FLOATING
C10206 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x4.A VSUBS 0.05733f $ **FLOATING
C10207 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.0341f $ **FLOATING
C10208 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x6.A VSUBS 0.03496f $ **FLOATING
C10209 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x1.A VSUBS 0.2605f $ **FLOATING
C10210 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x8.A VSUBS 0.2195f $ **FLOATING
C10211 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_8_0.tg_sw_8_8.SWN VSUBS 1.66072f $ **FLOATING
C10212 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27588f $ **FLOATING
C10213 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.x10.A VSUBS 0.27719f $ **FLOATING
C10214 a_5929_113881# VSUBS 0.05789f $ **FLOATING
C10215 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLK0 VSUBS 0.32373f $ **FLOATING
C10216 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.nooverlap_clk_0.CLKB0 VSUBS 0.63619f $ **FLOATING
C10217 a_5051_113018# VSUBS 0.16592f $ **FLOATING
C10218 sar10b_0.SWP[8] VSUBS 24.3683f $ **FLOATING
C10219 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[8] VSUBS 1.84658f $ **FLOATING
C10220 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x3.Y VSUBS 0.03563f $ **FLOATING
C10221 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWP VSUBS 1.36627f $ **FLOATING
C10222 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__nand2_1_0.Y VSUBS 0.06854f $ **FLOATING
C10223 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x4.A VSUBS 0.05733f $ **FLOATING
C10224 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_1_1.A VSUBS 0.03402f $ **FLOATING
C10225 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x6.A VSUBS 0.03496f $ **FLOATING
C10226 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x1.A VSUBS 0.21523f $ **FLOATING
C10227 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x8.A VSUBS 0.21886f $ **FLOATING
C10228 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_9_0.tg_sw_9_9.SWN VSUBS 1.26891f $ **FLOATING
C10229 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.sky130_fd_sc_hs__inv_8_0.A VSUBS 0.27607f $ **FLOATING
C10230 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.x10.A VSUBS 0.27893f $ **FLOATING
C10231 a_1127_114301# VSUBS 0.03736f $ **FLOATING
C10232 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLK0 VSUBS 0.19828f $ **FLOATING
C10233 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.nooverlap_clk_0.CLKB0 VSUBS 0.4974f $ **FLOATING
C10234 a_249_113874# VSUBS 0.09138f $ **FLOATING
C10235 sar10b_0.SWP[9] VSUBS 30.9434f $ **FLOATING
C10236 cdac_0.single_10b_cdac_1.x10b_cap_array_0.SW[9] VSUBS 1.7415f $ **FLOATING
C10237 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWP VSUBS 0.98472f $ **FLOATING
C10238 cdac_0.single_10b_cdac_1.cdac_sw_10b_0.cdac_sw_10_0.tg_sw_10_10.SWN VSUBS 0.88042f $ **FLOATING
C10239 w_n9655_56533# VSUBS 5.30723f $ **FLOATING
C10240 w_n9655_63119# VSUBS 5.32398f $ **FLOATING
.ends
