magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect 142 1527 148 1561
rect 182 1527 220 1561
rect 254 1527 292 1561
rect 326 1527 364 1561
rect 398 1527 436 1561
rect 470 1527 508 1561
rect 542 1527 580 1561
rect 614 1527 652 1561
rect 686 1527 724 1561
rect 758 1527 796 1561
rect 830 1527 868 1561
rect 902 1527 940 1561
rect 974 1527 1012 1561
rect 1046 1527 1084 1561
rect 1118 1527 1156 1561
rect 1190 1527 1228 1561
rect 1262 1527 1300 1561
rect 1334 1527 1372 1561
rect 1406 1527 1444 1561
rect 1478 1527 1516 1561
rect 1550 1527 1588 1561
rect 1622 1527 1660 1561
rect 1694 1527 1732 1561
rect 1766 1527 1804 1561
rect 1838 1527 1876 1561
rect 1910 1527 1948 1561
rect 1982 1527 2020 1561
rect 2054 1527 2092 1561
rect 2126 1527 2164 1561
rect 2198 1527 2236 1561
rect 2270 1527 2308 1561
rect 2342 1527 2380 1561
rect 2414 1527 2452 1561
rect 2486 1527 2524 1561
rect 2558 1527 2596 1561
rect 2630 1527 2668 1561
rect 2702 1527 2740 1561
rect 2774 1527 2812 1561
rect 2846 1527 2884 1561
rect 2918 1527 2956 1561
rect 2990 1527 3028 1561
rect 3062 1527 3100 1561
rect 3134 1527 3172 1561
rect 3206 1527 3244 1561
rect 3278 1527 3316 1561
rect 3350 1527 3388 1561
rect 3422 1527 3460 1561
rect 3494 1527 3532 1561
rect 3566 1527 3604 1561
rect 3638 1527 3676 1561
rect 3710 1527 3748 1561
rect 3782 1527 3820 1561
rect 3854 1527 3892 1561
rect 3926 1527 3964 1561
rect 3998 1527 4036 1561
rect 4070 1527 4108 1561
rect 4142 1527 4180 1561
rect 4214 1527 4252 1561
rect 4286 1527 4324 1561
rect 4358 1527 4396 1561
rect 4430 1527 4468 1561
rect 4502 1527 4540 1561
rect 4574 1527 4612 1561
rect 4646 1527 4684 1561
rect 4718 1527 4756 1561
rect 4790 1527 4828 1561
rect 4862 1527 4900 1561
rect 4934 1527 4972 1561
rect 5006 1527 5044 1561
rect 5078 1527 5116 1561
rect 5150 1527 5188 1561
rect 5222 1527 5260 1561
rect 5294 1527 5332 1561
rect 5366 1527 5404 1561
rect 5438 1527 5476 1561
rect 5510 1527 5516 1561
rect 142 -123 172 -89
rect 206 -123 244 -89
rect 278 -123 316 -89
rect 350 -123 388 -89
rect 422 -123 460 -89
rect 494 -123 532 -89
rect 566 -123 604 -89
rect 638 -123 676 -89
rect 710 -123 748 -89
rect 782 -123 820 -89
rect 854 -123 892 -89
rect 926 -123 964 -89
rect 998 -123 1036 -89
rect 1070 -123 1108 -89
rect 1142 -123 1180 -89
rect 1214 -123 1252 -89
rect 1286 -123 1324 -89
rect 1358 -123 1396 -89
rect 1430 -123 1468 -89
rect 1502 -123 1540 -89
rect 1574 -123 1612 -89
rect 1646 -123 1684 -89
rect 1718 -123 1756 -89
rect 1790 -123 1828 -89
rect 1862 -123 1900 -89
rect 1934 -123 1972 -89
rect 2006 -123 2044 -89
rect 2078 -123 2116 -89
rect 2150 -123 2188 -89
rect 2222 -123 2260 -89
rect 2294 -123 2332 -89
rect 2366 -123 2404 -89
rect 2438 -123 2476 -89
rect 2510 -123 2548 -89
rect 2582 -123 2620 -89
rect 2654 -123 2692 -89
rect 2726 -123 2764 -89
rect 2798 -123 2836 -89
rect 2870 -123 2900 -89
<< viali >>
rect 148 1527 182 1561
rect 220 1527 254 1561
rect 292 1527 326 1561
rect 364 1527 398 1561
rect 436 1527 470 1561
rect 508 1527 542 1561
rect 580 1527 614 1561
rect 652 1527 686 1561
rect 724 1527 758 1561
rect 796 1527 830 1561
rect 868 1527 902 1561
rect 940 1527 974 1561
rect 1012 1527 1046 1561
rect 1084 1527 1118 1561
rect 1156 1527 1190 1561
rect 1228 1527 1262 1561
rect 1300 1527 1334 1561
rect 1372 1527 1406 1561
rect 1444 1527 1478 1561
rect 1516 1527 1550 1561
rect 1588 1527 1622 1561
rect 1660 1527 1694 1561
rect 1732 1527 1766 1561
rect 1804 1527 1838 1561
rect 1876 1527 1910 1561
rect 1948 1527 1982 1561
rect 2020 1527 2054 1561
rect 2092 1527 2126 1561
rect 2164 1527 2198 1561
rect 2236 1527 2270 1561
rect 2308 1527 2342 1561
rect 2380 1527 2414 1561
rect 2452 1527 2486 1561
rect 2524 1527 2558 1561
rect 2596 1527 2630 1561
rect 2668 1527 2702 1561
rect 2740 1527 2774 1561
rect 2812 1527 2846 1561
rect 2884 1527 2918 1561
rect 2956 1527 2990 1561
rect 3028 1527 3062 1561
rect 3100 1527 3134 1561
rect 3172 1527 3206 1561
rect 3244 1527 3278 1561
rect 3316 1527 3350 1561
rect 3388 1527 3422 1561
rect 3460 1527 3494 1561
rect 3532 1527 3566 1561
rect 3604 1527 3638 1561
rect 3676 1527 3710 1561
rect 3748 1527 3782 1561
rect 3820 1527 3854 1561
rect 3892 1527 3926 1561
rect 3964 1527 3998 1561
rect 4036 1527 4070 1561
rect 4108 1527 4142 1561
rect 4180 1527 4214 1561
rect 4252 1527 4286 1561
rect 4324 1527 4358 1561
rect 4396 1527 4430 1561
rect 4468 1527 4502 1561
rect 4540 1527 4574 1561
rect 4612 1527 4646 1561
rect 4684 1527 4718 1561
rect 4756 1527 4790 1561
rect 4828 1527 4862 1561
rect 4900 1527 4934 1561
rect 4972 1527 5006 1561
rect 5044 1527 5078 1561
rect 5116 1527 5150 1561
rect 5188 1527 5222 1561
rect 5260 1527 5294 1561
rect 5332 1527 5366 1561
rect 5404 1527 5438 1561
rect 5476 1527 5510 1561
rect 172 -123 206 -89
rect 244 -123 278 -89
rect 316 -123 350 -89
rect 388 -123 422 -89
rect 460 -123 494 -89
rect 532 -123 566 -89
rect 604 -123 638 -89
rect 676 -123 710 -89
rect 748 -123 782 -89
rect 820 -123 854 -89
rect 892 -123 926 -89
rect 964 -123 998 -89
rect 1036 -123 1070 -89
rect 1108 -123 1142 -89
rect 1180 -123 1214 -89
rect 1252 -123 1286 -89
rect 1324 -123 1358 -89
rect 1396 -123 1430 -89
rect 1468 -123 1502 -89
rect 1540 -123 1574 -89
rect 1612 -123 1646 -89
rect 1684 -123 1718 -89
rect 1756 -123 1790 -89
rect 1828 -123 1862 -89
rect 1900 -123 1934 -89
rect 1972 -123 2006 -89
rect 2044 -123 2078 -89
rect 2116 -123 2150 -89
rect 2188 -123 2222 -89
rect 2260 -123 2294 -89
rect 2332 -123 2366 -89
rect 2404 -123 2438 -89
rect 2476 -123 2510 -89
rect 2548 -123 2582 -89
rect 2620 -123 2654 -89
rect 2692 -123 2726 -89
rect 2764 -123 2798 -89
rect 2836 -123 2870 -89
<< metal1 >>
rect 106 1561 5552 1597
rect 106 1527 148 1561
rect 182 1527 220 1561
rect 254 1527 292 1561
rect 326 1527 364 1561
rect 398 1527 436 1561
rect 470 1527 508 1561
rect 542 1527 580 1561
rect 614 1527 652 1561
rect 686 1527 724 1561
rect 758 1527 796 1561
rect 830 1527 868 1561
rect 902 1527 940 1561
rect 974 1527 1012 1561
rect 1046 1527 1084 1561
rect 1118 1527 1156 1561
rect 1190 1527 1228 1561
rect 1262 1527 1300 1561
rect 1334 1527 1372 1561
rect 1406 1527 1444 1561
rect 1478 1527 1516 1561
rect 1550 1527 1588 1561
rect 1622 1527 1660 1561
rect 1694 1527 1732 1561
rect 1766 1527 1804 1561
rect 1838 1527 1876 1561
rect 1910 1527 1948 1561
rect 1982 1527 2020 1561
rect 2054 1527 2092 1561
rect 2126 1527 2164 1561
rect 2198 1527 2236 1561
rect 2270 1527 2308 1561
rect 2342 1527 2380 1561
rect 2414 1527 2452 1561
rect 2486 1527 2524 1561
rect 2558 1527 2596 1561
rect 2630 1527 2668 1561
rect 2702 1527 2740 1561
rect 2774 1527 2812 1561
rect 2846 1527 2884 1561
rect 2918 1527 2956 1561
rect 2990 1527 3028 1561
rect 3062 1527 3100 1561
rect 3134 1527 3172 1561
rect 3206 1527 3244 1561
rect 3278 1527 3316 1561
rect 3350 1527 3388 1561
rect 3422 1527 3460 1561
rect 3494 1527 3532 1561
rect 3566 1527 3604 1561
rect 3638 1527 3676 1561
rect 3710 1527 3748 1561
rect 3782 1527 3820 1561
rect 3854 1527 3892 1561
rect 3926 1527 3964 1561
rect 3998 1527 4036 1561
rect 4070 1527 4108 1561
rect 4142 1527 4180 1561
rect 4214 1527 4252 1561
rect 4286 1527 4324 1561
rect 4358 1527 4396 1561
rect 4430 1527 4468 1561
rect 4502 1527 4540 1561
rect 4574 1527 4612 1561
rect 4646 1527 4684 1561
rect 4718 1527 4756 1561
rect 4790 1527 4828 1561
rect 4862 1527 4900 1561
rect 4934 1527 4972 1561
rect 5006 1527 5044 1561
rect 5078 1527 5116 1561
rect 5150 1527 5188 1561
rect 5222 1527 5260 1561
rect 5294 1527 5332 1561
rect 5366 1527 5404 1561
rect 5438 1527 5476 1561
rect 5510 1527 5552 1561
rect 106 1521 5552 1527
rect 325 1447 5333 1521
rect 106 1377 284 1401
rect 106 1325 176 1377
rect 228 1325 284 1377
rect 106 1301 284 1325
rect 325 1061 5333 1255
rect 106 915 284 1015
rect 106 569 5553 869
rect 106 423 284 523
rect 316 183 2726 377
rect 166 113 284 137
rect 166 61 176 113
rect 228 61 284 113
rect 166 37 284 61
rect 316 -83 2726 -9
rect 106 -89 5552 -83
rect 106 -123 172 -89
rect 206 -123 244 -89
rect 278 -123 316 -89
rect 350 -123 388 -89
rect 422 -123 460 -89
rect 494 -123 532 -89
rect 566 -123 604 -89
rect 638 -123 676 -89
rect 710 -123 748 -89
rect 782 -123 820 -89
rect 854 -123 892 -89
rect 926 -123 964 -89
rect 998 -123 1036 -89
rect 1070 -123 1108 -89
rect 1142 -123 1180 -89
rect 1214 -123 1252 -89
rect 1286 -123 1324 -89
rect 1358 -123 1396 -89
rect 1430 -123 1468 -89
rect 1502 -123 1540 -89
rect 1574 -123 1612 -89
rect 1646 -123 1684 -89
rect 1718 -123 1756 -89
rect 1790 -123 1828 -89
rect 1862 -123 1900 -89
rect 1934 -123 1972 -89
rect 2006 -123 2044 -89
rect 2078 -123 2116 -89
rect 2150 -123 2188 -89
rect 2222 -123 2260 -89
rect 2294 -123 2332 -89
rect 2366 -123 2404 -89
rect 2438 -123 2476 -89
rect 2510 -123 2548 -89
rect 2582 -123 2620 -89
rect 2654 -123 2692 -89
rect 2726 -123 2764 -89
rect 2798 -123 2836 -89
rect 2870 -123 5552 -89
rect 106 -159 5552 -123
<< via1 >>
rect 176 1325 228 1377
rect 176 61 228 113
<< metal2 >>
rect 176 1377 228 1411
rect 176 113 228 1325
rect 176 27 228 61
use sky130_fd_pr__nfet_01v8_PHNS9E  sky130_fd_pr__nfet_01v8_PHNS9E_0
timestamp 1750100919
transform 0 1 1521 -1 0 87
box -236 -1405 236 1405
use sky130_fd_pr__pfet_01v8_D9QVK3  sky130_fd_pr__pfet_01v8_D9QVK3_0
timestamp 1750100919
transform 0 1 2829 -1 0 965
box -246 -2723 246 2723
use sky130_fd_pr__pfet_01v8_D9QVK3  XM1
timestamp 1750100919
transform 0 1 2829 -1 0 1351
box -246 -2723 246 2723
use sky130_fd_pr__nfet_01v8_PHNS9E  XM3
timestamp 1750100919
transform 0 1 1521 -1 0 473
box -236 -1405 236 1405
<< labels >>
flabel metal1 s 118 1554 124 1560 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 119 1347 125 1353 0 FreeSans 500 0 0 0 IN
port 2 nsew
flabel metal1 s 122 961 128 967 0 FreeSans 500 0 0 0 CKB
port 3 nsew
flabel metal1 s 119 469 125 475 0 FreeSans 500 0 0 0 CK
port 4 nsew
flabel metal1 s 119 -127 125 -121 0 FreeSans 500 0 0 0 VSS
port 5 nsew
flabel metal1 s 5515 700 5521 706 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
