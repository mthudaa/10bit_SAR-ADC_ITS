magic
tech sky130A
magscale 1 2
timestamp 1749499571
<< dnwell >>
rect -10590 44364 -3793 76025
rect -2373 1624 49198 118766
rect 50479 58365 56127 62017
<< metal1 >>
rect 614 61819 624 61900
rect -4692 61563 624 61819
rect 44492 61563 49994 61900
rect 50046 61563 50056 61900
rect 49984 60282 49994 60334
rect 50046 60316 50056 60334
rect 50046 60282 50737 60316
rect 49984 60048 49994 60100
rect 50046 60066 50538 60100
rect 50046 60048 50056 60066
rect -4704 58571 624 58827
rect 614 58490 624 58571
rect 44492 58490 49994 58827
rect 50046 58490 50056 58827
<< via1 >>
rect 624 61563 44492 61900
rect 49994 61563 50046 61900
rect 49994 60282 50046 60334
rect 49994 60048 50046 60100
rect 624 58490 44492 58827
rect 49994 58490 50046 58827
<< metal2 >>
rect 624 61900 44492 61910
rect 624 61553 44492 61563
rect 49994 61900 50046 61910
rect 49994 60334 50046 61563
rect 49994 60272 50046 60282
rect 49994 60100 50046 60110
rect 624 58827 44492 58837
rect 624 58480 44492 58490
rect 49994 58827 50046 60048
rect 49994 58480 50046 58490
<< via2 >>
rect 624 61563 44492 61900
rect 624 58490 44492 58827
<< metal3 >>
rect 614 61900 44502 61905
rect 614 61563 624 61900
rect 44492 61563 44502 61900
rect 614 61558 44502 61563
rect 614 58827 44502 58832
rect 614 58490 624 58827
rect 44492 58490 44502 58827
rect 614 58485 44502 58490
<< via3 >>
rect 624 61563 44492 61900
rect 624 58490 44492 58827
<< metal4 >>
rect 623 61900 44493 61901
rect 623 61563 624 61900
rect 44492 61563 44493 61900
rect 623 61562 44493 61563
rect 623 58827 44493 58828
rect 623 58490 624 58827
rect 44492 58490 44493 58827
rect 623 58489 44493 58490
use cdac  cdac_0
timestamp 1749497408
transform 1 0 -1274 0 1 2329
box -1099 -705 50472 116437
use sar10b  sar10b_0
timestamp 1749411235
transform 1 0 56915 0 1 44953
box 0 0 11722 28874
use tdc  tdc_0
timestamp 1749411235
transform 1 0 50703 0 1 59011
box -224 -646 5424 3006
use th_dif_sw  th_dif_sw_0
timestamp 1749411235
transform 0 -1 -4206 1 0 44365
box -1 -413 31660 6384
<< end >>
