magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< metal1 >>
rect -228 1377 61 1400
rect -228 1325 -194 1377
rect -142 1325 61 1377
rect -228 1302 61 1325
rect -1628 1224 42 1228
rect -1628 1172 -1594 1224
rect -1542 1172 42 1224
rect -1628 1168 42 1172
rect -628 1073 42 1077
rect -628 1021 -594 1073
rect -542 1021 42 1073
rect -628 1017 42 1021
rect -828 897 51 901
rect -828 845 -794 897
rect -742 845 51 897
rect -828 841 51 845
rect -428 711 116 734
rect -428 659 -394 711
rect -342 659 116 711
rect -428 636 116 659
rect -1028 349 45 353
rect -1028 297 -994 349
rect -942 297 45 349
rect -1028 293 45 297
rect -1228 194 44 198
rect -1228 142 -1194 194
rect -1142 142 44 194
rect -1228 138 44 142
rect -228 39 91 68
rect -228 -13 -194 39
rect -142 -13 91 39
rect -228 -25 91 -13
rect -228 -77 -194 -25
rect -142 -77 91 -25
rect -228 -106 91 -77
rect -628 -636 67 -612
rect -628 -688 -594 -636
rect -542 -688 67 -636
rect -628 -712 67 -688
rect 1539 -786 3365 -758
rect 1539 -838 3279 -786
rect 3331 -838 3365 -786
rect 1539 -850 3365 -838
rect 1539 -902 3279 -850
rect 3331 -902 3365 -850
rect 1539 -914 3365 -902
rect 1539 -966 3279 -914
rect 3331 -966 3365 -914
rect 1539 -978 3365 -966
rect 1539 -1030 3279 -978
rect 3331 -1030 3365 -978
rect 1539 -1058 3365 -1030
rect -828 -1128 -18 -1104
rect -828 -1180 -794 -1128
rect -742 -1180 -18 -1128
rect -828 -1204 -18 -1180
rect -1828 -1514 49 -1490
rect -1828 -1566 -1794 -1514
rect -1742 -1566 49 -1514
rect -1828 -1590 49 -1566
rect -428 -1728 59 -1710
rect -428 -1780 -394 -1728
rect -342 -1780 59 -1728
rect -428 -1792 59 -1780
rect -428 -1844 -394 -1792
rect -342 -1844 59 -1792
rect -428 -1862 59 -1844
rect 3245 -1893 3365 -1868
rect 3245 -1902 3279 -1893
rect -27 -2006 93 -1986
rect -27 -2058 7 -2006
rect 59 -2058 93 -2006
rect -27 -2078 93 -2058
rect 1115 -2162 1149 -1903
rect 3018 -1936 3279 -1902
rect 3245 -1945 3279 -1936
rect 3331 -1945 3365 -1893
rect 3245 -1970 3365 -1945
rect 3045 -2006 3165 -1986
rect 3045 -2058 3079 -2006
rect 3131 -2058 3165 -2006
rect 3045 -2078 3165 -2058
rect -228 -2220 57 -2202
rect -228 -2272 -194 -2220
rect -142 -2272 57 -2220
rect -228 -2284 57 -2272
rect -228 -2336 -194 -2284
rect -142 -2336 57 -2284
rect -228 -2354 57 -2336
rect 3245 -2385 3365 -2360
rect 3245 -2394 3279 -2385
rect 3010 -2428 3279 -2394
rect 3245 -2437 3279 -2428
rect 3331 -2437 3365 -2385
rect 3245 -2462 3365 -2437
rect -1228 -2498 93 -2478
rect -1228 -2550 -1194 -2498
rect -1142 -2550 7 -2498
rect 59 -2550 93 -2498
rect -1228 -2570 93 -2550
rect 3045 -2498 3165 -2478
rect 3045 -2550 3079 -2498
rect 3131 -2550 3165 -2498
rect 3045 -2570 3165 -2550
rect -1428 -2611 -1308 -2586
rect -1428 -2663 -1394 -2611
rect -1342 -2620 -1308 -2611
rect -1342 -2654 126 -2620
rect -1342 -2663 -1308 -2654
rect -1428 -2688 -1308 -2663
rect -428 -2712 51 -2694
rect -428 -2764 -394 -2712
rect -342 -2764 51 -2712
rect -428 -2776 51 -2764
rect -428 -2828 -394 -2776
rect -342 -2828 51 -2776
rect -428 -2846 51 -2828
rect -27 -2990 93 -2970
rect -27 -3042 7 -2990
rect 59 -3042 93 -2990
rect -27 -3062 93 -3042
rect -1428 -3103 -1308 -3078
rect -1428 -3155 -1394 -3103
rect -1342 -3112 -1308 -3103
rect -1342 -3146 109 -3112
rect 1116 -3146 1150 -2902
rect 3045 -2990 3165 -2970
rect 3045 -3042 3079 -2990
rect 3131 -3042 3165 -2990
rect 3045 -3062 3165 -3042
rect -1342 -3155 -1308 -3146
rect -1428 -3180 -1308 -3155
rect -228 -3198 84 -3186
rect -228 -3250 -194 -3198
rect -142 -3250 84 -3198
rect -228 -3262 84 -3250
<< via1 >>
rect -194 1325 -142 1377
rect -1594 1172 -1542 1224
rect -594 1021 -542 1073
rect -794 845 -742 897
rect -394 659 -342 711
rect -994 297 -942 349
rect -1194 142 -1142 194
rect -194 -13 -142 39
rect -194 -77 -142 -25
rect -594 -688 -542 -636
rect 3279 -838 3331 -786
rect 3279 -902 3331 -850
rect 3279 -966 3331 -914
rect 3279 -1030 3331 -978
rect -794 -1180 -742 -1128
rect -1794 -1566 -1742 -1514
rect -394 -1780 -342 -1728
rect -394 -1844 -342 -1792
rect 7 -2058 59 -2006
rect 3279 -1945 3331 -1893
rect 3079 -2058 3131 -2006
rect -194 -2272 -142 -2220
rect -194 -2336 -142 -2284
rect 3279 -2437 3331 -2385
rect -1194 -2550 -1142 -2498
rect 7 -2550 59 -2498
rect 3079 -2550 3131 -2498
rect -1394 -2663 -1342 -2611
rect -394 -2764 -342 -2712
rect -394 -2828 -342 -2776
rect 7 -3042 59 -2990
rect -1394 -3155 -1342 -3103
rect 3079 -3042 3131 -2990
rect -194 -3250 -142 -3198
<< metal2 >>
rect -1818 -1514 -1718 1400
rect -1818 -1566 -1794 -1514
rect -1742 -1566 -1718 -1514
rect -1818 -3272 -1718 -1566
rect -1618 1224 -1518 1400
rect -1618 1172 -1594 1224
rect -1542 1172 -1518 1224
rect -1618 -3272 -1518 1172
rect -1418 -2611 -1318 1400
rect -1418 -2663 -1394 -2611
rect -1342 -2663 -1318 -2611
rect -1418 -3103 -1318 -2663
rect -1418 -3155 -1394 -3103
rect -1342 -3155 -1318 -3103
rect -1418 -3272 -1318 -3155
rect -1218 194 -1118 1400
rect -1218 142 -1194 194
rect -1142 142 -1118 194
rect -1218 -2498 -1118 142
rect -1218 -2550 -1194 -2498
rect -1142 -2550 -1118 -2498
rect -1218 -3272 -1118 -2550
rect -1018 349 -918 1400
rect -1018 297 -994 349
rect -942 297 -918 349
rect -1018 -2004 -918 297
rect -1018 -2060 -996 -2004
rect -940 -2060 -918 -2004
rect -1018 -3272 -918 -2060
rect -818 897 -718 1400
rect -818 845 -794 897
rect -742 845 -718 897
rect -818 -1128 -718 845
rect -818 -1180 -794 -1128
rect -742 -1180 -718 -1128
rect -818 -3272 -718 -1180
rect -618 1073 -518 1400
rect -618 1021 -594 1073
rect -542 1021 -518 1073
rect -618 -636 -518 1021
rect -618 -688 -594 -636
rect -542 -688 -518 -636
rect -618 -3272 -518 -688
rect -418 711 -318 1400
rect -418 659 -394 711
rect -342 659 -318 711
rect -418 -1728 -318 659
rect -418 -1780 -394 -1728
rect -342 -1780 -318 -1728
rect -418 -1792 -318 -1780
rect -418 -1844 -394 -1792
rect -342 -1844 -318 -1792
rect -418 -2712 -318 -1844
rect -418 -2764 -394 -2712
rect -342 -2764 -318 -2712
rect -418 -2776 -318 -2764
rect -418 -2828 -394 -2776
rect -342 -2828 -318 -2776
rect -418 -3272 -318 -2828
rect -218 1377 -118 1410
rect -218 1325 -194 1377
rect -142 1325 -118 1377
rect -218 39 -118 1325
rect -218 -13 -194 39
rect -142 -13 -118 39
rect -218 -25 -118 -13
rect -218 -77 -194 -25
rect -142 -77 -118 -25
rect -218 -2220 -118 -77
rect 3255 -786 3355 -748
rect 3255 -838 3279 -786
rect 3331 -838 3355 -786
rect 3255 -850 3355 -838
rect 3255 -902 3279 -850
rect 3331 -902 3355 -850
rect 3255 -914 3355 -902
rect 3255 -966 3279 -914
rect 3331 -966 3355 -914
rect 3255 -978 3355 -966
rect 3255 -1030 3279 -978
rect 3331 -1030 3355 -978
rect 3255 -1893 3355 -1030
rect 3255 -1945 3279 -1893
rect 3331 -1945 3355 -1893
rect -218 -2272 -194 -2220
rect -142 -2272 -118 -2220
rect -218 -2284 -118 -2272
rect -218 -2336 -194 -2284
rect -142 -2336 -118 -2284
rect -218 -3198 -118 -2336
rect -17 -2006 83 -1976
rect -17 -2058 7 -2006
rect 59 -2058 83 -2006
rect -17 -2498 83 -2058
rect -17 -2550 7 -2498
rect 59 -2550 83 -2498
rect -17 -2990 83 -2550
rect -17 -3042 7 -2990
rect 59 -3042 83 -2990
rect -17 -3072 83 -3042
rect 3055 -2004 3155 -1976
rect 3055 -2060 3077 -2004
rect 3133 -2060 3155 -2004
rect 3055 -2498 3155 -2060
rect 3255 -2385 3355 -1945
rect 3255 -2437 3279 -2385
rect 3331 -2437 3355 -2385
rect 3255 -2472 3355 -2437
rect 3055 -2550 3079 -2498
rect 3131 -2550 3155 -2498
rect 3055 -2990 3155 -2550
rect 3055 -3042 3079 -2990
rect 3131 -3042 3155 -2990
rect 3055 -3072 3155 -3042
rect -218 -3250 -194 -3198
rect -142 -3250 -118 -3198
rect -218 -3272 -118 -3250
<< via2 >>
rect -996 -2060 -940 -2004
rect 3077 -2006 3133 -2004
rect 3077 -2058 3079 -2006
rect 3079 -2058 3131 -2006
rect 3131 -2058 3133 -2006
rect 3077 -2060 3133 -2058
<< metal3 >>
rect -1028 -1986 -908 -1981
rect 3045 -1986 3165 -1981
rect -1028 -2004 3165 -1986
rect -1028 -2060 -996 -2004
rect -940 -2060 3077 -2004
rect 3133 -2060 3165 -2004
rect -1028 -2078 3165 -2060
rect -1028 -2083 -908 -2078
rect 3045 -2083 3165 -2078
use dac_sw_9  dac_sw_9_0
timestamp 1750100919
transform 1 0 -124 0 -1 -189
box 106 -159 2128 1597
use nooverlap_clk  nooverlap_clk_0
timestamp 1750100919
transform -1 0 2909 0 1 4745
box -701 -4775 2927 -3345
use tg_sw_9  tg_sw_9_0
timestamp 1750100919
transform -1 0 3101 0 1 -2225
box -53 -53 3119 439
use tg_sw_9  tg_sw_9_1
timestamp 1750100919
transform 1 0 36 0 -1 -2331
box -53 -53 3119 439
use tg_sw_9  tg_sw_9_9
timestamp 1750100919
transform -1 0 3102 0 1 -3209
box -53 -53 3119 439
<< labels >>
flabel metal1 s 3036 -973 3136 -839 0 FreeSans 500 0 0 0 DAC_OUT
port 1 nsew
flabel metal2 s -182 -393 -142 -353 0 FreeSans 600 0 0 0 VSSA
port 2 nsew
flabel metal2 s -393 -382 -353 -342 0 FreeSans 600 0 0 0 VDDA
port 3 nsew
flabel metal2 s -1384 -382 -1344 -342 0 FreeSans 600 0 0 0 VCM
port 4 nsew
flabel metal2 s -1593 -388 -1553 -348 0 FreeSans 600 0 0 0 CKI
port 5 nsew
flabel metal2 s -1786 -378 -1746 -338 0 FreeSans 600 0 0 0 BI
port 6 nsew
<< end >>
