magic
tech sky130A
magscale 1 2
timestamp 1748794220
<< viali >>
rect 142 1527 5516 1561
rect 142 -123 2900 -89
<< metal1 >>
rect 106 1561 5552 1597
rect 106 1527 142 1561
rect 5516 1527 5552 1561
rect 106 1521 5552 1527
rect 325 1447 5333 1521
rect 106 1301 176 1401
rect 228 1301 284 1401
rect 325 1061 5333 1255
rect 106 915 284 1015
rect 106 569 5553 869
rect 106 423 284 523
rect 316 183 2726 377
rect 166 37 176 137
rect 228 37 284 137
rect 316 -83 2726 -9
rect 106 -89 5552 -83
rect 106 -123 142 -89
rect 2900 -123 5552 -89
rect 106 -159 5552 -123
<< via1 >>
rect 176 1301 228 1401
rect 176 37 228 137
<< metal2 >>
rect 176 1401 228 1411
rect 176 137 228 1301
rect 176 27 228 37
use sky130_fd_pr__nfet_01v8_PHNS9E  sky130_fd_pr__nfet_01v8_PHNS9E_0
timestamp 1746381332
transform 0 1 1521 -1 0 87
box -246 -1415 246 1415
use sky130_fd_pr__pfet_01v8_D9QVK3  sky130_fd_pr__pfet_01v8_D9QVK3_0
timestamp 1746381332
transform 0 1 2829 -1 0 965
box -246 -2723 246 2723
use sky130_fd_pr__pfet_01v8_D9QVK3  XM1
timestamp 1746381332
transform 0 1 2829 -1 0 1351
box -246 -2723 246 2723
use sky130_fd_pr__nfet_01v8_PHNS9E  XM3
timestamp 1746381332
transform 0 1 1521 -1 0 473
box -246 -1415 246 1415
<< labels >>
flabel metal1 118 1554 124 1560 0 FreeSans 400 0 0 0 VDD
port 0 nsew
flabel metal1 119 1347 125 1353 0 FreeSans 400 0 0 0 IN
port 1 nsew
flabel metal1 122 961 128 967 0 FreeSans 400 0 0 0 CKB
port 2 nsew
flabel metal1 119 469 125 475 0 FreeSans 400 0 0 0 CK
port 3 nsew
flabel metal1 119 -127 125 -121 0 FreeSans 400 0 0 0 VSS
port 4 nsew
flabel metal1 5515 700 5521 706 0 FreeSans 400 0 0 0 OUT
port 6 nsew
<< end >>
