magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect 9509 4631 9667 6177
rect 10990 1253 11024 1282
rect 10990 1157 11024 1219
rect 10990 1061 11024 1123
rect 10990 965 11024 1027
rect 10990 869 11024 931
rect 10990 773 11024 835
rect 10990 677 11024 739
rect 10990 581 11024 643
rect 10990 485 11024 547
rect 10990 389 11024 451
rect 10990 293 11024 355
rect 10990 197 11024 259
rect 10959 163 10990 197
<< viali >>
rect 10990 1219 11024 1253
rect 10990 1123 11024 1157
rect 10990 1027 11024 1061
rect 10990 931 11024 965
rect 10990 835 11024 869
rect 10990 739 11024 773
rect 10990 643 11024 677
rect 10990 547 11024 581
rect 10990 451 11024 485
rect 10990 355 11024 389
rect 10990 259 11024 293
rect 10990 163 11024 197
<< metal1 >>
rect 9509 4631 9667 6177
rect 10801 2417 10811 2469
rect 10863 2417 10873 2469
rect 12803 2063 14615 2069
rect 12803 1819 12819 2063
rect 14599 1819 14615 2063
rect 12803 1813 14615 1819
rect 10724 1761 13069 1813
rect 12813 1666 13069 1761
rect 13325 1650 13581 1813
rect 13837 1666 14093 1813
rect 14349 1666 14605 1813
rect 10959 1253 11055 1282
rect 10959 1219 10990 1253
rect 11024 1219 11055 1253
rect 10959 1157 11055 1219
rect 10959 1123 10990 1157
rect 11024 1123 11055 1157
rect 10959 1061 11055 1123
rect 10959 1027 10990 1061
rect 11024 1027 11055 1061
rect 10959 965 11055 1027
rect 10959 931 10990 965
rect 11024 931 11055 965
rect 10959 869 11055 931
rect 10959 835 10990 869
rect 11024 835 11055 869
rect 10959 773 11055 835
rect 10959 739 10990 773
rect 11024 739 11055 773
rect 10801 668 10811 720
rect 10863 668 10873 720
rect 10959 677 11055 739
rect 10959 643 10990 677
rect 11024 643 11055 677
rect 10959 581 11055 643
rect 9667 197 9825 563
rect 10959 547 10990 581
rect 11024 547 11055 581
rect 10959 485 11055 547
rect 10959 451 10990 485
rect 11024 451 11055 485
rect 10959 389 11055 451
rect 10959 355 10990 389
rect 11024 355 11055 389
rect 10959 293 11055 355
rect 10959 259 10990 293
rect 11024 259 11055 293
rect 10959 197 11055 259
rect 10959 163 10990 197
rect 11024 163 11055 197
rect 10959 132 11055 163
rect 11789 388 12045 568
rect 12301 388 12557 568
rect 12813 388 13069 568
rect 13325 388 13581 568
rect 13837 388 14093 568
rect 14349 388 14605 568
rect 11789 132 14605 388
<< via1 >>
rect 10811 2417 10863 2469
rect 12819 1819 14599 2063
rect 10811 668 10863 720
<< metal2 >>
rect 12813 6223 14605 6253
rect 12813 6007 12841 6223
rect 14577 6007 14605 6223
rect 12813 5977 14605 6007
rect 10811 2469 10863 2479
rect 10811 1165 10863 2417
rect 12813 2063 14605 2079
rect 12813 1819 12819 2063
rect 14599 1819 14605 2063
rect 12813 1803 14605 1819
rect 10811 1113 11102 1165
rect 10811 797 11095 849
rect 10811 720 10863 797
rect 10811 36 10863 668
rect 10811 -16 15509 36
rect 10679 -66 10735 -56
rect 10801 -66 10857 -56
rect 10735 -120 10801 -68
rect 10679 -132 10735 -122
rect 10857 -120 15509 -68
rect 10801 -132 10857 -122
<< via2 >>
rect 12841 6007 14577 6223
rect 12841 1833 14577 2049
rect 10679 -122 10735 -66
rect 10801 -122 10857 -66
<< metal3 >>
rect 12803 6223 14615 6248
rect 12803 6007 12841 6223
rect 14577 6007 14615 6223
rect 12803 5982 14615 6007
rect 10735 -61 10801 4166
rect 12813 2074 13069 5982
rect 13325 2074 13581 5982
rect 13837 2074 14093 5982
rect 14349 2074 14605 5982
rect 12803 2049 14615 2074
rect 12803 1833 12841 2049
rect 14577 1833 14615 2049
rect 12803 1808 14615 1833
rect 10669 -66 10867 -61
rect 10669 -122 10679 -66
rect 10735 -122 10801 -66
rect 10857 -122 10867 -66
rect 10669 -127 10867 -122
use bootstrap  bootstrap_0
timestamp 1750100919
transform 1 0 9430 0 1 4264
box -9799 -4132 4107 1978
use th_sw_main  th_sw_main_0
timestamp 1750100919
transform 0 -1 13127 1 0 -16
box 584 -2382 1726 2168
<< labels >>
flabel metal1 s 9562 5504 9596 5538 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 9730 378 9764 412 0 FreeSans 500 0 0 0 VSS
port 2 nsew
flabel metal3 s 13156 6124 13190 6158 0 FreeSans 500 0 0 0 IN
port 3 nsew
flabel metal1 s 13165 281 13199 315 0 FreeSans 500 0 0 0 OUT
port 4 nsew
flabel metal2 s 15468 -7 15502 27 0 FreeSans 500 0 0 0 CK
port 5 nsew
flabel metal2 s 15467 -109 15501 -75 0 FreeSans 500 0 0 0 CKB
port 6 nsew
<< end >>
