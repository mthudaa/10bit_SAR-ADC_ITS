magic
tech sky130A
magscale 1 2
timestamp 1749310734
<< error_p >>
rect -29 -86 29 -80
rect -29 -120 -17 -86
rect -29 -126 29 -120
<< nwell >>
rect -211 -259 211 259
<< pmos >>
rect -15 -39 15 111
<< pdiff >>
rect -73 99 -15 111
rect -73 -27 -61 99
rect -27 -27 -15 99
rect -73 -39 -15 -27
rect 15 99 73 111
rect 15 -27 27 99
rect 61 -27 73 99
rect 15 -39 73 -27
<< pdiffc >>
rect -61 -27 -27 99
rect 27 -27 61 99
<< nsubdiff >>
rect -175 189 -79 223
rect 79 189 175 223
rect -175 126 -141 189
rect 141 126 175 189
rect -175 -189 -141 -126
rect 141 -189 175 -126
rect -175 -223 -79 -189
rect 79 -223 175 -189
<< nsubdiffcont >>
rect -79 189 79 223
rect -175 -126 -141 126
rect 141 -126 175 126
rect -79 -223 79 -189
<< poly >>
rect -15 111 15 137
rect -15 -70 15 -39
rect -33 -86 33 -70
rect -33 -120 -17 -86
rect 17 -120 33 -86
rect -33 -136 33 -120
<< polycont >>
rect -17 -120 17 -86
<< locali >>
rect -175 189 -79 223
rect 79 189 175 223
rect -175 126 -141 189
rect 141 126 175 189
rect -61 99 -27 115
rect -61 -43 -27 -27
rect 27 99 61 115
rect 27 -43 61 -27
rect -33 -120 -17 -86
rect 17 -120 33 -86
rect -175 -189 -141 -126
rect 141 -189 175 -126
rect -175 -223 -79 -189
rect 79 -223 175 -189
<< viali >>
rect -61 -27 -27 99
rect 27 -27 61 99
rect -17 -120 17 -86
<< metal1 >>
rect -67 99 -21 111
rect -67 -27 -61 99
rect -27 -27 -21 99
rect -67 -39 -21 -27
rect 21 99 67 111
rect 21 -27 27 99
rect 61 -27 67 99
rect 21 -39 67 -27
rect -29 -86 29 -80
rect -29 -120 -17 -86
rect 17 -120 29 -86
rect -29 -126 29 -120
<< properties >>
string FIXED_BBOX -158 -206 158 206
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.75 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
