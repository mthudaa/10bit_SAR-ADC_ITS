magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect -17 369 -15 403
rect 19 369 57 403
rect 91 369 129 403
rect 163 369 201 403
rect 235 369 273 403
rect 307 369 345 403
rect 379 369 417 403
rect 451 369 489 403
rect 523 369 561 403
rect 595 369 633 403
rect 667 369 705 403
rect 739 369 777 403
rect 811 369 849 403
rect 883 369 921 403
rect 955 369 993 403
rect 1027 369 1065 403
rect 1099 369 1137 403
rect 1171 369 1209 403
rect 1243 369 1281 403
rect 1315 369 1353 403
rect 1387 369 1425 403
rect 1459 369 1497 403
rect 1531 369 1569 403
rect 1603 369 1641 403
rect 1675 369 1713 403
rect 1747 369 1785 403
rect 1819 369 1857 403
rect 1891 369 1929 403
rect 1963 369 2001 403
rect 2035 369 2073 403
rect 2107 369 2145 403
rect 2179 369 2217 403
rect 2251 369 2289 403
rect 2323 369 2361 403
rect 2395 369 2433 403
rect 2467 369 2505 403
rect 2539 369 2577 403
rect 2611 369 2649 403
rect 2683 369 2721 403
rect 2755 369 2793 403
rect 2827 369 2865 403
rect 2899 369 2937 403
rect 2971 369 3009 403
rect 3043 369 3081 403
rect 3115 369 3153 403
rect 3187 369 3225 403
rect 3259 369 3297 403
rect 3331 369 3369 403
rect 3403 369 3441 403
rect 3475 369 3513 403
rect 3547 369 3585 403
rect 3619 369 3657 403
rect 3691 369 3729 403
rect 3763 369 3801 403
rect 3835 369 3873 403
rect 3907 369 3945 403
rect 3979 369 4017 403
rect 4051 369 4089 403
rect 4123 369 4161 403
rect 4195 369 4233 403
rect 4267 369 4305 403
rect 4339 369 4377 403
rect 4411 369 4449 403
rect 4483 369 4521 403
rect 4555 369 4593 403
rect 4627 369 4665 403
rect 4699 369 4737 403
rect 4771 369 4809 403
rect 4843 369 4881 403
rect 4915 369 4953 403
rect 4987 369 5025 403
rect 5059 369 5097 403
rect 5131 369 5169 403
rect 5203 369 5241 403
rect 5275 369 5313 403
rect 5347 369 5385 403
rect 5419 369 5457 403
rect 5491 369 5529 403
rect 5563 369 5601 403
rect 5635 369 5673 403
rect 5707 369 5745 403
rect 5779 369 5817 403
rect 5851 369 5889 403
rect 5923 369 5961 403
rect 5995 369 6033 403
rect 6067 369 6105 403
rect 6139 369 6177 403
rect 6211 369 6213 403
rect 6285 -17 6309 17
rect 6343 -17 6381 17
rect 6415 -17 6453 17
rect 6487 -17 6525 17
rect 6559 -17 6597 17
rect 6631 -17 6669 17
rect 6703 -17 6741 17
rect 6775 -17 6813 17
rect 6847 -17 6885 17
rect 6919 -17 6957 17
rect 6991 -17 7029 17
rect 7063 -17 7101 17
rect 7135 -17 7173 17
rect 7207 -17 7245 17
rect 7279 -17 7317 17
rect 7351 -17 7389 17
rect 7423 -17 7461 17
rect 7495 -17 7533 17
rect 7567 -17 7605 17
rect 7639 -17 7677 17
rect 7711 -17 7749 17
rect 7783 -17 7821 17
rect 7855 -17 7893 17
rect 7927 -17 7965 17
rect 7999 -17 8037 17
rect 8071 -17 8109 17
rect 8143 -17 8181 17
rect 8215 -17 8253 17
rect 8287 -17 8325 17
rect 8359 -17 8397 17
rect 8431 -17 8469 17
rect 8503 -17 8541 17
rect 8575 -17 8613 17
rect 8647 -17 8685 17
rect 8719 -17 8757 17
rect 8791 -17 8829 17
rect 8863 -17 8901 17
rect 8935 -17 8973 17
rect 9007 -17 9045 17
rect 9079 -17 9117 17
rect 9151 -17 9189 17
rect 9223 -17 9261 17
rect 9295 -17 9333 17
rect 9367 -17 9405 17
rect 9439 -17 9463 17
<< viali >>
rect -15 369 19 403
rect 57 369 91 403
rect 129 369 163 403
rect 201 369 235 403
rect 273 369 307 403
rect 345 369 379 403
rect 417 369 451 403
rect 489 369 523 403
rect 561 369 595 403
rect 633 369 667 403
rect 705 369 739 403
rect 777 369 811 403
rect 849 369 883 403
rect 921 369 955 403
rect 993 369 1027 403
rect 1065 369 1099 403
rect 1137 369 1171 403
rect 1209 369 1243 403
rect 1281 369 1315 403
rect 1353 369 1387 403
rect 1425 369 1459 403
rect 1497 369 1531 403
rect 1569 369 1603 403
rect 1641 369 1675 403
rect 1713 369 1747 403
rect 1785 369 1819 403
rect 1857 369 1891 403
rect 1929 369 1963 403
rect 2001 369 2035 403
rect 2073 369 2107 403
rect 2145 369 2179 403
rect 2217 369 2251 403
rect 2289 369 2323 403
rect 2361 369 2395 403
rect 2433 369 2467 403
rect 2505 369 2539 403
rect 2577 369 2611 403
rect 2649 369 2683 403
rect 2721 369 2755 403
rect 2793 369 2827 403
rect 2865 369 2899 403
rect 2937 369 2971 403
rect 3009 369 3043 403
rect 3081 369 3115 403
rect 3153 369 3187 403
rect 3225 369 3259 403
rect 3297 369 3331 403
rect 3369 369 3403 403
rect 3441 369 3475 403
rect 3513 369 3547 403
rect 3585 369 3619 403
rect 3657 369 3691 403
rect 3729 369 3763 403
rect 3801 369 3835 403
rect 3873 369 3907 403
rect 3945 369 3979 403
rect 4017 369 4051 403
rect 4089 369 4123 403
rect 4161 369 4195 403
rect 4233 369 4267 403
rect 4305 369 4339 403
rect 4377 369 4411 403
rect 4449 369 4483 403
rect 4521 369 4555 403
rect 4593 369 4627 403
rect 4665 369 4699 403
rect 4737 369 4771 403
rect 4809 369 4843 403
rect 4881 369 4915 403
rect 4953 369 4987 403
rect 5025 369 5059 403
rect 5097 369 5131 403
rect 5169 369 5203 403
rect 5241 369 5275 403
rect 5313 369 5347 403
rect 5385 369 5419 403
rect 5457 369 5491 403
rect 5529 369 5563 403
rect 5601 369 5635 403
rect 5673 369 5707 403
rect 5745 369 5779 403
rect 5817 369 5851 403
rect 5889 369 5923 403
rect 5961 369 5995 403
rect 6033 369 6067 403
rect 6105 369 6139 403
rect 6177 369 6211 403
rect 6309 -17 6343 17
rect 6381 -17 6415 17
rect 6453 -17 6487 17
rect 6525 -17 6559 17
rect 6597 -17 6631 17
rect 6669 -17 6703 17
rect 6741 -17 6775 17
rect 6813 -17 6847 17
rect 6885 -17 6919 17
rect 6957 -17 6991 17
rect 7029 -17 7063 17
rect 7101 -17 7135 17
rect 7173 -17 7207 17
rect 7245 -17 7279 17
rect 7317 -17 7351 17
rect 7389 -17 7423 17
rect 7461 -17 7495 17
rect 7533 -17 7567 17
rect 7605 -17 7639 17
rect 7677 -17 7711 17
rect 7749 -17 7783 17
rect 7821 -17 7855 17
rect 7893 -17 7927 17
rect 7965 -17 7999 17
rect 8037 -17 8071 17
rect 8109 -17 8143 17
rect 8181 -17 8215 17
rect 8253 -17 8287 17
rect 8325 -17 8359 17
rect 8397 -17 8431 17
rect 8469 -17 8503 17
rect 8541 -17 8575 17
rect 8613 -17 8647 17
rect 8685 -17 8719 17
rect 8757 -17 8791 17
rect 8829 -17 8863 17
rect 8901 -17 8935 17
rect 8973 -17 9007 17
rect 9045 -17 9079 17
rect 9117 -17 9151 17
rect 9189 -17 9223 17
rect 9261 -17 9295 17
rect 9333 -17 9367 17
rect 9405 -17 9439 17
<< metal1 >>
rect -53 403 9499 439
rect -53 369 -15 403
rect 19 369 57 403
rect 91 369 129 403
rect 163 369 201 403
rect 235 369 273 403
rect 307 369 345 403
rect 379 369 417 403
rect 451 369 489 403
rect 523 369 561 403
rect 595 369 633 403
rect 667 369 705 403
rect 739 369 777 403
rect 811 369 849 403
rect 883 369 921 403
rect 955 369 993 403
rect 1027 369 1065 403
rect 1099 369 1137 403
rect 1171 369 1209 403
rect 1243 369 1281 403
rect 1315 369 1353 403
rect 1387 369 1425 403
rect 1459 369 1497 403
rect 1531 369 1569 403
rect 1603 369 1641 403
rect 1675 369 1713 403
rect 1747 369 1785 403
rect 1819 369 1857 403
rect 1891 369 1929 403
rect 1963 369 2001 403
rect 2035 369 2073 403
rect 2107 369 2145 403
rect 2179 369 2217 403
rect 2251 369 2289 403
rect 2323 369 2361 403
rect 2395 369 2433 403
rect 2467 369 2505 403
rect 2539 369 2577 403
rect 2611 369 2649 403
rect 2683 369 2721 403
rect 2755 369 2793 403
rect 2827 369 2865 403
rect 2899 369 2937 403
rect 2971 369 3009 403
rect 3043 369 3081 403
rect 3115 369 3153 403
rect 3187 369 3225 403
rect 3259 369 3297 403
rect 3331 369 3369 403
rect 3403 369 3441 403
rect 3475 369 3513 403
rect 3547 369 3585 403
rect 3619 369 3657 403
rect 3691 369 3729 403
rect 3763 369 3801 403
rect 3835 369 3873 403
rect 3907 369 3945 403
rect 3979 369 4017 403
rect 4051 369 4089 403
rect 4123 369 4161 403
rect 4195 369 4233 403
rect 4267 369 4305 403
rect 4339 369 4377 403
rect 4411 369 4449 403
rect 4483 369 4521 403
rect 4555 369 4593 403
rect 4627 369 4665 403
rect 4699 369 4737 403
rect 4771 369 4809 403
rect 4843 369 4881 403
rect 4915 369 4953 403
rect 4987 369 5025 403
rect 5059 369 5097 403
rect 5131 369 5169 403
rect 5203 369 5241 403
rect 5275 369 5313 403
rect 5347 369 5385 403
rect 5419 369 5457 403
rect 5491 369 5529 403
rect 5563 369 5601 403
rect 5635 369 5673 403
rect 5707 369 5745 403
rect 5779 369 5817 403
rect 5851 369 5889 403
rect 5923 369 5961 403
rect 5995 369 6033 403
rect 6067 369 6105 403
rect 6139 369 6177 403
rect 6211 369 9499 403
rect -53 363 9499 369
rect -53 289 9289 323
rect -53 143 119 243
rect 9327 143 9499 243
rect 166 63 9499 97
rect -53 17 9499 23
rect -53 -17 6309 17
rect 6343 -17 6381 17
rect 6415 -17 6453 17
rect 6487 -17 6525 17
rect 6559 -17 6597 17
rect 6631 -17 6669 17
rect 6703 -17 6741 17
rect 6775 -17 6813 17
rect 6847 -17 6885 17
rect 6919 -17 6957 17
rect 6991 -17 7029 17
rect 7063 -17 7101 17
rect 7135 -17 7173 17
rect 7207 -17 7245 17
rect 7279 -17 7317 17
rect 7351 -17 7389 17
rect 7423 -17 7461 17
rect 7495 -17 7533 17
rect 7567 -17 7605 17
rect 7639 -17 7677 17
rect 7711 -17 7749 17
rect 7783 -17 7821 17
rect 7855 -17 7893 17
rect 7927 -17 7965 17
rect 7999 -17 8037 17
rect 8071 -17 8109 17
rect 8143 -17 8181 17
rect 8215 -17 8253 17
rect 8287 -17 8325 17
rect 8359 -17 8397 17
rect 8431 -17 8469 17
rect 8503 -17 8541 17
rect 8575 -17 8613 17
rect 8647 -17 8685 17
rect 8719 -17 8757 17
rect 8791 -17 8829 17
rect 8863 -17 8901 17
rect 8935 -17 8973 17
rect 9007 -17 9045 17
rect 9079 -17 9117 17
rect 9151 -17 9189 17
rect 9223 -17 9261 17
rect 9295 -17 9333 17
rect 9367 -17 9405 17
rect 9439 -17 9499 17
rect -53 -53 9499 -17
use sky130_fd_pr__pfet_01v8_D9Q956  XM1
timestamp 1750100919
transform 0 1 3098 -1 0 193
box -246 -3151 246 3151
use sky130_fd_pr__nfet_01v8_H9ZN2D  XM2
timestamp 1750100919
transform 0 1 7874 -1 0 193
box -236 -1615 236 1615
<< labels >>
flabel metal1 s -32 391 -15 407 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s -33 -34 -16 -18 0 FreeSans 500 0 0 0 VSS
port 2 nsew
flabel metal1 s -43 300 -26 316 0 FreeSans 500 0 0 0 IN
port 3 nsew
flabel metal1 s -42 184 -25 200 0 FreeSans 500 0 0 0 SWP
port 4 nsew
flabel metal1 s 9472 178 9490 195 0 FreeSans 500 0 0 0 SWN
port 5 nsew
flabel metal1 s 9474 73 9492 90 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
