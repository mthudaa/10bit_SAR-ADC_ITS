magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect 142 1527 144 1561
rect 178 1527 216 1561
rect 250 1527 288 1561
rect 322 1527 360 1561
rect 394 1527 432 1561
rect 466 1527 504 1561
rect 538 1527 576 1561
rect 610 1527 648 1561
rect 682 1527 720 1561
rect 754 1527 792 1561
rect 826 1527 864 1561
rect 898 1527 936 1561
rect 970 1527 1008 1561
rect 1042 1527 1080 1561
rect 1114 1527 1152 1561
rect 1186 1527 1224 1561
rect 1258 1527 1296 1561
rect 1330 1527 1368 1561
rect 1402 1527 1440 1561
rect 1474 1527 1512 1561
rect 1546 1527 1584 1561
rect 1618 1527 1656 1561
rect 1690 1527 1728 1561
rect 1762 1527 1800 1561
rect 1834 1527 1872 1561
rect 1906 1527 1944 1561
rect 1978 1527 2016 1561
rect 2050 1527 2088 1561
rect 2122 1527 2160 1561
rect 2194 1527 2232 1561
rect 2266 1527 2304 1561
rect 2338 1527 2376 1561
rect 2410 1527 2448 1561
rect 2482 1527 2520 1561
rect 2554 1527 2592 1561
rect 2626 1527 2664 1561
rect 2698 1527 2736 1561
rect 2770 1527 2808 1561
rect 2842 1527 2880 1561
rect 2914 1527 2952 1561
rect 2986 1527 3024 1561
rect 3058 1527 3096 1561
rect 3130 1527 3168 1561
rect 3202 1527 3240 1561
rect 3274 1527 3312 1561
rect 3346 1527 3384 1561
rect 3418 1527 3456 1561
rect 3490 1527 3528 1561
rect 3562 1527 3600 1561
rect 3634 1527 3672 1561
rect 3706 1527 3744 1561
rect 3778 1527 3816 1561
rect 3850 1527 3888 1561
rect 3922 1527 3960 1561
rect 3994 1527 4032 1561
rect 4066 1527 4104 1561
rect 4138 1527 4176 1561
rect 4210 1527 4248 1561
rect 4282 1527 4320 1561
rect 4354 1527 4392 1561
rect 4426 1527 4464 1561
rect 4498 1527 4536 1561
rect 4570 1527 4608 1561
rect 4642 1527 4680 1561
rect 4714 1527 4752 1561
rect 4786 1527 4824 1561
rect 4858 1527 4896 1561
rect 4930 1527 4968 1561
rect 5002 1527 5040 1561
rect 5074 1527 5112 1561
rect 5146 1527 5184 1561
rect 5218 1527 5256 1561
rect 5290 1527 5328 1561
rect 5362 1527 5400 1561
rect 5434 1527 5472 1561
rect 5506 1527 5544 1561
rect 5578 1527 5616 1561
rect 5650 1527 5688 1561
rect 5722 1527 5760 1561
rect 5794 1527 5832 1561
rect 5866 1527 5904 1561
rect 5938 1527 5976 1561
rect 6010 1527 6048 1561
rect 6082 1527 6120 1561
rect 6154 1527 6192 1561
rect 6226 1527 6264 1561
rect 6298 1527 6336 1561
rect 6370 1527 6372 1561
rect 142 -123 166 -89
rect 200 -123 238 -89
rect 272 -123 310 -89
rect 344 -123 382 -89
rect 416 -123 454 -89
rect 488 -123 526 -89
rect 560 -123 598 -89
rect 632 -123 670 -89
rect 704 -123 742 -89
rect 776 -123 814 -89
rect 848 -123 886 -89
rect 920 -123 958 -89
rect 992 -123 1030 -89
rect 1064 -123 1102 -89
rect 1136 -123 1174 -89
rect 1208 -123 1246 -89
rect 1280 -123 1318 -89
rect 1352 -123 1390 -89
rect 1424 -123 1462 -89
rect 1496 -123 1534 -89
rect 1568 -123 1606 -89
rect 1640 -123 1678 -89
rect 1712 -123 1750 -89
rect 1784 -123 1822 -89
rect 1856 -123 1894 -89
rect 1928 -123 1966 -89
rect 2000 -123 2038 -89
rect 2072 -123 2110 -89
rect 2144 -123 2182 -89
rect 2216 -123 2254 -89
rect 2288 -123 2326 -89
rect 2360 -123 2398 -89
rect 2432 -123 2470 -89
rect 2504 -123 2542 -89
rect 2576 -123 2614 -89
rect 2648 -123 2686 -89
rect 2720 -123 2758 -89
rect 2792 -123 2830 -89
rect 2864 -123 2902 -89
rect 2936 -123 2974 -89
rect 3008 -123 3046 -89
rect 3080 -123 3118 -89
rect 3152 -123 3190 -89
rect 3224 -123 3262 -89
rect 3296 -123 3320 -89
<< viali >>
rect 144 1527 178 1561
rect 216 1527 250 1561
rect 288 1527 322 1561
rect 360 1527 394 1561
rect 432 1527 466 1561
rect 504 1527 538 1561
rect 576 1527 610 1561
rect 648 1527 682 1561
rect 720 1527 754 1561
rect 792 1527 826 1561
rect 864 1527 898 1561
rect 936 1527 970 1561
rect 1008 1527 1042 1561
rect 1080 1527 1114 1561
rect 1152 1527 1186 1561
rect 1224 1527 1258 1561
rect 1296 1527 1330 1561
rect 1368 1527 1402 1561
rect 1440 1527 1474 1561
rect 1512 1527 1546 1561
rect 1584 1527 1618 1561
rect 1656 1527 1690 1561
rect 1728 1527 1762 1561
rect 1800 1527 1834 1561
rect 1872 1527 1906 1561
rect 1944 1527 1978 1561
rect 2016 1527 2050 1561
rect 2088 1527 2122 1561
rect 2160 1527 2194 1561
rect 2232 1527 2266 1561
rect 2304 1527 2338 1561
rect 2376 1527 2410 1561
rect 2448 1527 2482 1561
rect 2520 1527 2554 1561
rect 2592 1527 2626 1561
rect 2664 1527 2698 1561
rect 2736 1527 2770 1561
rect 2808 1527 2842 1561
rect 2880 1527 2914 1561
rect 2952 1527 2986 1561
rect 3024 1527 3058 1561
rect 3096 1527 3130 1561
rect 3168 1527 3202 1561
rect 3240 1527 3274 1561
rect 3312 1527 3346 1561
rect 3384 1527 3418 1561
rect 3456 1527 3490 1561
rect 3528 1527 3562 1561
rect 3600 1527 3634 1561
rect 3672 1527 3706 1561
rect 3744 1527 3778 1561
rect 3816 1527 3850 1561
rect 3888 1527 3922 1561
rect 3960 1527 3994 1561
rect 4032 1527 4066 1561
rect 4104 1527 4138 1561
rect 4176 1527 4210 1561
rect 4248 1527 4282 1561
rect 4320 1527 4354 1561
rect 4392 1527 4426 1561
rect 4464 1527 4498 1561
rect 4536 1527 4570 1561
rect 4608 1527 4642 1561
rect 4680 1527 4714 1561
rect 4752 1527 4786 1561
rect 4824 1527 4858 1561
rect 4896 1527 4930 1561
rect 4968 1527 5002 1561
rect 5040 1527 5074 1561
rect 5112 1527 5146 1561
rect 5184 1527 5218 1561
rect 5256 1527 5290 1561
rect 5328 1527 5362 1561
rect 5400 1527 5434 1561
rect 5472 1527 5506 1561
rect 5544 1527 5578 1561
rect 5616 1527 5650 1561
rect 5688 1527 5722 1561
rect 5760 1527 5794 1561
rect 5832 1527 5866 1561
rect 5904 1527 5938 1561
rect 5976 1527 6010 1561
rect 6048 1527 6082 1561
rect 6120 1527 6154 1561
rect 6192 1527 6226 1561
rect 6264 1527 6298 1561
rect 6336 1527 6370 1561
rect 166 -123 200 -89
rect 238 -123 272 -89
rect 310 -123 344 -89
rect 382 -123 416 -89
rect 454 -123 488 -89
rect 526 -123 560 -89
rect 598 -123 632 -89
rect 670 -123 704 -89
rect 742 -123 776 -89
rect 814 -123 848 -89
rect 886 -123 920 -89
rect 958 -123 992 -89
rect 1030 -123 1064 -89
rect 1102 -123 1136 -89
rect 1174 -123 1208 -89
rect 1246 -123 1280 -89
rect 1318 -123 1352 -89
rect 1390 -123 1424 -89
rect 1462 -123 1496 -89
rect 1534 -123 1568 -89
rect 1606 -123 1640 -89
rect 1678 -123 1712 -89
rect 1750 -123 1784 -89
rect 1822 -123 1856 -89
rect 1894 -123 1928 -89
rect 1966 -123 2000 -89
rect 2038 -123 2072 -89
rect 2110 -123 2144 -89
rect 2182 -123 2216 -89
rect 2254 -123 2288 -89
rect 2326 -123 2360 -89
rect 2398 -123 2432 -89
rect 2470 -123 2504 -89
rect 2542 -123 2576 -89
rect 2614 -123 2648 -89
rect 2686 -123 2720 -89
rect 2758 -123 2792 -89
rect 2830 -123 2864 -89
rect 2902 -123 2936 -89
rect 2974 -123 3008 -89
rect 3046 -123 3080 -89
rect 3118 -123 3152 -89
rect 3190 -123 3224 -89
rect 3262 -123 3296 -89
<< metal1 >>
rect 106 1561 6408 1597
rect 106 1527 144 1561
rect 178 1527 216 1561
rect 250 1527 288 1561
rect 322 1527 360 1561
rect 394 1527 432 1561
rect 466 1527 504 1561
rect 538 1527 576 1561
rect 610 1527 648 1561
rect 682 1527 720 1561
rect 754 1527 792 1561
rect 826 1527 864 1561
rect 898 1527 936 1561
rect 970 1527 1008 1561
rect 1042 1527 1080 1561
rect 1114 1527 1152 1561
rect 1186 1527 1224 1561
rect 1258 1527 1296 1561
rect 1330 1527 1368 1561
rect 1402 1527 1440 1561
rect 1474 1527 1512 1561
rect 1546 1527 1584 1561
rect 1618 1527 1656 1561
rect 1690 1527 1728 1561
rect 1762 1527 1800 1561
rect 1834 1527 1872 1561
rect 1906 1527 1944 1561
rect 1978 1527 2016 1561
rect 2050 1527 2088 1561
rect 2122 1527 2160 1561
rect 2194 1527 2232 1561
rect 2266 1527 2304 1561
rect 2338 1527 2376 1561
rect 2410 1527 2448 1561
rect 2482 1527 2520 1561
rect 2554 1527 2592 1561
rect 2626 1527 2664 1561
rect 2698 1527 2736 1561
rect 2770 1527 2808 1561
rect 2842 1527 2880 1561
rect 2914 1527 2952 1561
rect 2986 1527 3024 1561
rect 3058 1527 3096 1561
rect 3130 1527 3168 1561
rect 3202 1527 3240 1561
rect 3274 1527 3312 1561
rect 3346 1527 3384 1561
rect 3418 1527 3456 1561
rect 3490 1527 3528 1561
rect 3562 1527 3600 1561
rect 3634 1527 3672 1561
rect 3706 1527 3744 1561
rect 3778 1527 3816 1561
rect 3850 1527 3888 1561
rect 3922 1527 3960 1561
rect 3994 1527 4032 1561
rect 4066 1527 4104 1561
rect 4138 1527 4176 1561
rect 4210 1527 4248 1561
rect 4282 1527 4320 1561
rect 4354 1527 4392 1561
rect 4426 1527 4464 1561
rect 4498 1527 4536 1561
rect 4570 1527 4608 1561
rect 4642 1527 4680 1561
rect 4714 1527 4752 1561
rect 4786 1527 4824 1561
rect 4858 1527 4896 1561
rect 4930 1527 4968 1561
rect 5002 1527 5040 1561
rect 5074 1527 5112 1561
rect 5146 1527 5184 1561
rect 5218 1527 5256 1561
rect 5290 1527 5328 1561
rect 5362 1527 5400 1561
rect 5434 1527 5472 1561
rect 5506 1527 5544 1561
rect 5578 1527 5616 1561
rect 5650 1527 5688 1561
rect 5722 1527 5760 1561
rect 5794 1527 5832 1561
rect 5866 1527 5904 1561
rect 5938 1527 5976 1561
rect 6010 1527 6048 1561
rect 6082 1527 6120 1561
rect 6154 1527 6192 1561
rect 6226 1527 6264 1561
rect 6298 1527 6336 1561
rect 6370 1527 6408 1561
rect 106 1521 6408 1527
rect 325 1447 6189 1521
rect 106 1377 284 1401
rect 106 1325 176 1377
rect 228 1325 284 1377
rect 106 1301 284 1325
rect 325 1061 6189 1255
rect 106 915 284 1015
rect 106 569 6408 869
rect 106 423 284 523
rect 316 183 3146 377
rect 166 113 284 137
rect 166 61 176 113
rect 228 61 284 113
rect 166 37 284 61
rect 316 -83 3146 -9
rect 106 -89 6408 -83
rect 106 -123 166 -89
rect 200 -123 238 -89
rect 272 -123 310 -89
rect 344 -123 382 -89
rect 416 -123 454 -89
rect 488 -123 526 -89
rect 560 -123 598 -89
rect 632 -123 670 -89
rect 704 -123 742 -89
rect 776 -123 814 -89
rect 848 -123 886 -89
rect 920 -123 958 -89
rect 992 -123 1030 -89
rect 1064 -123 1102 -89
rect 1136 -123 1174 -89
rect 1208 -123 1246 -89
rect 1280 -123 1318 -89
rect 1352 -123 1390 -89
rect 1424 -123 1462 -89
rect 1496 -123 1534 -89
rect 1568 -123 1606 -89
rect 1640 -123 1678 -89
rect 1712 -123 1750 -89
rect 1784 -123 1822 -89
rect 1856 -123 1894 -89
rect 1928 -123 1966 -89
rect 2000 -123 2038 -89
rect 2072 -123 2110 -89
rect 2144 -123 2182 -89
rect 2216 -123 2254 -89
rect 2288 -123 2326 -89
rect 2360 -123 2398 -89
rect 2432 -123 2470 -89
rect 2504 -123 2542 -89
rect 2576 -123 2614 -89
rect 2648 -123 2686 -89
rect 2720 -123 2758 -89
rect 2792 -123 2830 -89
rect 2864 -123 2902 -89
rect 2936 -123 2974 -89
rect 3008 -123 3046 -89
rect 3080 -123 3118 -89
rect 3152 -123 3190 -89
rect 3224 -123 3262 -89
rect 3296 -123 6408 -89
rect 106 -159 6408 -123
<< via1 >>
rect 176 1325 228 1377
rect 176 61 228 113
<< metal2 >>
rect 176 1377 228 1411
rect 176 113 228 1325
rect 176 27 228 61
use sky130_fd_pr__nfet_01v8_H9ZN2D  sky130_fd_pr__nfet_01v8_H9ZN2D_0
timestamp 1750100919
transform 0 1 1731 -1 0 87
box -236 -1615 236 1615
use sky130_fd_pr__pfet_01v8_D9Q956  sky130_fd_pr__pfet_01v8_D9Q956_0
timestamp 1750100919
transform 0 1 3257 -1 0 965
box -246 -3151 246 3151
use sky130_fd_pr__pfet_01v8_D9Q956  XM1
timestamp 1750100919
transform 0 1 3257 -1 0 1351
box -246 -3151 246 3151
use sky130_fd_pr__nfet_01v8_H9ZN2D  XM3
timestamp 1750100919
transform 0 1 1731 -1 0 473
box -236 -1615 236 1615
<< labels >>
flabel metal1 s 113 1556 120 1563 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 119 1345 126 1352 0 FreeSans 500 0 0 0 IN
port 2 nsew
flabel metal1 s 119 960 126 967 0 FreeSans 500 0 0 0 CKB
port 3 nsew
flabel metal1 s 119 469 126 476 0 FreeSans 500 0 0 0 CK
port 4 nsew
flabel metal1 s 122 -125 129 -118 0 FreeSans 500 0 0 0 VSS
port 5 nsew
flabel metal1 s 6347 690 6354 697 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
