magic
tech sky130A
magscale 1 2
timestamp 1749657747
<< dnwell >>
rect -10590 64857 -3793 76025
rect -7487 55533 -3793 64857
rect -10580 44365 -3783 55533
rect -2373 1624 49198 118766
rect 50479 58365 56127 62017
rect 59127 45909 70849 74783
<< metal1 >>
rect -11103 121841 61079 122097
rect 61479 121841 67079 122097
rect 67479 121841 71105 122097
rect -11103 121329 -10580 121585
rect -10484 121329 -3901 121585
rect -3803 121329 50489 121585
rect 50585 121329 56021 121585
rect 56117 121329 71105 121585
rect -11103 120816 46777 121072
rect 46917 120816 71105 121072
rect -2083 115221 -1943 120816
rect -1333 120461 70091 120561
rect 70147 120461 70157 120561
rect -1333 118607 -1233 120461
rect 3469 120261 68939 120361
rect 68995 120261 69005 120361
rect 3469 118690 3569 120261
rect 8271 120061 67787 120161
rect 67843 120061 67853 120161
rect 8271 118659 8371 120061
rect 13073 119861 66635 119961
rect 66691 119861 66701 119961
rect 13073 118671 13173 119861
rect 17875 119661 65483 119761
rect 65539 119661 65549 119761
rect 17875 118665 17975 119661
rect 22677 119461 64331 119561
rect 64387 119461 64397 119561
rect 22677 118632 22777 119461
rect 27479 119261 63179 119361
rect 63235 119261 63245 119361
rect 27479 118674 27579 119261
rect 32281 119061 62027 119161
rect 62083 119061 62093 119161
rect 32281 118632 32381 119061
rect 37083 118861 60875 118961
rect 60931 118861 60941 118961
rect 37083 118613 37183 118861
rect 41885 118661 59723 118761
rect 59779 118661 59789 118761
rect -2093 115081 -2083 115221
rect -1943 115081 -1933 115221
rect -10590 76025 -10580 76121
rect -10484 76025 -10474 76121
rect -4251 67457 -4241 67509
rect -4189 67457 -4179 67509
rect -10581 61051 -10325 63867
rect 614 61819 624 61900
rect -4692 61563 624 61819
rect 44492 61563 49994 61900
rect 50046 61563 50056 61900
rect -3739 61371 -3729 61435
rect -3665 61371 49261 61435
rect 49325 61371 49335 61435
rect -4576 60582 -4566 60678
rect -4470 60582 50681 60678
rect 50777 60582 50787 60678
rect 50367 60347 50377 60399
rect 50429 60390 50439 60399
rect 50429 60356 50623 60390
rect 50429 60347 50439 60356
rect 49984 60282 49994 60334
rect 50046 60316 50056 60334
rect 50046 60282 50737 60316
rect 49984 60048 49994 60100
rect 50046 60066 50538 60100
rect 50046 60048 50056 60066
rect 55955 59899 58407 59939
rect 58397 59887 58407 59899
rect 58527 59887 58537 59939
rect -3911 59778 -3901 59874
rect -3805 59778 50489 59874
rect 50585 59778 50595 59874
rect 58637 59727 58647 59779
rect 58767 59727 58777 59779
rect 55964 59687 58777 59727
rect 55930 59608 58777 59648
rect 58637 59556 58647 59608
rect 58767 59556 58777 59608
rect -10581 56523 -10325 59339
rect -3739 58955 -3729 59019
rect -3665 58955 49262 59019
rect 49326 58955 49336 59019
rect -4704 58571 624 58827
rect 614 58490 624 58571
rect 44492 58490 49994 58827
rect 50046 58490 50056 58827
rect -4251 52881 -4241 52933
rect -4189 52881 -4179 52933
rect -4576 44269 -4566 44365
rect -4470 44269 -4460 44365
rect -10590 43955 -3336 44075
rect -3216 43955 -3206 44075
rect -10590 43715 -2362 43835
rect -2222 43715 -2212 43835
rect -10590 43475 -3469 43595
rect -3349 43475 -3339 43595
rect -1813 5369 -1803 5509
rect -1663 5369 -1653 5509
rect -1803 -432 -1663 5369
rect -1332 -76 -1232 1737
rect 3470 124 3570 1737
rect 8272 324 8372 1698
rect 13074 524 13174 1688
rect 17876 724 17976 1748
rect 22678 924 22778 1743
rect 27480 1124 27580 1798
rect 32282 1324 32382 1700
rect 37084 1524 37184 1680
rect 41886 1624 59723 1724
rect 59779 1624 59789 1724
rect 37084 1424 60875 1524
rect 60931 1424 60941 1524
rect 32282 1224 62027 1324
rect 62083 1224 62093 1324
rect 27480 1024 63179 1124
rect 63235 1024 63245 1124
rect 22678 824 64331 924
rect 64387 824 64397 924
rect 17876 624 65483 724
rect 65539 624 65549 724
rect 13074 424 66635 524
rect 66691 424 66701 524
rect 8272 224 67787 324
rect 67843 224 67853 324
rect 3470 24 68939 124
rect 68995 24 69005 124
rect -1332 -176 70091 -76
rect 70147 -176 70157 -76
rect -11102 -688 46497 -432
rect 46638 -688 71106 -432
rect -11102 -1200 -4566 -944
rect -4470 -1200 50681 -944
rect 50777 -1200 55829 -944
rect 55925 -1200 71106 -944
rect -11102 -1713 64079 -1457
rect 64479 -1713 71106 -1457
<< via1 >>
rect 61079 121841 61479 122097
rect 67079 121841 67479 122097
rect -10580 121329 -10484 121585
rect -3901 121329 -3803 121585
rect 50489 121329 50585 121585
rect 56021 121329 56117 121585
rect 46777 120816 46917 121072
rect 70091 120461 70147 120561
rect 68939 120261 68995 120361
rect 67787 120061 67843 120161
rect 66635 119861 66691 119961
rect 65483 119661 65539 119761
rect 64331 119461 64387 119561
rect 63179 119261 63235 119361
rect 62027 119061 62083 119161
rect 60875 118861 60931 118961
rect 59723 118661 59779 118761
rect -2083 115081 -1943 115221
rect -10580 76025 -10484 76121
rect -4241 67457 -4189 67509
rect 624 61563 44492 61900
rect 49994 61563 50046 61900
rect -3729 61371 -3665 61435
rect 49261 61371 49325 61435
rect -4566 60582 -4470 60678
rect 50681 60582 50777 60678
rect 50377 60347 50429 60399
rect 49994 60282 50046 60334
rect 49994 60048 50046 60100
rect 58407 59887 58527 59939
rect -3901 59778 -3805 59874
rect 50489 59778 50585 59874
rect 58647 59727 58767 59779
rect 58647 59556 58767 59608
rect -3729 58955 -3665 59019
rect 49262 58955 49326 59019
rect 624 58490 44492 58827
rect 49994 58490 50046 58827
rect -4241 52881 -4189 52933
rect -4566 44269 -4470 44365
rect -3336 43955 -3216 44075
rect -2362 43715 -2222 43835
rect -3469 43475 -3349 43595
rect -1803 5369 -1663 5509
rect 59723 1624 59779 1724
rect 60875 1424 60931 1524
rect 62027 1224 62083 1324
rect 63179 1024 63235 1124
rect 64331 824 64387 924
rect 65483 624 65539 724
rect 66635 424 66691 524
rect 67787 224 67843 324
rect 68939 24 68995 124
rect 70091 -176 70147 -76
rect 46497 -688 46638 -432
rect -4566 -1200 -4470 -944
rect 50681 -1200 50777 -944
rect 55829 -1200 55925 -944
rect 64079 -1713 64479 -1457
<< metal2 >>
rect 61079 122097 61479 122107
rect 61079 121831 61479 121841
rect 67079 122097 67479 122107
rect 67079 121831 67479 121841
rect -10580 121585 -10484 121595
rect -10580 76121 -10484 121329
rect -3901 121585 -3803 121595
rect -3901 121319 -3803 121329
rect 50489 121585 50585 121595
rect 46777 121072 46917 121082
rect 46777 120806 46917 120816
rect -2083 115221 -1943 115231
rect -2083 115071 -1943 115081
rect 46777 115221 46917 115231
rect 46777 115071 46917 115081
rect -10580 76015 -10484 76025
rect 49261 72091 49325 72101
rect 49097 69131 49217 69141
rect 49097 69001 49217 69011
rect 48897 67651 49017 67661
rect -4241 67509 -4189 67519
rect -3729 67515 -3665 67525
rect 48897 67521 49017 67531
rect -4189 67457 -3729 67509
rect -4241 67447 -4189 67457
rect -3665 67457 -3621 67509
rect -3729 67441 -3665 67451
rect 48697 66171 48817 66181
rect 48697 66041 48817 66051
rect 48497 64691 48617 64701
rect 48497 64561 48617 64571
rect 48297 63211 48417 63221
rect 48297 63081 48417 63091
rect 48097 62611 48217 62621
rect 48097 62481 48217 62491
rect 624 61900 44492 61910
rect 624 61553 44492 61563
rect -3729 61435 -3665 61445
rect -3729 61361 -3665 61371
rect 49261 61435 49325 71971
rect 49261 61361 49325 61371
rect 49994 61900 50046 61910
rect 50489 61753 50585 121329
rect 56021 121585 56117 121595
rect 56021 61765 56117 121329
rect 70091 120561 70147 120571
rect 68939 120361 68995 120371
rect 67787 120161 67843 120171
rect 66635 119961 66691 119971
rect 65483 119761 65539 119771
rect 64331 119561 64387 119571
rect 63179 119361 63235 119371
rect 62027 119161 62083 119171
rect 60875 118961 60931 118971
rect 59723 118761 59779 118771
rect 59723 74724 59779 118661
rect 60875 74579 60931 118861
rect 62027 74727 62083 119061
rect 63179 74697 63235 119261
rect 64331 74694 64387 119461
rect 65483 74727 65539 119661
rect 66635 74707 66691 119861
rect 67787 74718 67843 120061
rect 68939 74701 68995 120261
rect 70091 74726 70147 120461
rect 58647 70611 58767 70621
rect -4566 60678 -4470 60688
rect -4566 60572 -4470 60582
rect 49994 60334 50046 61563
rect 50681 60678 50777 60688
rect 50681 60572 50777 60582
rect 49994 60272 50046 60282
rect 50377 60399 50429 60409
rect 50377 60234 50429 60347
rect -3280 60224 -3216 60234
rect -3901 59874 -3805 59884
rect -3901 59768 -3805 59778
rect -3729 59019 -3665 59029
rect -3729 58945 -3665 58955
rect -4241 52933 -4189 52943
rect -3729 52939 -3665 52949
rect -4189 52881 -3729 52933
rect -4241 52871 -4189 52881
rect -3729 52865 -3665 52875
rect -4566 44365 -4470 44375
rect -4566 -944 -4470 44269
rect -3280 44085 -3216 60160
rect 50365 60224 50429 60234
rect 50365 60150 50429 60160
rect 49994 60100 50046 60110
rect 49262 59019 49326 59029
rect 624 58827 44492 58837
rect 624 58480 44492 58490
rect 47898 58251 48018 58261
rect 47898 58121 48018 58131
rect 47698 57891 47818 57901
rect 47698 57761 47818 57771
rect 47498 57291 47618 57301
rect 47498 57161 47618 57171
rect 47298 55811 47418 55821
rect 47298 55681 47418 55691
rect 49262 48411 49326 58955
rect 49994 58827 50046 60048
rect 49994 58480 50046 58490
rect 50377 51381 50429 60150
rect 58407 59939 58527 59949
rect 50489 59874 50585 59884
rect 50489 59768 50585 59778
rect 50375 51371 50431 51381
rect 50375 51241 50431 51251
rect 49262 48281 49326 48291
rect 49686 49891 49806 49901
rect -3336 44075 -3216 44085
rect -3336 43945 -3216 43955
rect -2362 43835 -2222 43845
rect -2362 43705 -2222 43715
rect -3469 43595 -3349 43605
rect -3469 43465 -3349 43475
rect -1803 5509 -1663 5519
rect -1803 5359 -1663 5369
rect 46497 5510 46638 5520
rect 46497 5359 46638 5369
rect -3469 -240 -3349 -230
rect 49686 -240 49806 49771
rect -3349 -360 49806 -240
rect -3469 -370 -3349 -360
rect 46497 -432 46638 -422
rect 46497 -698 46638 -688
rect -4566 -1210 -4470 -1200
rect 50681 -944 50777 59494
rect 50681 -1210 50777 -1200
rect 55829 -944 55925 58910
rect 58407 52851 58527 59887
rect 58647 59779 58767 70491
rect 59127 62611 59247 62621
rect 59127 61731 59247 62491
rect 59127 61601 59247 61611
rect 58647 59687 58767 59727
rect 58887 60251 59007 60261
rect 58647 59608 58767 59648
rect 58647 54331 58767 59556
rect 58887 58251 59007 60131
rect 58887 58121 59007 58131
rect 59127 58771 59247 58781
rect 59127 57891 59247 58651
rect 59127 57761 59247 57771
rect 58647 54201 58767 54211
rect 58407 52721 58527 52731
rect 59723 1724 59779 46402
rect 59723 1614 59779 1624
rect 60875 1524 60931 46402
rect 60875 1414 60931 1424
rect 62027 1324 62083 46402
rect 62027 1214 62083 1224
rect 63179 1124 63235 46402
rect 63179 1014 63235 1024
rect 64331 924 64387 46402
rect 64331 814 64387 824
rect 65483 724 65539 46402
rect 65483 614 65539 624
rect 66635 524 66691 46402
rect 66635 414 66691 424
rect 67787 324 67843 46402
rect 67787 214 67843 224
rect 68939 124 68995 46402
rect 68939 14 68995 24
rect 70091 -76 70147 46402
rect 70091 -186 70147 -176
rect 55829 -1210 55925 -1200
rect 64079 -1457 64479 -1447
rect 64079 -1723 64479 -1713
<< via2 >>
rect 61079 121841 61479 122097
rect 67079 121841 67479 122097
rect -3901 121329 -3803 121585
rect 46777 120816 46917 121072
rect 46777 115081 46917 115221
rect 49261 71971 49325 72091
rect 49097 69011 49217 69131
rect 48897 67531 49017 67651
rect -3729 67451 -3665 67515
rect 48697 66051 48817 66171
rect 48497 64571 48617 64691
rect 48297 63091 48417 63211
rect 48097 62491 48217 62611
rect 624 61563 44492 61900
rect -3729 61371 -3665 61435
rect 58647 70491 58767 70611
rect -4566 60582 -4470 60678
rect -3280 60160 -3216 60224
rect -3901 59778 -3805 59874
rect -3729 58955 -3665 59019
rect -3729 52875 -3665 52939
rect 50365 60160 50429 60224
rect 624 58490 44492 58827
rect 47898 58131 48018 58251
rect 47698 57771 47818 57891
rect 47498 57171 47618 57291
rect 47298 55691 47418 55811
rect 50375 51251 50431 51371
rect 49262 48291 49326 48411
rect 49686 49771 49806 49891
rect -3469 43475 -3349 43595
rect 46497 5369 46638 5510
rect -3469 -360 -3349 -240
rect 46497 -688 46638 -432
rect 59127 62491 59247 62611
rect 59127 61611 59247 61731
rect 58887 60131 59007 60251
rect 58887 58131 59007 58251
rect 59127 58651 59247 58771
rect 59127 57771 59247 57891
rect 58647 54211 58767 54331
rect 58407 52731 58527 52851
rect 64079 -1713 64479 -1457
<< metal3 >>
rect 61069 122097 61489 122102
rect 61069 121841 61079 122097
rect 61479 121841 61489 122097
rect 61069 121836 61489 121841
rect 67069 122097 67489 122102
rect 67069 121841 67079 122097
rect 67479 121841 67489 122097
rect 67069 121836 67489 121841
rect -3911 121585 -3793 121590
rect -3911 121329 -3901 121585
rect -3803 121329 -3793 121585
rect -3911 121324 -3793 121329
rect -3901 64788 -3803 121324
rect 46767 121072 46927 121077
rect 46767 120816 46777 121072
rect 46917 120816 46927 121072
rect 46767 120811 46927 120816
rect 46777 115226 46917 120811
rect 46767 115221 46927 115226
rect 46767 115081 46777 115221
rect 46917 115081 46927 115221
rect 46767 115076 46927 115081
rect 70049 73155 70849 73275
rect 49251 72091 49335 72096
rect 49251 71971 49261 72091
rect 49325 71971 59263 72091
rect 49251 71966 49335 71971
rect 58637 70611 58777 70616
rect 58637 70491 58647 70611
rect 58767 70491 59127 70611
rect 58637 70486 58777 70491
rect 49087 69131 49227 69136
rect 49087 69011 49097 69131
rect 49217 69011 59247 69131
rect 49087 69006 49227 69011
rect 70049 68419 70849 68539
rect 48887 67651 49027 67656
rect 48887 67531 48897 67651
rect 49017 67531 59267 67651
rect 48887 67526 49027 67531
rect -3739 67515 -3655 67520
rect -3739 67451 -3729 67515
rect -3665 67451 -3655 67515
rect -3739 67446 -3655 67451
rect -3729 61440 -3665 67446
rect 48687 66171 48827 66176
rect 48687 66051 48697 66171
rect 48817 66051 59247 66171
rect 70049 66051 70849 66171
rect 48687 66046 48827 66051
rect 48487 64691 48627 64696
rect 48487 64571 48497 64691
rect 48617 64571 59247 64691
rect 48487 64566 48627 64571
rect 70049 63683 70849 63803
rect 48287 63211 48427 63216
rect 48287 63091 48297 63211
rect 48417 63091 59247 63211
rect 48287 63086 48427 63091
rect 48087 62611 48227 62616
rect 59117 62611 59257 62616
rect 48087 62491 48097 62611
rect 48217 62491 59127 62611
rect 59247 62491 59257 62611
rect 48087 62486 48227 62491
rect 59117 62486 59257 62491
rect 614 61900 44502 61905
rect 614 61563 624 61900
rect 44492 61563 44502 61900
rect 59117 61731 59257 61736
rect 59117 61611 59127 61731
rect 59247 61611 59257 61731
rect 59117 61606 59257 61611
rect 614 61558 44502 61563
rect -3739 61435 -3655 61440
rect -3739 61371 -3729 61435
rect -3665 61371 -3655 61435
rect -3739 61366 -3655 61371
rect 70049 61315 70849 61435
rect -4576 60678 -4460 60683
rect -4576 60582 -4566 60678
rect -4470 60582 -4460 60678
rect -4576 60577 -4460 60582
rect 58877 60251 59017 60256
rect -3290 60224 -3206 60229
rect 50355 60224 50439 60229
rect -3290 60160 -3280 60224
rect -3216 60160 50365 60224
rect 50429 60160 50439 60224
rect -3290 60155 -3206 60160
rect 50355 60155 50439 60160
rect 58877 60131 58887 60251
rect 59007 60131 59127 60251
rect 58877 60126 59017 60131
rect -3911 59874 -3795 59879
rect -3911 59778 -3901 59874
rect -3805 59778 -3795 59874
rect -3911 59773 -3795 59778
rect -3739 59019 -3655 59024
rect -3739 58955 -3729 59019
rect -3665 58955 -3655 59019
rect -3739 58950 -3655 58955
rect -3729 52944 -3665 58950
rect 70049 58947 70849 59067
rect 614 58827 44502 58832
rect 614 58490 624 58827
rect 44492 58490 44502 58827
rect 59117 58771 59257 58776
rect 59117 58651 59127 58771
rect 59247 58651 59257 58771
rect 59117 58646 59257 58651
rect 614 58485 44502 58490
rect 47888 58251 48028 58256
rect 58877 58251 59017 58256
rect 47888 58131 47898 58251
rect 48018 58131 58887 58251
rect 59007 58131 59017 58251
rect 47888 58126 48028 58131
rect 58877 58126 59017 58131
rect 47688 57891 47828 57896
rect 59117 57891 59257 57896
rect 47688 57771 47698 57891
rect 47818 57771 59127 57891
rect 59247 57771 59257 57891
rect 47688 57766 47828 57771
rect 59117 57766 59257 57771
rect 47488 57291 47628 57296
rect 47488 57171 47498 57291
rect 47618 57171 59247 57291
rect 47488 57166 47628 57171
rect 70049 56579 70849 56699
rect 47288 55811 47428 55816
rect 47288 55691 47298 55811
rect 47418 55691 59248 55811
rect 47288 55686 47428 55691
rect 58637 54331 58777 54336
rect 58637 54211 58647 54331
rect 58767 54211 59127 54331
rect 70049 54211 70849 54331
rect 58637 54206 58777 54211
rect -3739 52939 -3655 52944
rect -3739 52875 -3729 52939
rect -3665 52875 -3655 52939
rect -3739 52870 -3655 52875
rect 58397 52851 58537 52856
rect 58397 52731 58407 52851
rect 58527 52731 59127 52851
rect 58397 52726 58537 52731
rect 70049 51843 70849 51963
rect 50365 51371 50441 51376
rect 50365 51251 50375 51371
rect 50431 51251 59288 51371
rect 50365 51246 50441 51251
rect 49676 49891 49816 49896
rect 49676 49771 49686 49891
rect 49806 49771 59279 49891
rect 49676 49766 49816 49771
rect 70049 49475 70849 49595
rect 49252 48411 49336 48416
rect 49252 48291 49262 48411
rect 49326 48291 59391 48411
rect 49252 48286 49336 48291
rect 70049 47107 70849 47227
rect -3479 43595 -3339 43600
rect -3479 43475 -3469 43595
rect -3349 43475 -3339 43595
rect -3479 43470 -3339 43475
rect -3469 -235 -3349 43470
rect 46487 5510 46648 5515
rect 46487 5369 46497 5510
rect 46638 5369 46648 5510
rect 46487 5364 46648 5369
rect -3479 -240 -3339 -235
rect -3479 -360 -3469 -240
rect -3349 -360 -3339 -240
rect -3479 -365 -3339 -360
rect 46497 -427 46638 5364
rect 46487 -432 46648 -427
rect 46487 -688 46497 -432
rect 46638 -688 46648 -432
rect 46487 -693 46648 -688
rect 64069 -1457 64489 -1452
rect 64069 -1713 64079 -1457
rect 64479 -1713 64489 -1457
rect 64069 -1718 64489 -1713
<< via3 >>
rect 61079 121841 61479 122097
rect 67079 121841 67479 122097
rect 624 61563 44492 61900
rect 624 58490 44492 58827
rect 64079 -1713 64479 -1457
<< metal4 >>
rect 61078 122097 61480 122098
rect 61078 121841 61079 122097
rect 61479 121841 61480 122097
rect 61078 121840 61480 121841
rect 67078 122097 67480 122098
rect 67078 121841 67079 122097
rect 67479 121841 67480 122097
rect 67078 121840 67480 121841
rect 61079 71451 61479 121840
rect 67079 71328 67479 121840
rect 623 61900 44493 61901
rect 623 61563 624 61900
rect 44492 61563 44493 61900
rect 623 61562 44493 61563
rect 623 58827 44493 58828
rect 623 58490 624 58827
rect 44492 58490 44493 58827
rect 623 58489 44493 58490
rect 64079 -1456 64479 49005
rect 64078 -1457 64480 -1456
rect 64078 -1713 64079 -1457
rect 64479 -1713 64480 -1457
rect 64078 -1714 64480 -1713
use cdac  cdac_0
timestamp 1749497408
transform 1 0 -1274 0 1 2329
box -1099 -705 50472 116437
use sar10b  sar10b_0
timestamp 1749574357
transform 1 0 59127 0 1 45909
box 0 0 11722 28874
use tdc  tdc_0
timestamp 1749411235
transform 1 0 50703 0 1 59011
box -224 -646 5424 3006
use th_dif_sw  th_dif_sw_0
timestamp 1749656470
transform 0 -1 -4206 1 0 44365
box -1 -413 31660 6384
<< labels >>
flabel metal1 -10590 43715 -10470 43835 0 FreeSans 800 0 0 0 VCM
port 0 nsew
flabel metal1 -10590 43475 -10470 43595 0 FreeSans 800 0 0 0 EN
port 1 nsew
flabel metal1 -11103 121329 -10847 121585 0 FreeSans 800 0 0 0 VDDA
port 3 nsew
flabel metal1 -11103 120816 -10847 121072 0 FreeSans 800 0 0 0 VDDR
port 4 nsew
flabel metal1 -10590 43955 -10470 44075 0 FreeSans 800 0 0 0 CLK
port 10 nsew
flabel metal3 70729 73155 70849 73275 0 FreeSans 800 0 0 0 CKO
port 11 nsew
flabel metal3 70729 66051 70849 66171 0 FreeSans 800 0 0 0 DATA[8]
port 13 nsew
flabel metal3 70729 63683 70849 63803 0 FreeSans 800 0 0 0 DATA[7]
port 14 nsew
flabel metal3 70729 61315 70849 61435 0 FreeSans 800 0 0 0 DATA[6]
port 15 nsew
flabel metal3 70729 58947 70849 59067 0 FreeSans 800 0 0 0 DATA[5]
port 16 nsew
flabel metal3 70729 56579 70849 56699 0 FreeSans 800 0 0 0 DATA[4]
port 17 nsew
flabel metal3 70729 54211 70849 54331 0 FreeSans 800 0 0 0 DATA[3]
port 18 nsew
flabel metal3 70729 51843 70849 51963 0 FreeSans 800 0 0 0 DATA[2]
port 20 nsew
flabel metal3 70729 49475 70849 49595 0 FreeSans 800 0 0 0 DATA[1]
port 21 nsew
flabel metal3 70729 47107 70849 47227 0 FreeSans 800 0 0 0 DATA[0]
port 22 nsew
flabel metal1 -10426 61158 -10396 61188 0 FreeSans 800 0 0 0 VINP
port 23 nsew
flabel metal1 -10422 59192 -10392 59222 0 FreeSans 800 0 0 0 VINN
port 24 nsew
flabel metal1 -11102 -688 -10846 -432 0 FreeSans 400 0 0 0 VSSR
port 25 nsew
flabel metal1 -11102 -1200 -10846 -944 0 FreeSans 400 0 0 0 VSSA
port 26 nsew
flabel metal1 -11102 -1713 -10846 -1457 0 FreeSans 400 0 0 0 VSSD
port 27 nsew
flabel metal1 -11039 121933 -10943 122029 0 FreeSans 400 0 0 0 VDDD
port 28 nsew
flabel metal3 70777 68452 70822 68500 0 FreeSans 400 0 0 0 DATA[9]
port 29 nsew
<< end >>
