magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect 238 1527 260 1561
rect 294 1527 332 1561
rect 366 1527 404 1561
rect 438 1527 476 1561
rect 510 1527 548 1561
rect 582 1527 620 1561
rect 654 1527 692 1561
rect 726 1527 764 1561
rect 798 1527 836 1561
rect 870 1527 908 1561
rect 942 1527 980 1561
rect 1014 1527 1052 1561
rect 1086 1527 1124 1561
rect 1158 1527 1196 1561
rect 1230 1527 1268 1561
rect 1302 1527 1340 1561
rect 1374 1527 1412 1561
rect 1446 1527 1484 1561
rect 1518 1527 1556 1561
rect 1590 1527 1628 1561
rect 1662 1527 1700 1561
rect 1734 1527 1772 1561
rect 1806 1527 1844 1561
rect 1878 1527 1916 1561
rect 1950 1527 1988 1561
rect 2022 1527 2060 1561
rect 2094 1527 2132 1561
rect 2166 1527 2204 1561
rect 2238 1527 2276 1561
rect 2310 1527 2348 1561
rect 2382 1527 2420 1561
rect 2454 1527 2492 1561
rect 2526 1527 2564 1561
rect 2598 1527 2636 1561
rect 2670 1527 2708 1561
rect 2742 1527 2780 1561
rect 2814 1527 2852 1561
rect 2886 1527 2924 1561
rect 2958 1527 2996 1561
rect 3030 1527 3068 1561
rect 3102 1527 3140 1561
rect 3174 1527 3212 1561
rect 3246 1527 3284 1561
rect 3318 1527 3356 1561
rect 3390 1527 3428 1561
rect 3462 1527 3500 1561
rect 3534 1527 3572 1561
rect 3606 1527 3644 1561
rect 3678 1527 3716 1561
rect 3750 1527 3788 1561
rect 3822 1527 3860 1561
rect 3894 1527 3932 1561
rect 3966 1527 4004 1561
rect 4038 1527 4076 1561
rect 4110 1527 4148 1561
rect 4182 1527 4220 1561
rect 4254 1527 4292 1561
rect 4326 1527 4364 1561
rect 4398 1527 4436 1561
rect 4470 1527 4508 1561
rect 4542 1527 4564 1561
rect 238 -123 250 -89
rect 284 -123 322 -89
rect 356 -123 394 -89
rect 428 -123 466 -89
rect 500 -123 538 -89
rect 572 -123 610 -89
rect 644 -123 682 -89
rect 716 -123 754 -89
rect 788 -123 826 -89
rect 860 -123 898 -89
rect 932 -123 970 -89
rect 1004 -123 1042 -89
rect 1076 -123 1114 -89
rect 1148 -123 1186 -89
rect 1220 -123 1258 -89
rect 1292 -123 1330 -89
rect 1364 -123 1402 -89
rect 1436 -123 1474 -89
rect 1508 -123 1546 -89
rect 1580 -123 1618 -89
rect 1652 -123 1690 -89
rect 1724 -123 1762 -89
rect 1796 -123 1834 -89
rect 1868 -123 1906 -89
rect 1940 -123 1978 -89
rect 2012 -123 2050 -89
rect 2084 -123 2122 -89
rect 2156 -123 2194 -89
rect 2228 -123 2266 -89
rect 2300 -123 2338 -89
rect 2372 -123 2384 -89
<< viali >>
rect 260 1527 294 1561
rect 332 1527 366 1561
rect 404 1527 438 1561
rect 476 1527 510 1561
rect 548 1527 582 1561
rect 620 1527 654 1561
rect 692 1527 726 1561
rect 764 1527 798 1561
rect 836 1527 870 1561
rect 908 1527 942 1561
rect 980 1527 1014 1561
rect 1052 1527 1086 1561
rect 1124 1527 1158 1561
rect 1196 1527 1230 1561
rect 1268 1527 1302 1561
rect 1340 1527 1374 1561
rect 1412 1527 1446 1561
rect 1484 1527 1518 1561
rect 1556 1527 1590 1561
rect 1628 1527 1662 1561
rect 1700 1527 1734 1561
rect 1772 1527 1806 1561
rect 1844 1527 1878 1561
rect 1916 1527 1950 1561
rect 1988 1527 2022 1561
rect 2060 1527 2094 1561
rect 2132 1527 2166 1561
rect 2204 1527 2238 1561
rect 2276 1527 2310 1561
rect 2348 1527 2382 1561
rect 2420 1527 2454 1561
rect 2492 1527 2526 1561
rect 2564 1527 2598 1561
rect 2636 1527 2670 1561
rect 2708 1527 2742 1561
rect 2780 1527 2814 1561
rect 2852 1527 2886 1561
rect 2924 1527 2958 1561
rect 2996 1527 3030 1561
rect 3068 1527 3102 1561
rect 3140 1527 3174 1561
rect 3212 1527 3246 1561
rect 3284 1527 3318 1561
rect 3356 1527 3390 1561
rect 3428 1527 3462 1561
rect 3500 1527 3534 1561
rect 3572 1527 3606 1561
rect 3644 1527 3678 1561
rect 3716 1527 3750 1561
rect 3788 1527 3822 1561
rect 3860 1527 3894 1561
rect 3932 1527 3966 1561
rect 4004 1527 4038 1561
rect 4076 1527 4110 1561
rect 4148 1527 4182 1561
rect 4220 1527 4254 1561
rect 4292 1527 4326 1561
rect 4364 1527 4398 1561
rect 4436 1527 4470 1561
rect 4508 1527 4542 1561
rect 250 -123 284 -89
rect 322 -123 356 -89
rect 394 -123 428 -89
rect 466 -123 500 -89
rect 538 -123 572 -89
rect 610 -123 644 -89
rect 682 -123 716 -89
rect 754 -123 788 -89
rect 826 -123 860 -89
rect 898 -123 932 -89
rect 970 -123 1004 -89
rect 1042 -123 1076 -89
rect 1114 -123 1148 -89
rect 1186 -123 1220 -89
rect 1258 -123 1292 -89
rect 1330 -123 1364 -89
rect 1402 -123 1436 -89
rect 1474 -123 1508 -89
rect 1546 -123 1580 -89
rect 1618 -123 1652 -89
rect 1690 -123 1724 -89
rect 1762 -123 1796 -89
rect 1834 -123 1868 -89
rect 1906 -123 1940 -89
rect 1978 -123 2012 -89
rect 2050 -123 2084 -89
rect 2122 -123 2156 -89
rect 2194 -123 2228 -89
rect 2266 -123 2300 -89
rect 2338 -123 2372 -89
<< metal1 >>
rect 106 1561 4696 1597
rect 106 1527 260 1561
rect 294 1527 332 1561
rect 366 1527 404 1561
rect 438 1527 476 1561
rect 510 1527 548 1561
rect 582 1527 620 1561
rect 654 1527 692 1561
rect 726 1527 764 1561
rect 798 1527 836 1561
rect 870 1527 908 1561
rect 942 1527 980 1561
rect 1014 1527 1052 1561
rect 1086 1527 1124 1561
rect 1158 1527 1196 1561
rect 1230 1527 1268 1561
rect 1302 1527 1340 1561
rect 1374 1527 1412 1561
rect 1446 1527 1484 1561
rect 1518 1527 1556 1561
rect 1590 1527 1628 1561
rect 1662 1527 1700 1561
rect 1734 1527 1772 1561
rect 1806 1527 1844 1561
rect 1878 1527 1916 1561
rect 1950 1527 1988 1561
rect 2022 1527 2060 1561
rect 2094 1527 2132 1561
rect 2166 1527 2204 1561
rect 2238 1527 2276 1561
rect 2310 1527 2348 1561
rect 2382 1527 2420 1561
rect 2454 1527 2492 1561
rect 2526 1527 2564 1561
rect 2598 1527 2636 1561
rect 2670 1527 2708 1561
rect 2742 1527 2780 1561
rect 2814 1527 2852 1561
rect 2886 1527 2924 1561
rect 2958 1527 2996 1561
rect 3030 1527 3068 1561
rect 3102 1527 3140 1561
rect 3174 1527 3212 1561
rect 3246 1527 3284 1561
rect 3318 1527 3356 1561
rect 3390 1527 3428 1561
rect 3462 1527 3500 1561
rect 3534 1527 3572 1561
rect 3606 1527 3644 1561
rect 3678 1527 3716 1561
rect 3750 1527 3788 1561
rect 3822 1527 3860 1561
rect 3894 1527 3932 1561
rect 3966 1527 4004 1561
rect 4038 1527 4076 1561
rect 4110 1527 4148 1561
rect 4182 1527 4220 1561
rect 4254 1527 4292 1561
rect 4326 1527 4364 1561
rect 4398 1527 4436 1561
rect 4470 1527 4508 1561
rect 4542 1527 4696 1561
rect 106 1521 4696 1527
rect 325 1447 4477 1521
rect 106 1377 284 1401
rect 106 1325 176 1377
rect 228 1325 284 1377
rect 106 1301 284 1325
rect 325 1061 4477 1255
rect 106 915 284 1015
rect 316 569 4696 869
rect 106 423 284 523
rect 316 183 2306 377
rect 166 113 284 137
rect 166 61 176 113
rect 228 61 284 113
rect 166 37 284 61
rect 316 -83 2306 -9
rect 106 -89 4696 -83
rect 106 -123 250 -89
rect 284 -123 322 -89
rect 356 -123 394 -89
rect 428 -123 466 -89
rect 500 -123 538 -89
rect 572 -123 610 -89
rect 644 -123 682 -89
rect 716 -123 754 -89
rect 788 -123 826 -89
rect 860 -123 898 -89
rect 932 -123 970 -89
rect 1004 -123 1042 -89
rect 1076 -123 1114 -89
rect 1148 -123 1186 -89
rect 1220 -123 1258 -89
rect 1292 -123 1330 -89
rect 1364 -123 1402 -89
rect 1436 -123 1474 -89
rect 1508 -123 1546 -89
rect 1580 -123 1618 -89
rect 1652 -123 1690 -89
rect 1724 -123 1762 -89
rect 1796 -123 1834 -89
rect 1868 -123 1906 -89
rect 1940 -123 1978 -89
rect 2012 -123 2050 -89
rect 2084 -123 2122 -89
rect 2156 -123 2194 -89
rect 2228 -123 2266 -89
rect 2300 -123 2338 -89
rect 2372 -123 4696 -89
rect 106 -159 4696 -123
<< via1 >>
rect 176 1325 228 1377
rect 176 61 228 113
<< metal2 >>
rect 176 1377 228 1411
rect 176 113 228 1325
rect 176 27 228 61
use sky130_fd_pr__nfet_01v8_55NS9E  sky130_fd_pr__nfet_01v8_55NS9E_0
timestamp 1750100919
transform 0 1 1311 -1 0 87
box -236 -1195 236 1195
use sky130_fd_pr__pfet_01v8_D9QZ56  sky130_fd_pr__pfet_01v8_D9QZ56_0
timestamp 1750100919
transform 0 1 2401 -1 0 965
box -246 -2295 246 2295
use sky130_fd_pr__pfet_01v8_D9QZ56  XM1
timestamp 1750100919
transform 0 1 2401 -1 0 1351
box -246 -2295 246 2295
use sky130_fd_pr__nfet_01v8_55NS9E  XM3
timestamp 1750100919
transform 0 1 1311 -1 0 473
box -236 -1195 236 1195
<< labels >>
flabel metal1 s 106 1521 238 1597 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 106 1301 176 1401 0 FreeSans 500 0 0 0 IN
port 2 nsew
flabel metal1 s 106 915 284 1015 0 FreeSans 500 0 0 0 CKB
port 3 nsew
flabel metal1 s 106 423 284 523 0 FreeSans 500 0 0 0 CK
port 4 nsew
flabel metal1 s 106 -159 238 -83 0 FreeSans 500 0 0 0 VSS
port 5 nsew
flabel metal1 s 4514 655 4628 703 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
