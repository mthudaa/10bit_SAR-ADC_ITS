magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< nwell >>
rect 3369 -56 4107 1053
rect 3369 -115 4033 -56
<< locali >>
rect -9799 1913 -9768 1947
rect -9734 1913 -9672 1947
rect -9638 1913 -9576 1947
rect -9542 1913 -9480 1947
rect -9446 1913 -9384 1947
rect -9350 1913 -9288 1947
rect -9254 1913 -9192 1947
rect -9158 1913 -9096 1947
rect -9062 1913 -9000 1947
rect -8966 1913 -8904 1947
rect -8870 1913 -8808 1947
rect -8774 1913 -8712 1947
rect -8678 1913 -8616 1947
rect -8582 1913 -8520 1947
rect -8486 1913 -8424 1947
rect -8390 1913 -8328 1947
rect -8294 1913 -8232 1947
rect -8198 1913 -8136 1947
rect -8102 1913 -8040 1947
rect -8006 1913 -7944 1947
rect -7910 1913 -7848 1947
rect -7814 1913 -7752 1947
rect -7718 1913 -7656 1947
rect -7622 1913 -7560 1947
rect -7526 1913 -7464 1947
rect -7430 1913 -7368 1947
rect -7334 1913 -7272 1947
rect -7238 1913 -7176 1947
rect -7142 1913 -7080 1947
rect -7046 1913 -6984 1947
rect -6950 1913 -6888 1947
rect -6854 1913 -6792 1947
rect -6758 1913 -6696 1947
rect -6662 1913 -6600 1947
rect -6566 1913 -6504 1947
rect -6470 1913 -6408 1947
rect -6374 1913 -6312 1947
rect -6278 1913 -6216 1947
rect -6182 1913 -6120 1947
rect -6086 1913 -6024 1947
rect -5990 1913 -5928 1947
rect -5894 1913 -5832 1947
rect -5798 1913 -5736 1947
rect -5702 1913 -5640 1947
rect -5606 1913 -5544 1947
rect -5510 1913 -5448 1947
rect -5414 1913 -5352 1947
rect -5318 1913 -5256 1947
rect -5222 1913 -5160 1947
rect -5126 1913 -5064 1947
rect -5030 1913 -4968 1947
rect -4934 1913 -4872 1947
rect -4838 1913 -4776 1947
rect -4742 1913 -4680 1947
rect -4646 1913 -4584 1947
rect -4550 1913 -4488 1947
rect -4454 1913 -4392 1947
rect -4358 1913 -4296 1947
rect -4262 1913 -4200 1947
rect -4166 1913 -4104 1947
rect -4070 1913 -4008 1947
rect -3974 1913 -3912 1947
rect -3878 1913 -3816 1947
rect -3782 1913 -3720 1947
rect -3686 1913 -3624 1947
rect -3590 1913 -3528 1947
rect -3494 1913 -3432 1947
rect -3398 1913 -3336 1947
rect -3302 1913 -3240 1947
rect -3206 1913 -3144 1947
rect -3110 1913 -3048 1947
rect -3014 1913 -2952 1947
rect -2918 1913 -2856 1947
rect -2822 1913 -2760 1947
rect -2726 1913 -2664 1947
rect -2630 1913 -2568 1947
rect -2534 1913 -2472 1947
rect -2438 1913 -2376 1947
rect -2342 1913 -2280 1947
rect -2246 1913 -2184 1947
rect -2150 1913 -2088 1947
rect -2054 1913 -1992 1947
rect -1958 1913 -1896 1947
rect -1862 1913 -1800 1947
rect -1766 1913 -1704 1947
rect -1670 1913 -1608 1947
rect -1574 1913 -1512 1947
rect -1478 1913 -1416 1947
rect -1382 1913 -1320 1947
rect -1286 1913 -1224 1947
rect -1190 1913 -1128 1947
rect -1094 1913 -1032 1947
rect -998 1913 -936 1947
rect -902 1913 -840 1947
rect -806 1913 -744 1947
rect -710 1913 -648 1947
rect -614 1913 -552 1947
rect -518 1913 -456 1947
rect -422 1913 -360 1947
rect -326 1913 -264 1947
rect -230 1913 -168 1947
rect -134 1913 -72 1947
rect -38 1913 24 1947
rect 58 1913 120 1947
rect 154 1913 216 1947
rect 250 1913 312 1947
rect 346 1913 408 1947
rect 442 1913 504 1947
rect 538 1913 600 1947
rect 634 1913 696 1947
rect 730 1913 792 1947
rect 826 1913 888 1947
rect 922 1913 984 1947
rect 1018 1913 1080 1947
rect 1114 1913 1176 1947
rect 1210 1913 1272 1947
rect 1306 1913 1368 1947
rect 1402 1913 1464 1947
rect 1498 1913 1529 1947
rect 79 367 237 1913
rect 79 333 105 367
rect 139 333 177 367
rect 211 333 237 367
rect 3721 466 3755 471
rect 3721 394 3755 432
rect 3721 322 3755 360
rect 3721 250 3755 288
rect 3721 178 3755 216
rect 3721 139 3755 144
rect 237 -3689 263 -3655
rect 297 -3689 335 -3655
rect 369 -3689 395 -3655
rect -9799 -4101 -9768 -4067
rect -9734 -4101 -9672 -4067
rect -9638 -4101 -9576 -4067
rect -9542 -4101 -9480 -4067
rect -9446 -4101 -9384 -4067
rect -9350 -4101 -9288 -4067
rect -9254 -4101 -9192 -4067
rect -9158 -4101 -9096 -4067
rect -9062 -4101 -9000 -4067
rect -8966 -4101 -8904 -4067
rect -8870 -4101 -8808 -4067
rect -8774 -4101 -8712 -4067
rect -8678 -4101 -8616 -4067
rect -8582 -4101 -8520 -4067
rect -8486 -4101 -8424 -4067
rect -8390 -4101 -8328 -4067
rect -8294 -4101 -8232 -4067
rect -8198 -4101 -8136 -4067
rect -8102 -4101 -8040 -4067
rect -8006 -4101 -7944 -4067
rect -7910 -4101 -7848 -4067
rect -7814 -4101 -7752 -4067
rect -7718 -4101 -7656 -4067
rect -7622 -4101 -7560 -4067
rect -7526 -4101 -7464 -4067
rect -7430 -4101 -7368 -4067
rect -7334 -4101 -7272 -4067
rect -7238 -4101 -7176 -4067
rect -7142 -4101 -7080 -4067
rect -7046 -4101 -6984 -4067
rect -6950 -4101 -6888 -4067
rect -6854 -4101 -6792 -4067
rect -6758 -4101 -6696 -4067
rect -6662 -4101 -6600 -4067
rect -6566 -4101 -6504 -4067
rect -6470 -4101 -6408 -4067
rect -6374 -4101 -6312 -4067
rect -6278 -4101 -6216 -4067
rect -6182 -4101 -6120 -4067
rect -6086 -4101 -6024 -4067
rect -5990 -4101 -5928 -4067
rect -5894 -4101 -5832 -4067
rect -5798 -4101 -5736 -4067
rect -5702 -4101 -5640 -4067
rect -5606 -4101 -5544 -4067
rect -5510 -4101 -5448 -4067
rect -5414 -4101 -5352 -4067
rect -5318 -4101 -5256 -4067
rect -5222 -4101 -5160 -4067
rect -5126 -4101 -5064 -4067
rect -5030 -4101 -4968 -4067
rect -4934 -4101 -4872 -4067
rect -4838 -4101 -4776 -4067
rect -4742 -4101 -4680 -4067
rect -4646 -4101 -4584 -4067
rect -4550 -4101 -4488 -4067
rect -4454 -4101 -4392 -4067
rect -4358 -4101 -4296 -4067
rect -4262 -4101 -4200 -4067
rect -4166 -4101 -4104 -4067
rect -4070 -4101 -4008 -4067
rect -3974 -4101 -3912 -4067
rect -3878 -4101 -3816 -4067
rect -3782 -4101 -3720 -4067
rect -3686 -4101 -3624 -4067
rect -3590 -4101 -3528 -4067
rect -3494 -4101 -3432 -4067
rect -3398 -4101 -3336 -4067
rect -3302 -4101 -3240 -4067
rect -3206 -4101 -3144 -4067
rect -3110 -4101 -3048 -4067
rect -3014 -4101 -2952 -4067
rect -2918 -4101 -2856 -4067
rect -2822 -4101 -2760 -4067
rect -2726 -4101 -2664 -4067
rect -2630 -4101 -2568 -4067
rect -2534 -4101 -2472 -4067
rect -2438 -4101 -2376 -4067
rect -2342 -4101 -2280 -4067
rect -2246 -4101 -2184 -4067
rect -2150 -4101 -2088 -4067
rect -2054 -4101 -1992 -4067
rect -1958 -4101 -1896 -4067
rect -1862 -4101 -1800 -4067
rect -1766 -4101 -1704 -4067
rect -1670 -4101 -1608 -4067
rect -1574 -4101 -1512 -4067
rect -1478 -4101 -1416 -4067
rect -1382 -4101 -1320 -4067
rect -1286 -4101 -1224 -4067
rect -1190 -4101 -1128 -4067
rect -1094 -4101 -1032 -4067
rect -998 -4101 -936 -4067
rect -902 -4101 -840 -4067
rect -806 -4101 -744 -4067
rect -710 -4101 -648 -4067
rect -614 -4101 -552 -4067
rect -518 -4101 -456 -4067
rect -422 -4101 -360 -4067
rect -326 -4101 -264 -4067
rect -230 -4101 -168 -4067
rect -134 -4101 -72 -4067
rect -38 -4101 24 -4067
rect 58 -4101 120 -4067
rect 154 -4101 216 -4067
rect 250 -4101 312 -4067
rect 346 -4101 408 -4067
rect 442 -4101 504 -4067
rect 538 -4101 600 -4067
rect 634 -4101 696 -4067
rect 730 -4101 792 -4067
rect 826 -4101 888 -4067
rect 922 -4101 984 -4067
rect 1018 -4101 1080 -4067
rect 1114 -4101 1176 -4067
rect 1210 -4101 1272 -4067
rect 1306 -4101 1368 -4067
rect 1402 -4101 1464 -4067
rect 1498 -4101 1529 -4067
<< viali >>
rect -9768 1913 -9734 1947
rect -9672 1913 -9638 1947
rect -9576 1913 -9542 1947
rect -9480 1913 -9446 1947
rect -9384 1913 -9350 1947
rect -9288 1913 -9254 1947
rect -9192 1913 -9158 1947
rect -9096 1913 -9062 1947
rect -9000 1913 -8966 1947
rect -8904 1913 -8870 1947
rect -8808 1913 -8774 1947
rect -8712 1913 -8678 1947
rect -8616 1913 -8582 1947
rect -8520 1913 -8486 1947
rect -8424 1913 -8390 1947
rect -8328 1913 -8294 1947
rect -8232 1913 -8198 1947
rect -8136 1913 -8102 1947
rect -8040 1913 -8006 1947
rect -7944 1913 -7910 1947
rect -7848 1913 -7814 1947
rect -7752 1913 -7718 1947
rect -7656 1913 -7622 1947
rect -7560 1913 -7526 1947
rect -7464 1913 -7430 1947
rect -7368 1913 -7334 1947
rect -7272 1913 -7238 1947
rect -7176 1913 -7142 1947
rect -7080 1913 -7046 1947
rect -6984 1913 -6950 1947
rect -6888 1913 -6854 1947
rect -6792 1913 -6758 1947
rect -6696 1913 -6662 1947
rect -6600 1913 -6566 1947
rect -6504 1913 -6470 1947
rect -6408 1913 -6374 1947
rect -6312 1913 -6278 1947
rect -6216 1913 -6182 1947
rect -6120 1913 -6086 1947
rect -6024 1913 -5990 1947
rect -5928 1913 -5894 1947
rect -5832 1913 -5798 1947
rect -5736 1913 -5702 1947
rect -5640 1913 -5606 1947
rect -5544 1913 -5510 1947
rect -5448 1913 -5414 1947
rect -5352 1913 -5318 1947
rect -5256 1913 -5222 1947
rect -5160 1913 -5126 1947
rect -5064 1913 -5030 1947
rect -4968 1913 -4934 1947
rect -4872 1913 -4838 1947
rect -4776 1913 -4742 1947
rect -4680 1913 -4646 1947
rect -4584 1913 -4550 1947
rect -4488 1913 -4454 1947
rect -4392 1913 -4358 1947
rect -4296 1913 -4262 1947
rect -4200 1913 -4166 1947
rect -4104 1913 -4070 1947
rect -4008 1913 -3974 1947
rect -3912 1913 -3878 1947
rect -3816 1913 -3782 1947
rect -3720 1913 -3686 1947
rect -3624 1913 -3590 1947
rect -3528 1913 -3494 1947
rect -3432 1913 -3398 1947
rect -3336 1913 -3302 1947
rect -3240 1913 -3206 1947
rect -3144 1913 -3110 1947
rect -3048 1913 -3014 1947
rect -2952 1913 -2918 1947
rect -2856 1913 -2822 1947
rect -2760 1913 -2726 1947
rect -2664 1913 -2630 1947
rect -2568 1913 -2534 1947
rect -2472 1913 -2438 1947
rect -2376 1913 -2342 1947
rect -2280 1913 -2246 1947
rect -2184 1913 -2150 1947
rect -2088 1913 -2054 1947
rect -1992 1913 -1958 1947
rect -1896 1913 -1862 1947
rect -1800 1913 -1766 1947
rect -1704 1913 -1670 1947
rect -1608 1913 -1574 1947
rect -1512 1913 -1478 1947
rect -1416 1913 -1382 1947
rect -1320 1913 -1286 1947
rect -1224 1913 -1190 1947
rect -1128 1913 -1094 1947
rect -1032 1913 -998 1947
rect -936 1913 -902 1947
rect -840 1913 -806 1947
rect -744 1913 -710 1947
rect -648 1913 -614 1947
rect -552 1913 -518 1947
rect -456 1913 -422 1947
rect -360 1913 -326 1947
rect -264 1913 -230 1947
rect -168 1913 -134 1947
rect -72 1913 -38 1947
rect 24 1913 58 1947
rect 120 1913 154 1947
rect 216 1913 250 1947
rect 312 1913 346 1947
rect 408 1913 442 1947
rect 504 1913 538 1947
rect 600 1913 634 1947
rect 696 1913 730 1947
rect 792 1913 826 1947
rect 888 1913 922 1947
rect 984 1913 1018 1947
rect 1080 1913 1114 1947
rect 1176 1913 1210 1947
rect 1272 1913 1306 1947
rect 1368 1913 1402 1947
rect 1464 1913 1498 1947
rect 105 333 139 367
rect 177 333 211 367
rect 3721 432 3755 466
rect 3721 360 3755 394
rect 3721 288 3755 322
rect 3721 216 3755 250
rect 3721 144 3755 178
rect 263 -3689 297 -3655
rect 335 -3689 369 -3655
rect -9768 -4101 -9734 -4067
rect -9672 -4101 -9638 -4067
rect -9576 -4101 -9542 -4067
rect -9480 -4101 -9446 -4067
rect -9384 -4101 -9350 -4067
rect -9288 -4101 -9254 -4067
rect -9192 -4101 -9158 -4067
rect -9096 -4101 -9062 -4067
rect -9000 -4101 -8966 -4067
rect -8904 -4101 -8870 -4067
rect -8808 -4101 -8774 -4067
rect -8712 -4101 -8678 -4067
rect -8616 -4101 -8582 -4067
rect -8520 -4101 -8486 -4067
rect -8424 -4101 -8390 -4067
rect -8328 -4101 -8294 -4067
rect -8232 -4101 -8198 -4067
rect -8136 -4101 -8102 -4067
rect -8040 -4101 -8006 -4067
rect -7944 -4101 -7910 -4067
rect -7848 -4101 -7814 -4067
rect -7752 -4101 -7718 -4067
rect -7656 -4101 -7622 -4067
rect -7560 -4101 -7526 -4067
rect -7464 -4101 -7430 -4067
rect -7368 -4101 -7334 -4067
rect -7272 -4101 -7238 -4067
rect -7176 -4101 -7142 -4067
rect -7080 -4101 -7046 -4067
rect -6984 -4101 -6950 -4067
rect -6888 -4101 -6854 -4067
rect -6792 -4101 -6758 -4067
rect -6696 -4101 -6662 -4067
rect -6600 -4101 -6566 -4067
rect -6504 -4101 -6470 -4067
rect -6408 -4101 -6374 -4067
rect -6312 -4101 -6278 -4067
rect -6216 -4101 -6182 -4067
rect -6120 -4101 -6086 -4067
rect -6024 -4101 -5990 -4067
rect -5928 -4101 -5894 -4067
rect -5832 -4101 -5798 -4067
rect -5736 -4101 -5702 -4067
rect -5640 -4101 -5606 -4067
rect -5544 -4101 -5510 -4067
rect -5448 -4101 -5414 -4067
rect -5352 -4101 -5318 -4067
rect -5256 -4101 -5222 -4067
rect -5160 -4101 -5126 -4067
rect -5064 -4101 -5030 -4067
rect -4968 -4101 -4934 -4067
rect -4872 -4101 -4838 -4067
rect -4776 -4101 -4742 -4067
rect -4680 -4101 -4646 -4067
rect -4584 -4101 -4550 -4067
rect -4488 -4101 -4454 -4067
rect -4392 -4101 -4358 -4067
rect -4296 -4101 -4262 -4067
rect -4200 -4101 -4166 -4067
rect -4104 -4101 -4070 -4067
rect -4008 -4101 -3974 -4067
rect -3912 -4101 -3878 -4067
rect -3816 -4101 -3782 -4067
rect -3720 -4101 -3686 -4067
rect -3624 -4101 -3590 -4067
rect -3528 -4101 -3494 -4067
rect -3432 -4101 -3398 -4067
rect -3336 -4101 -3302 -4067
rect -3240 -4101 -3206 -4067
rect -3144 -4101 -3110 -4067
rect -3048 -4101 -3014 -4067
rect -2952 -4101 -2918 -4067
rect -2856 -4101 -2822 -4067
rect -2760 -4101 -2726 -4067
rect -2664 -4101 -2630 -4067
rect -2568 -4101 -2534 -4067
rect -2472 -4101 -2438 -4067
rect -2376 -4101 -2342 -4067
rect -2280 -4101 -2246 -4067
rect -2184 -4101 -2150 -4067
rect -2088 -4101 -2054 -4067
rect -1992 -4101 -1958 -4067
rect -1896 -4101 -1862 -4067
rect -1800 -4101 -1766 -4067
rect -1704 -4101 -1670 -4067
rect -1608 -4101 -1574 -4067
rect -1512 -4101 -1478 -4067
rect -1416 -4101 -1382 -4067
rect -1320 -4101 -1286 -4067
rect -1224 -4101 -1190 -4067
rect -1128 -4101 -1094 -4067
rect -1032 -4101 -998 -4067
rect -936 -4101 -902 -4067
rect -840 -4101 -806 -4067
rect -744 -4101 -710 -4067
rect -648 -4101 -614 -4067
rect -552 -4101 -518 -4067
rect -456 -4101 -422 -4067
rect -360 -4101 -326 -4067
rect -264 -4101 -230 -4067
rect -168 -4101 -134 -4067
rect -72 -4101 -38 -4067
rect 24 -4101 58 -4067
rect 120 -4101 154 -4067
rect 216 -4101 250 -4067
rect 312 -4101 346 -4067
rect 408 -4101 442 -4067
rect 504 -4101 538 -4067
rect 600 -4101 634 -4067
rect 696 -4101 730 -4067
rect 792 -4101 826 -4067
rect 888 -4101 922 -4067
rect 984 -4101 1018 -4067
rect 1080 -4101 1114 -4067
rect 1176 -4101 1210 -4067
rect 1272 -4101 1306 -4067
rect 1368 -4101 1402 -4067
rect 1464 -4101 1498 -4067
<< metal1 >>
rect -9799 1947 1529 1978
rect -9799 1913 -9768 1947
rect -9734 1913 -9672 1947
rect -9638 1913 -9576 1947
rect -9542 1913 -9480 1947
rect -9446 1913 -9384 1947
rect -9350 1913 -9288 1947
rect -9254 1913 -9192 1947
rect -9158 1913 -9096 1947
rect -9062 1913 -9000 1947
rect -8966 1913 -8904 1947
rect -8870 1913 -8808 1947
rect -8774 1913 -8712 1947
rect -8678 1913 -8616 1947
rect -8582 1913 -8520 1947
rect -8486 1913 -8424 1947
rect -8390 1913 -8328 1947
rect -8294 1913 -8232 1947
rect -8198 1913 -8136 1947
rect -8102 1913 -8040 1947
rect -8006 1913 -7944 1947
rect -7910 1913 -7848 1947
rect -7814 1913 -7752 1947
rect -7718 1913 -7656 1947
rect -7622 1913 -7560 1947
rect -7526 1913 -7464 1947
rect -7430 1913 -7368 1947
rect -7334 1913 -7272 1947
rect -7238 1913 -7176 1947
rect -7142 1913 -7080 1947
rect -7046 1913 -6984 1947
rect -6950 1913 -6888 1947
rect -6854 1913 -6792 1947
rect -6758 1913 -6696 1947
rect -6662 1913 -6600 1947
rect -6566 1913 -6504 1947
rect -6470 1913 -6408 1947
rect -6374 1913 -6312 1947
rect -6278 1913 -6216 1947
rect -6182 1913 -6120 1947
rect -6086 1913 -6024 1947
rect -5990 1913 -5928 1947
rect -5894 1913 -5832 1947
rect -5798 1913 -5736 1947
rect -5702 1913 -5640 1947
rect -5606 1913 -5544 1947
rect -5510 1913 -5448 1947
rect -5414 1913 -5352 1947
rect -5318 1913 -5256 1947
rect -5222 1913 -5160 1947
rect -5126 1913 -5064 1947
rect -5030 1913 -4968 1947
rect -4934 1913 -4872 1947
rect -4838 1913 -4776 1947
rect -4742 1913 -4680 1947
rect -4646 1913 -4584 1947
rect -4550 1913 -4488 1947
rect -4454 1913 -4392 1947
rect -4358 1913 -4296 1947
rect -4262 1913 -4200 1947
rect -4166 1913 -4104 1947
rect -4070 1913 -4008 1947
rect -3974 1913 -3912 1947
rect -3878 1913 -3816 1947
rect -3782 1913 -3720 1947
rect -3686 1913 -3624 1947
rect -3590 1913 -3528 1947
rect -3494 1913 -3432 1947
rect -3398 1913 -3336 1947
rect -3302 1913 -3240 1947
rect -3206 1913 -3144 1947
rect -3110 1913 -3048 1947
rect -3014 1913 -2952 1947
rect -2918 1913 -2856 1947
rect -2822 1913 -2760 1947
rect -2726 1913 -2664 1947
rect -2630 1913 -2568 1947
rect -2534 1913 -2472 1947
rect -2438 1913 -2376 1947
rect -2342 1913 -2280 1947
rect -2246 1913 -2184 1947
rect -2150 1913 -2088 1947
rect -2054 1913 -1992 1947
rect -1958 1913 -1896 1947
rect -1862 1913 -1800 1947
rect -1766 1913 -1704 1947
rect -1670 1913 -1608 1947
rect -1574 1913 -1512 1947
rect -1478 1913 -1416 1947
rect -1382 1913 -1320 1947
rect -1286 1913 -1224 1947
rect -1190 1913 -1128 1947
rect -1094 1913 -1032 1947
rect -998 1913 -936 1947
rect -902 1913 -840 1947
rect -806 1913 -744 1947
rect -710 1913 -648 1947
rect -614 1913 -552 1947
rect -518 1913 -456 1947
rect -422 1913 -360 1947
rect -326 1913 -264 1947
rect -230 1913 -168 1947
rect -134 1913 -72 1947
rect -38 1913 24 1947
rect 58 1913 120 1947
rect 154 1913 216 1947
rect 250 1913 312 1947
rect 346 1913 408 1947
rect 442 1913 504 1947
rect 538 1913 600 1947
rect 634 1913 696 1947
rect 730 1913 792 1947
rect 826 1913 888 1947
rect 922 1913 984 1947
rect 1018 1913 1080 1947
rect 1114 1913 1176 1947
rect 1210 1913 1272 1947
rect 1306 1913 1368 1947
rect 1402 1913 1464 1947
rect 1498 1913 1529 1947
rect -9799 1882 1529 1913
rect 79 1053 237 1882
rect 79 981 3523 1053
rect 79 507 237 981
rect 79 455 448 507
rect 500 455 510 507
rect 79 373 237 455
rect 67 367 249 373
rect 67 333 105 367
rect 139 333 177 367
rect 211 333 249 367
rect 67 327 249 333
rect 91 220 137 327
rect 215 237 287 254
rect 215 185 225 237
rect 277 185 287 237
rect 215 173 287 185
rect 215 121 225 173
rect 277 121 287 173
rect 215 104 287 121
rect -281 33 -157 59
rect -281 -19 -245 33
rect -193 -19 -157 33
rect 122 11 132 63
rect 184 11 194 63
rect 3451 33 3523 981
rect 3551 874 3963 926
rect 4015 874 4025 926
rect 3607 466 3870 505
rect 3607 459 3721 466
rect 3755 459 3870 466
rect 3607 407 3712 459
rect 3764 407 3870 459
rect 3607 395 3870 407
rect 3607 343 3712 395
rect 3764 343 3870 395
rect 3607 331 3870 343
rect 3607 279 3712 331
rect 3764 279 3870 331
rect 3607 267 3870 279
rect 3607 215 3712 267
rect 3764 215 3870 267
rect 3607 203 3870 215
rect 3607 151 3712 203
rect 3764 151 3870 203
rect 3607 144 3721 151
rect 3755 144 3870 151
rect 3607 105 3870 144
rect 3953 491 4025 505
rect 3953 439 3963 491
rect 4015 439 4025 491
rect 3953 427 4025 439
rect 3953 375 3963 427
rect 4015 375 4025 427
rect 3953 363 4025 375
rect 3953 311 3963 363
rect 4015 311 4025 363
rect 3953 299 4025 311
rect 3953 247 3963 299
rect 4015 247 4025 299
rect 3953 235 4025 247
rect 3953 183 3963 235
rect 4015 183 4025 235
rect 3953 171 4025 183
rect 3953 119 3963 171
rect 4015 119 4025 171
rect 3953 105 4025 119
rect 3860 12 3870 64
rect 3922 12 3932 64
rect -281 -45 -157 -19
rect -281 -97 3712 -45
rect 3764 -97 3774 -45
rect -281 -123 -157 -97
rect -281 -175 -245 -123
rect -193 -175 -157 -123
rect -281 -201 -157 -175
rect 215 -201 225 -149
rect 277 -201 857 -149
rect 909 -201 3870 -149
rect 3922 -201 3932 -149
rect 122 -293 132 -241
rect 184 -293 194 -241
rect 438 -293 448 -241
rect 500 -293 510 -241
rect 29 -349 101 -325
rect 29 -401 39 -349
rect 91 -401 101 -349
rect 29 -425 101 -401
rect 215 -349 287 -325
rect 215 -401 225 -349
rect 277 -401 287 -349
rect 215 -425 287 -401
rect 345 -345 417 -325
rect 345 -397 355 -345
rect 407 -397 417 -345
rect 345 -409 417 -397
rect 345 -461 355 -409
rect 407 -461 417 -409
rect 345 -473 417 -461
rect 345 -525 355 -473
rect 407 -525 417 -473
rect 345 -537 417 -525
rect 345 -589 355 -537
rect 407 -589 417 -537
rect 345 -601 417 -589
rect 345 -653 355 -601
rect 407 -653 417 -601
rect 345 -665 417 -653
rect 345 -717 355 -665
rect 407 -717 417 -665
rect 345 -729 417 -717
rect 345 -781 355 -729
rect 407 -781 417 -729
rect 345 -793 417 -781
rect 345 -845 355 -793
rect 407 -845 417 -793
rect 345 -857 417 -845
rect 345 -909 355 -857
rect 407 -909 417 -857
rect 345 -921 417 -909
rect 345 -973 355 -921
rect 407 -973 417 -921
rect 345 -985 417 -973
rect 345 -1037 355 -985
rect 407 -1037 417 -985
rect 345 -1049 417 -1037
rect 345 -1101 355 -1049
rect 407 -1101 417 -1049
rect 345 -1113 417 -1101
rect 345 -1165 355 -1113
rect 407 -1165 417 -1113
rect 345 -1177 417 -1165
rect 345 -1229 355 -1177
rect 407 -1229 417 -1177
rect 345 -1241 417 -1229
rect 345 -1293 355 -1241
rect 407 -1293 417 -1241
rect 345 -1305 417 -1293
rect 345 -1357 355 -1305
rect 407 -1357 417 -1305
rect 345 -1369 417 -1357
rect 345 -1421 355 -1369
rect 407 -1421 417 -1369
rect 345 -1433 417 -1421
rect 345 -1485 355 -1433
rect 407 -1485 417 -1433
rect 345 -1497 417 -1485
rect 345 -1549 355 -1497
rect 407 -1549 417 -1497
rect 345 -1561 417 -1549
rect 345 -1613 355 -1561
rect 407 -1613 417 -1561
rect 345 -1625 417 -1613
rect 345 -1677 355 -1625
rect 407 -1677 417 -1625
rect 345 -1689 417 -1677
rect 345 -1741 355 -1689
rect 407 -1741 417 -1689
rect 345 -1753 417 -1741
rect 345 -1805 355 -1753
rect 407 -1805 417 -1753
rect 345 -1825 417 -1805
rect 531 -356 3963 -325
rect 531 -408 541 -356
rect 593 -377 3963 -356
rect 4015 -377 4025 -325
rect 593 -408 603 -377
rect 531 -420 603 -408
rect 531 -472 541 -420
rect 593 -472 603 -420
rect 531 -484 603 -472
rect 531 -536 541 -484
rect 593 -536 603 -484
rect 531 -548 603 -536
rect 531 -600 541 -548
rect 593 -600 603 -548
rect 531 -612 603 -600
rect 531 -664 541 -612
rect 593 -664 603 -612
rect 531 -676 603 -664
rect 531 -728 541 -676
rect 593 -728 603 -676
rect 531 -740 603 -728
rect 531 -792 541 -740
rect 593 -792 603 -740
rect 531 -804 603 -792
rect 531 -856 541 -804
rect 593 -856 603 -804
rect 531 -868 603 -856
rect 531 -920 541 -868
rect 593 -920 603 -868
rect 531 -932 603 -920
rect 531 -984 541 -932
rect 593 -984 603 -932
rect 531 -996 603 -984
rect 531 -1048 541 -996
rect 593 -1048 603 -996
rect 531 -1060 603 -1048
rect 531 -1112 541 -1060
rect 593 -1112 603 -1060
rect 531 -1124 603 -1112
rect 531 -1176 541 -1124
rect 593 -1176 603 -1124
rect 531 -1188 603 -1176
rect 531 -1240 541 -1188
rect 593 -1240 603 -1188
rect 531 -1252 603 -1240
rect 531 -1304 541 -1252
rect 593 -1304 603 -1252
rect 531 -1316 603 -1304
rect 531 -1368 541 -1316
rect 593 -1368 603 -1316
rect 531 -1380 603 -1368
rect 531 -1432 541 -1380
rect 593 -1432 603 -1380
rect 531 -1444 603 -1432
rect 531 -1496 541 -1444
rect 593 -1496 603 -1444
rect 531 -1508 603 -1496
rect 531 -1560 541 -1508
rect 593 -1560 603 -1508
rect 531 -1572 603 -1560
rect 531 -1624 541 -1572
rect 593 -1624 603 -1572
rect 531 -1636 603 -1624
rect 531 -1688 541 -1636
rect 593 -1688 603 -1636
rect 531 -1700 603 -1688
rect 531 -1752 541 -1700
rect 593 -1752 603 -1700
rect 531 -1764 603 -1752
rect 661 -985 733 -963
rect 661 -1037 671 -985
rect 723 -1037 733 -985
rect 661 -1049 733 -1037
rect 661 -1101 671 -1049
rect 723 -1101 733 -1049
rect 661 -1113 733 -1101
rect 661 -1165 671 -1113
rect 723 -1165 733 -1113
rect 661 -1177 733 -1165
rect 661 -1229 671 -1177
rect 723 -1229 733 -1177
rect 661 -1241 733 -1229
rect 661 -1293 671 -1241
rect 723 -1293 733 -1241
rect 661 -1305 733 -1293
rect 661 -1357 671 -1305
rect 723 -1357 733 -1305
rect 661 -1369 733 -1357
rect 661 -1421 671 -1369
rect 723 -1421 733 -1369
rect 661 -1433 733 -1421
rect 661 -1485 671 -1433
rect 723 -1485 733 -1433
rect 661 -1497 733 -1485
rect 661 -1549 671 -1497
rect 723 -1549 733 -1497
rect 661 -1561 733 -1549
rect 661 -1613 671 -1561
rect 723 -1613 733 -1561
rect 661 -1625 733 -1613
rect 661 -1677 671 -1625
rect 723 -1677 733 -1625
rect 661 -1689 733 -1677
rect 661 -1741 671 -1689
rect 723 -1741 733 -1689
rect 661 -1763 733 -1741
rect 847 -985 919 -963
rect 847 -1037 857 -985
rect 909 -1037 919 -985
rect 847 -1049 919 -1037
rect 847 -1101 857 -1049
rect 909 -1101 919 -1049
rect 847 -1113 919 -1101
rect 847 -1165 857 -1113
rect 909 -1165 919 -1113
rect 847 -1177 919 -1165
rect 847 -1229 857 -1177
rect 909 -1229 919 -1177
rect 847 -1241 919 -1229
rect 847 -1293 857 -1241
rect 909 -1293 919 -1241
rect 847 -1305 919 -1293
rect 847 -1357 857 -1305
rect 909 -1357 919 -1305
rect 847 -1369 919 -1357
rect 847 -1421 857 -1369
rect 909 -1421 919 -1369
rect 847 -1433 919 -1421
rect 847 -1485 857 -1433
rect 909 -1485 919 -1433
rect 847 -1497 919 -1485
rect 847 -1549 857 -1497
rect 909 -1549 919 -1497
rect 847 -1561 919 -1549
rect 847 -1613 857 -1561
rect 909 -1613 919 -1561
rect 847 -1625 919 -1613
rect 847 -1677 857 -1625
rect 909 -1677 919 -1625
rect 847 -1689 919 -1677
rect 847 -1741 857 -1689
rect 909 -1741 919 -1689
rect 847 -1763 919 -1741
rect 531 -1816 541 -1764
rect 593 -1795 603 -1764
rect 593 -1816 764 -1795
rect 531 -1847 764 -1816
rect 816 -1847 1433 -1795
rect 29 -1955 39 -1903
rect 91 -1955 671 -1903
rect 723 -1955 733 -1903
rect 345 -2035 417 -2015
rect 345 -2087 355 -2035
rect 407 -2087 417 -2035
rect 345 -2099 417 -2087
rect 345 -2151 355 -2099
rect 407 -2151 417 -2099
rect 345 -2163 417 -2151
rect 345 -2215 355 -2163
rect 407 -2215 417 -2163
rect 345 -2227 417 -2215
rect 345 -2279 355 -2227
rect 407 -2279 417 -2227
rect 345 -2291 417 -2279
rect 345 -2343 355 -2291
rect 407 -2343 417 -2291
rect 345 -2355 417 -2343
rect 345 -2407 355 -2355
rect 407 -2407 417 -2355
rect 345 -2419 417 -2407
rect 345 -2471 355 -2419
rect 407 -2471 417 -2419
rect 345 -2483 417 -2471
rect 345 -2535 355 -2483
rect 407 -2535 417 -2483
rect 345 -2547 417 -2535
rect 345 -2599 355 -2547
rect 407 -2599 417 -2547
rect 345 -2611 417 -2599
rect 345 -2663 355 -2611
rect 407 -2663 417 -2611
rect 345 -2675 417 -2663
rect 345 -2727 355 -2675
rect 407 -2727 417 -2675
rect 345 -2739 417 -2727
rect 345 -2791 355 -2739
rect 407 -2791 417 -2739
rect 345 -2803 417 -2791
rect 345 -2855 355 -2803
rect 407 -2855 417 -2803
rect 345 -2867 417 -2855
rect 345 -2919 355 -2867
rect 407 -2919 417 -2867
rect 345 -2931 417 -2919
rect 345 -2983 355 -2931
rect 407 -2983 417 -2931
rect 345 -2995 417 -2983
rect 345 -3047 355 -2995
rect 407 -3047 417 -2995
rect 345 -3059 417 -3047
rect 345 -3111 355 -3059
rect 407 -3111 417 -3059
rect 29 -3129 101 -3115
rect 29 -3181 39 -3129
rect 91 -3181 101 -3129
rect 29 -3193 101 -3181
rect 29 -3245 39 -3193
rect 91 -3245 101 -3193
rect 29 -3257 101 -3245
rect 29 -3309 39 -3257
rect 91 -3309 101 -3257
rect 29 -3321 101 -3309
rect 29 -3373 39 -3321
rect 91 -3373 101 -3321
rect 29 -3385 101 -3373
rect 29 -3437 39 -3385
rect 91 -3437 101 -3385
rect 29 -3449 101 -3437
rect 29 -3501 39 -3449
rect 91 -3501 101 -3449
rect 29 -3515 101 -3501
rect 215 -3129 287 -3115
rect 215 -3181 225 -3129
rect 277 -3181 287 -3129
rect 215 -3193 287 -3181
rect 215 -3245 225 -3193
rect 277 -3245 287 -3193
rect 215 -3257 287 -3245
rect 215 -3309 225 -3257
rect 277 -3309 287 -3257
rect 215 -3321 287 -3309
rect 215 -3373 225 -3321
rect 277 -3373 287 -3321
rect 215 -3385 287 -3373
rect 215 -3437 225 -3385
rect 277 -3437 287 -3385
rect 215 -3449 287 -3437
rect 215 -3501 225 -3449
rect 277 -3501 287 -3449
rect 215 -3515 287 -3501
rect 345 -3123 417 -3111
rect 345 -3175 355 -3123
rect 407 -3175 417 -3123
rect 345 -3187 417 -3175
rect 345 -3239 355 -3187
rect 407 -3239 417 -3187
rect 345 -3251 417 -3239
rect 345 -3303 355 -3251
rect 407 -3303 417 -3251
rect 345 -3315 417 -3303
rect 345 -3367 355 -3315
rect 407 -3367 417 -3315
rect 345 -3379 417 -3367
rect 345 -3431 355 -3379
rect 407 -3431 417 -3379
rect 345 -3443 417 -3431
rect 345 -3495 355 -3443
rect 407 -3495 417 -3443
rect 345 -3515 417 -3495
rect 531 -2035 603 -2015
rect 531 -2087 541 -2035
rect 593 -2087 603 -2035
rect 754 -2045 764 -1993
rect 816 -2045 826 -1993
rect 531 -2099 603 -2087
rect 531 -2151 541 -2099
rect 593 -2151 603 -2099
rect 531 -2163 603 -2151
rect 531 -2215 541 -2163
rect 593 -2215 603 -2163
rect 531 -2227 603 -2215
rect 531 -2279 541 -2227
rect 593 -2279 603 -2227
rect 531 -2291 603 -2279
rect 531 -2343 541 -2291
rect 593 -2343 603 -2291
rect 531 -2355 603 -2343
rect 531 -2407 541 -2355
rect 593 -2407 603 -2355
rect 531 -2419 603 -2407
rect 531 -2471 541 -2419
rect 593 -2471 603 -2419
rect 531 -2483 603 -2471
rect 531 -2535 541 -2483
rect 593 -2535 603 -2483
rect 531 -2547 603 -2535
rect 531 -2599 541 -2547
rect 593 -2599 603 -2547
rect 531 -2611 603 -2599
rect 531 -2663 541 -2611
rect 593 -2663 603 -2611
rect 531 -2675 603 -2663
rect 531 -2727 541 -2675
rect 593 -2727 603 -2675
rect 531 -2739 603 -2727
rect 531 -2791 541 -2739
rect 593 -2791 603 -2739
rect 531 -2803 603 -2791
rect 531 -2855 541 -2803
rect 593 -2855 603 -2803
rect 531 -2867 603 -2855
rect 531 -2919 541 -2867
rect 593 -2919 603 -2867
rect 661 -2099 733 -2077
rect 661 -2151 671 -2099
rect 723 -2151 733 -2099
rect 661 -2163 733 -2151
rect 661 -2215 671 -2163
rect 723 -2215 733 -2163
rect 661 -2227 733 -2215
rect 661 -2279 671 -2227
rect 723 -2279 733 -2227
rect 661 -2291 733 -2279
rect 661 -2343 671 -2291
rect 723 -2343 733 -2291
rect 661 -2355 733 -2343
rect 661 -2407 671 -2355
rect 723 -2407 733 -2355
rect 661 -2419 733 -2407
rect 661 -2471 671 -2419
rect 723 -2471 733 -2419
rect 661 -2483 733 -2471
rect 661 -2535 671 -2483
rect 723 -2535 733 -2483
rect 817 -2451 851 -2443
rect 817 -2503 1433 -2451
rect 817 -2511 851 -2503
rect 661 -2547 733 -2535
rect 661 -2599 671 -2547
rect 723 -2599 733 -2547
rect 661 -2611 733 -2599
rect 661 -2663 671 -2611
rect 723 -2663 733 -2611
rect 661 -2675 733 -2663
rect 661 -2727 671 -2675
rect 723 -2727 733 -2675
rect 661 -2739 733 -2727
rect 661 -2791 671 -2739
rect 723 -2791 733 -2739
rect 661 -2803 733 -2791
rect 661 -2855 671 -2803
rect 723 -2855 733 -2803
rect 661 -2877 733 -2855
rect 531 -2931 603 -2919
rect 531 -2983 541 -2931
rect 593 -2983 603 -2931
rect 531 -2995 603 -2983
rect 531 -3047 541 -2995
rect 593 -3047 603 -2995
rect 531 -3059 603 -3047
rect 531 -3111 541 -3059
rect 593 -3111 603 -3059
rect 531 -3123 603 -3111
rect 531 -3175 541 -3123
rect 593 -3175 603 -3123
rect 531 -3187 603 -3175
rect 531 -3239 541 -3187
rect 593 -3239 603 -3187
rect 531 -3251 603 -3239
rect 531 -3303 541 -3251
rect 593 -3303 603 -3251
rect 531 -3315 603 -3303
rect 531 -3367 541 -3315
rect 593 -3367 603 -3315
rect 531 -3379 603 -3367
rect 531 -3431 541 -3379
rect 593 -3431 603 -3379
rect 531 -3443 603 -3431
rect 531 -3495 541 -3443
rect 593 -3495 603 -3443
rect 531 -3515 603 -3495
rect 129 -3587 1433 -3553
rect 215 -3701 225 -3649
rect 277 -3655 541 -3649
rect 297 -3689 335 -3655
rect 369 -3689 541 -3655
rect 277 -3701 541 -3689
rect 593 -3701 603 -3649
rect 237 -4036 395 -3701
rect -9799 -4067 1529 -4036
rect -9799 -4101 -9768 -4067
rect -9734 -4101 -9672 -4067
rect -9638 -4101 -9576 -4067
rect -9542 -4101 -9480 -4067
rect -9446 -4101 -9384 -4067
rect -9350 -4101 -9288 -4067
rect -9254 -4101 -9192 -4067
rect -9158 -4101 -9096 -4067
rect -9062 -4101 -9000 -4067
rect -8966 -4101 -8904 -4067
rect -8870 -4101 -8808 -4067
rect -8774 -4101 -8712 -4067
rect -8678 -4101 -8616 -4067
rect -8582 -4101 -8520 -4067
rect -8486 -4101 -8424 -4067
rect -8390 -4101 -8328 -4067
rect -8294 -4101 -8232 -4067
rect -8198 -4101 -8136 -4067
rect -8102 -4101 -8040 -4067
rect -8006 -4101 -7944 -4067
rect -7910 -4101 -7848 -4067
rect -7814 -4101 -7752 -4067
rect -7718 -4101 -7656 -4067
rect -7622 -4101 -7560 -4067
rect -7526 -4101 -7464 -4067
rect -7430 -4101 -7368 -4067
rect -7334 -4101 -7272 -4067
rect -7238 -4101 -7176 -4067
rect -7142 -4101 -7080 -4067
rect -7046 -4101 -6984 -4067
rect -6950 -4101 -6888 -4067
rect -6854 -4101 -6792 -4067
rect -6758 -4101 -6696 -4067
rect -6662 -4101 -6600 -4067
rect -6566 -4101 -6504 -4067
rect -6470 -4101 -6408 -4067
rect -6374 -4101 -6312 -4067
rect -6278 -4101 -6216 -4067
rect -6182 -4101 -6120 -4067
rect -6086 -4101 -6024 -4067
rect -5990 -4101 -5928 -4067
rect -5894 -4101 -5832 -4067
rect -5798 -4101 -5736 -4067
rect -5702 -4101 -5640 -4067
rect -5606 -4101 -5544 -4067
rect -5510 -4101 -5448 -4067
rect -5414 -4101 -5352 -4067
rect -5318 -4101 -5256 -4067
rect -5222 -4101 -5160 -4067
rect -5126 -4101 -5064 -4067
rect -5030 -4101 -4968 -4067
rect -4934 -4101 -4872 -4067
rect -4838 -4101 -4776 -4067
rect -4742 -4101 -4680 -4067
rect -4646 -4101 -4584 -4067
rect -4550 -4101 -4488 -4067
rect -4454 -4101 -4392 -4067
rect -4358 -4101 -4296 -4067
rect -4262 -4101 -4200 -4067
rect -4166 -4101 -4104 -4067
rect -4070 -4101 -4008 -4067
rect -3974 -4101 -3912 -4067
rect -3878 -4101 -3816 -4067
rect -3782 -4101 -3720 -4067
rect -3686 -4101 -3624 -4067
rect -3590 -4101 -3528 -4067
rect -3494 -4101 -3432 -4067
rect -3398 -4101 -3336 -4067
rect -3302 -4101 -3240 -4067
rect -3206 -4101 -3144 -4067
rect -3110 -4101 -3048 -4067
rect -3014 -4101 -2952 -4067
rect -2918 -4101 -2856 -4067
rect -2822 -4101 -2760 -4067
rect -2726 -4101 -2664 -4067
rect -2630 -4101 -2568 -4067
rect -2534 -4101 -2472 -4067
rect -2438 -4101 -2376 -4067
rect -2342 -4101 -2280 -4067
rect -2246 -4101 -2184 -4067
rect -2150 -4101 -2088 -4067
rect -2054 -4101 -1992 -4067
rect -1958 -4101 -1896 -4067
rect -1862 -4101 -1800 -4067
rect -1766 -4101 -1704 -4067
rect -1670 -4101 -1608 -4067
rect -1574 -4101 -1512 -4067
rect -1478 -4101 -1416 -4067
rect -1382 -4101 -1320 -4067
rect -1286 -4101 -1224 -4067
rect -1190 -4101 -1128 -4067
rect -1094 -4101 -1032 -4067
rect -998 -4101 -936 -4067
rect -902 -4101 -840 -4067
rect -806 -4101 -744 -4067
rect -710 -4101 -648 -4067
rect -614 -4101 -552 -4067
rect -518 -4101 -456 -4067
rect -422 -4101 -360 -4067
rect -326 -4101 -264 -4067
rect -230 -4101 -168 -4067
rect -134 -4101 -72 -4067
rect -38 -4101 24 -4067
rect 58 -4101 120 -4067
rect 154 -4101 216 -4067
rect 250 -4101 312 -4067
rect 346 -4101 408 -4067
rect 442 -4101 504 -4067
rect 538 -4101 600 -4067
rect 634 -4101 696 -4067
rect 730 -4101 792 -4067
rect 826 -4101 888 -4067
rect 922 -4101 984 -4067
rect 1018 -4101 1080 -4067
rect 1114 -4101 1176 -4067
rect 1210 -4101 1272 -4067
rect 1306 -4101 1368 -4067
rect 1402 -4101 1464 -4067
rect 1498 -4101 1529 -4067
rect -9799 -4132 1529 -4101
<< via1 >>
rect 448 455 500 507
rect 225 185 277 237
rect 225 121 277 173
rect -245 -19 -193 33
rect 132 11 184 63
rect 3963 874 4015 926
rect 3712 432 3721 459
rect 3721 432 3755 459
rect 3755 432 3764 459
rect 3712 407 3764 432
rect 3712 394 3764 395
rect 3712 360 3721 394
rect 3721 360 3755 394
rect 3755 360 3764 394
rect 3712 343 3764 360
rect 3712 322 3764 331
rect 3712 288 3721 322
rect 3721 288 3755 322
rect 3755 288 3764 322
rect 3712 279 3764 288
rect 3712 250 3764 267
rect 3712 216 3721 250
rect 3721 216 3755 250
rect 3755 216 3764 250
rect 3712 215 3764 216
rect 3712 178 3764 203
rect 3712 151 3721 178
rect 3721 151 3755 178
rect 3755 151 3764 178
rect 3963 439 4015 491
rect 3963 375 4015 427
rect 3963 311 4015 363
rect 3963 247 4015 299
rect 3963 183 4015 235
rect 3963 119 4015 171
rect 3870 12 3922 64
rect 3712 -97 3764 -45
rect -245 -175 -193 -123
rect 225 -201 277 -149
rect 857 -201 909 -149
rect 3870 -201 3922 -149
rect 132 -293 184 -241
rect 448 -293 500 -241
rect 39 -401 91 -349
rect 225 -401 277 -349
rect 355 -397 407 -345
rect 355 -461 407 -409
rect 355 -525 407 -473
rect 355 -589 407 -537
rect 355 -653 407 -601
rect 355 -717 407 -665
rect 355 -781 407 -729
rect 355 -845 407 -793
rect 355 -909 407 -857
rect 355 -973 407 -921
rect 355 -1037 407 -985
rect 355 -1101 407 -1049
rect 355 -1165 407 -1113
rect 355 -1229 407 -1177
rect 355 -1293 407 -1241
rect 355 -1357 407 -1305
rect 355 -1421 407 -1369
rect 355 -1485 407 -1433
rect 355 -1549 407 -1497
rect 355 -1613 407 -1561
rect 355 -1677 407 -1625
rect 355 -1741 407 -1689
rect 355 -1805 407 -1753
rect 541 -408 593 -356
rect 3963 -377 4015 -325
rect 541 -472 593 -420
rect 541 -536 593 -484
rect 541 -600 593 -548
rect 541 -664 593 -612
rect 541 -728 593 -676
rect 541 -792 593 -740
rect 541 -856 593 -804
rect 541 -920 593 -868
rect 541 -984 593 -932
rect 541 -1048 593 -996
rect 541 -1112 593 -1060
rect 541 -1176 593 -1124
rect 541 -1240 593 -1188
rect 541 -1304 593 -1252
rect 541 -1368 593 -1316
rect 541 -1432 593 -1380
rect 541 -1496 593 -1444
rect 541 -1560 593 -1508
rect 541 -1624 593 -1572
rect 541 -1688 593 -1636
rect 541 -1752 593 -1700
rect 671 -1037 723 -985
rect 671 -1101 723 -1049
rect 671 -1165 723 -1113
rect 671 -1229 723 -1177
rect 671 -1293 723 -1241
rect 671 -1357 723 -1305
rect 671 -1421 723 -1369
rect 671 -1485 723 -1433
rect 671 -1549 723 -1497
rect 671 -1613 723 -1561
rect 671 -1677 723 -1625
rect 671 -1741 723 -1689
rect 857 -1037 909 -985
rect 857 -1101 909 -1049
rect 857 -1165 909 -1113
rect 857 -1229 909 -1177
rect 857 -1293 909 -1241
rect 857 -1357 909 -1305
rect 857 -1421 909 -1369
rect 857 -1485 909 -1433
rect 857 -1549 909 -1497
rect 857 -1613 909 -1561
rect 857 -1677 909 -1625
rect 857 -1741 909 -1689
rect 541 -1816 593 -1764
rect 764 -1847 816 -1795
rect 39 -1955 91 -1903
rect 671 -1955 723 -1903
rect 355 -2087 407 -2035
rect 355 -2151 407 -2099
rect 355 -2215 407 -2163
rect 355 -2279 407 -2227
rect 355 -2343 407 -2291
rect 355 -2407 407 -2355
rect 355 -2471 407 -2419
rect 355 -2535 407 -2483
rect 355 -2599 407 -2547
rect 355 -2663 407 -2611
rect 355 -2727 407 -2675
rect 355 -2791 407 -2739
rect 355 -2855 407 -2803
rect 355 -2919 407 -2867
rect 355 -2983 407 -2931
rect 355 -3047 407 -2995
rect 355 -3111 407 -3059
rect 39 -3181 91 -3129
rect 39 -3245 91 -3193
rect 39 -3309 91 -3257
rect 39 -3373 91 -3321
rect 39 -3437 91 -3385
rect 39 -3501 91 -3449
rect 225 -3181 277 -3129
rect 225 -3245 277 -3193
rect 225 -3309 277 -3257
rect 225 -3373 277 -3321
rect 225 -3437 277 -3385
rect 225 -3501 277 -3449
rect 355 -3175 407 -3123
rect 355 -3239 407 -3187
rect 355 -3303 407 -3251
rect 355 -3367 407 -3315
rect 355 -3431 407 -3379
rect 355 -3495 407 -3443
rect 541 -2087 593 -2035
rect 764 -2045 816 -1993
rect 541 -2151 593 -2099
rect 541 -2215 593 -2163
rect 541 -2279 593 -2227
rect 541 -2343 593 -2291
rect 541 -2407 593 -2355
rect 541 -2471 593 -2419
rect 541 -2535 593 -2483
rect 541 -2599 593 -2547
rect 541 -2663 593 -2611
rect 541 -2727 593 -2675
rect 541 -2791 593 -2739
rect 541 -2855 593 -2803
rect 541 -2919 593 -2867
rect 671 -2151 723 -2099
rect 671 -2215 723 -2163
rect 671 -2279 723 -2227
rect 671 -2343 723 -2291
rect 671 -2407 723 -2355
rect 671 -2471 723 -2419
rect 671 -2535 723 -2483
rect 671 -2599 723 -2547
rect 671 -2663 723 -2611
rect 671 -2727 723 -2675
rect 671 -2791 723 -2739
rect 671 -2855 723 -2803
rect 541 -2983 593 -2931
rect 541 -3047 593 -2995
rect 541 -3111 593 -3059
rect 541 -3175 593 -3123
rect 541 -3239 593 -3187
rect 541 -3303 593 -3251
rect 541 -3367 593 -3315
rect 541 -3431 593 -3379
rect 541 -3495 593 -3443
rect 225 -3655 277 -3649
rect 225 -3689 263 -3655
rect 263 -3689 277 -3655
rect 225 -3701 277 -3689
rect 541 -3701 593 -3649
<< metal2 >>
rect 3963 926 4015 936
rect 448 507 500 517
rect 3963 491 4015 874
rect 225 237 277 264
rect 225 173 277 185
rect -271 35 -167 69
rect -271 -21 -247 35
rect -191 -21 -167 35
rect -271 -55 -167 -21
rect 132 63 184 73
rect 132 -77 184 11
rect 128 -87 184 -77
rect -271 -121 -167 -87
rect -271 -177 -247 -121
rect -191 -177 -167 -121
rect 128 -153 184 -143
rect -271 -211 -167 -177
rect 132 -241 184 -153
rect 132 -303 184 -293
rect 225 -149 277 121
rect 39 -349 91 -315
rect 39 -1903 91 -401
rect 225 -349 277 -201
rect 448 -241 500 455
rect 3712 459 3764 481
rect 3712 395 3764 407
rect 3712 331 3764 343
rect 3712 267 3764 279
rect 3712 203 3764 215
rect 3712 -45 3764 151
rect 3963 427 4015 439
rect 3963 363 4015 375
rect 3963 299 4015 311
rect 3963 235 4015 247
rect 3963 171 4015 183
rect 3712 -107 3764 -97
rect 3870 64 3922 74
rect 448 -303 500 -293
rect 857 -149 909 -139
rect 225 -435 277 -401
rect 355 -345 407 -315
rect 355 -409 407 -397
rect 39 -2543 91 -1955
rect 35 -2553 91 -2543
rect 35 -2713 91 -2609
rect 35 -2779 91 -2769
rect 39 -3129 91 -2779
rect 355 -473 407 -461
rect 355 -537 407 -525
rect 355 -601 407 -589
rect 355 -665 407 -653
rect 355 -729 407 -717
rect 355 -793 407 -781
rect 355 -857 407 -845
rect 355 -921 407 -909
rect 355 -985 407 -973
rect 355 -1049 407 -1037
rect 355 -1113 407 -1101
rect 355 -1177 407 -1165
rect 355 -1241 407 -1229
rect 355 -1305 407 -1293
rect 355 -1369 407 -1357
rect 355 -1433 407 -1421
rect 355 -1497 407 -1485
rect 355 -1561 407 -1549
rect 355 -1625 407 -1613
rect 355 -1689 407 -1677
rect 355 -1753 407 -1741
rect 355 -2035 407 -1805
rect 541 -356 593 -315
rect 541 -420 593 -408
rect 541 -484 593 -472
rect 541 -548 593 -536
rect 541 -612 593 -600
rect 541 -676 593 -664
rect 541 -740 593 -728
rect 541 -804 593 -792
rect 541 -868 593 -856
rect 541 -932 593 -920
rect 541 -996 593 -984
rect 541 -1060 593 -1048
rect 541 -1124 593 -1112
rect 541 -1188 593 -1176
rect 541 -1252 593 -1240
rect 541 -1316 593 -1304
rect 541 -1380 593 -1368
rect 541 -1444 593 -1432
rect 541 -1508 593 -1496
rect 541 -1572 593 -1560
rect 541 -1636 593 -1624
rect 541 -1700 593 -1688
rect 541 -1764 593 -1752
rect 541 -1857 593 -1816
rect 671 -985 723 -953
rect 671 -1049 723 -1037
rect 671 -1113 723 -1101
rect 671 -1177 723 -1165
rect 671 -1241 723 -1229
rect 671 -1305 723 -1293
rect 671 -1369 723 -1357
rect 671 -1433 723 -1421
rect 671 -1497 723 -1485
rect 671 -1561 723 -1549
rect 671 -1625 723 -1613
rect 671 -1689 723 -1677
rect 671 -1903 723 -1741
rect 857 -985 909 -201
rect 3870 -149 3922 12
rect 3870 -211 3922 -201
rect 3963 -325 4015 119
rect 3963 -387 4015 -377
rect 857 -1049 909 -1037
rect 857 -1113 909 -1101
rect 857 -1177 909 -1165
rect 857 -1241 909 -1229
rect 857 -1305 909 -1293
rect 857 -1369 909 -1357
rect 857 -1433 909 -1421
rect 857 -1497 909 -1485
rect 857 -1561 909 -1549
rect 857 -1625 909 -1613
rect 857 -1689 909 -1677
rect 857 -1773 909 -1741
rect 355 -2099 407 -2087
rect 355 -2163 407 -2151
rect 355 -2227 407 -2215
rect 355 -2291 407 -2279
rect 355 -2355 407 -2343
rect 355 -2419 407 -2407
rect 355 -2483 407 -2471
rect 355 -2547 407 -2535
rect 355 -2611 407 -2599
rect 355 -2675 407 -2663
rect 355 -2739 407 -2727
rect 355 -2803 407 -2791
rect 355 -2867 407 -2855
rect 355 -2931 407 -2919
rect 355 -2995 407 -2983
rect 355 -3059 407 -3047
rect 39 -3193 91 -3181
rect 39 -3257 91 -3245
rect 39 -3321 91 -3309
rect 39 -3385 91 -3373
rect 39 -3449 91 -3437
rect 39 -3525 91 -3501
rect 225 -3129 277 -3105
rect 225 -3193 277 -3181
rect 225 -3257 277 -3245
rect 225 -3321 277 -3309
rect 225 -3385 277 -3373
rect 225 -3449 277 -3437
rect 225 -3649 277 -3501
rect 355 -3123 407 -3111
rect 355 -3187 407 -3175
rect 355 -3251 407 -3239
rect 355 -3315 407 -3303
rect 355 -3379 407 -3367
rect 355 -3443 407 -3431
rect 355 -3525 407 -3495
rect 541 -2035 593 -2005
rect 541 -2099 593 -2087
rect 541 -2163 593 -2151
rect 541 -2227 593 -2215
rect 541 -2291 593 -2279
rect 541 -2355 593 -2343
rect 541 -2419 593 -2407
rect 541 -2483 593 -2471
rect 541 -2547 593 -2535
rect 541 -2611 593 -2599
rect 541 -2675 593 -2663
rect 541 -2739 593 -2727
rect 541 -2803 593 -2791
rect 541 -2867 593 -2855
rect 671 -2099 723 -1955
rect 764 -1795 816 -1785
rect 764 -1993 816 -1847
rect 764 -2055 816 -2045
rect 671 -2163 723 -2151
rect 671 -2227 723 -2215
rect 671 -2291 723 -2279
rect 671 -2355 723 -2343
rect 671 -2419 723 -2407
rect 671 -2483 723 -2471
rect 671 -2547 723 -2535
rect 671 -2611 723 -2599
rect 671 -2675 723 -2663
rect 671 -2739 723 -2727
rect 671 -2803 723 -2791
rect 671 -2887 723 -2855
rect 541 -2931 593 -2919
rect 541 -2995 593 -2983
rect 541 -3059 593 -3047
rect 541 -3123 593 -3111
rect 541 -3187 593 -3175
rect 541 -3251 593 -3239
rect 541 -3315 593 -3303
rect 541 -3379 593 -3367
rect 541 -3443 593 -3431
rect 225 -3711 277 -3701
rect 541 -3649 593 -3495
rect 541 -3711 593 -3701
<< via2 >>
rect -247 33 -191 35
rect -247 -19 -245 33
rect -245 -19 -193 33
rect -193 -19 -191 33
rect -247 -21 -191 -19
rect -247 -123 -191 -121
rect -247 -175 -245 -123
rect -245 -175 -193 -123
rect -193 -175 -191 -123
rect -247 -177 -191 -175
rect 128 -143 184 -87
rect 35 -2609 91 -2553
rect 35 -2769 91 -2713
<< metal3 >>
rect -281 39 -157 64
rect -281 -25 -251 39
rect -187 -25 -157 39
rect -281 -117 -157 -25
rect -281 -181 -251 -117
rect -187 -181 -157 -117
rect 118 -87 1433 -82
rect 118 -143 128 -87
rect 184 -143 1433 -87
rect 118 -148 1433 -143
rect -281 -206 -157 -181
rect 25 -2553 101 -2548
rect 25 -2609 35 -2553
rect 91 -2609 101 -2553
rect -505 -2629 101 -2609
rect -505 -2693 -467 -2629
rect -403 -2693 101 -2629
rect -505 -2713 101 -2693
rect 25 -2769 35 -2713
rect 91 -2769 101 -2713
rect 25 -2774 101 -2769
<< via3 >>
rect -251 35 -187 39
rect -251 -21 -247 35
rect -247 -21 -191 35
rect -191 -21 -187 35
rect -251 -25 -187 -21
rect -251 -121 -187 -117
rect -251 -177 -247 -121
rect -247 -177 -191 -121
rect -191 -177 -187 -121
rect -251 -181 -187 -177
rect -467 -2693 -403 -2629
<< metal4 >>
rect -9543 1523 -9335 1627
rect -9543 215 -9439 1523
rect -375 843 -167 947
rect -9543 111 -9229 215
rect -9543 -1197 -9439 111
rect -271 60 -167 843
rect -272 39 -166 60
rect -272 -25 -251 39
rect -187 -25 -166 39
rect -272 -117 -166 -25
rect -272 -181 -251 -117
rect -187 -181 -166 -117
rect -272 -202 -166 -181
rect -271 -465 -167 -202
rect -375 -569 -167 -465
rect -9543 -1301 -9224 -1197
rect -9543 -2609 -9439 -1301
rect -271 -1877 -167 -569
rect -375 -1981 -167 -1877
rect -9543 -2713 -9231 -2609
rect -496 -2629 -374 -2608
rect -496 -2693 -467 -2629
rect -403 -2693 -374 -2629
rect -496 -2714 -374 -2693
rect -271 -3289 -167 -1981
rect -375 -3393 -167 -3289
use sky130_fd_pr__nfet_01v8_J4Y94J  sky130_fd_pr__nfet_01v8_J4Y94J_0
timestamp 1750100919
transform 1 0 790 0 1 -2446
box -201 -569 201 569
use sky130_fd_pr__cap_mim_m3_1_9XU9T9  XC1
timestamp 1750100919
transform 0 1 -4855 1 0 -1077
box -2704 -4480 2704 4480
use sky130_fd_pr__pfet_01v8_27QFPY  XM1
timestamp 1750100919
transform 1 0 158 0 1 144
box -211 -259 211 259
use sky130_fd_pr__pfet_01v8_MGASDN  XM2
timestamp 1750100919
transform 1 0 3580 0 1 469
box -211 -584 211 584
use sky130_fd_pr__pfet_01v8_LGMQDL  XM3
timestamp 1750100919
transform 1 0 3896 0 1 269
box -211 -384 211 384
use sky130_fd_pr__nfet_01v8_CQKS6Z  XM4
timestamp 1750100919
transform 1 0 158 0 1 -344
box -201 -219 201 219
use sky130_fd_pr__nfet_01v8_46WN23  XM5
timestamp 1750100919
transform 1 0 158 0 1 -3346
box -201 -369 201 369
use sky130_fd_pr__nfet_01v8_J47Z3J  XM6
timestamp 1750100919
transform 1 0 790 0 1 -1394
box -201 -569 201 569
use sky130_fd_pr__nfet_01v8_D4Y996  XM8
timestamp 1750100919
transform 1 0 474 0 1 -1044
box -201 -919 201 919
use sky130_fd_pr__nfet_01v8_D47ZC5  XM9
timestamp 1750100919
transform 1 0 474 0 1 -2796
box -201 -919 201 919
<< labels >>
flabel metal1 s 1464 1913 1498 1947 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 1464 -4101 1498 -4067 0 FreeSans 500 0 0 0 VSS
port 2 nsew
flabel metal1 s 1390 -2494 1424 -2460 0 FreeSans 500 0 0 0 IN
port 3 nsew
flabel metal1 s 1389 -1839 1423 -1805 0 FreeSans 500 0 0 0 VGS
port 4 nsew
flabel metal1 s 1399 -3587 1433 -3553 0 FreeSans 500 0 0 0 CK
port 5 nsew
flabel metal3 s 1378 -139 1412 -105 0 FreeSans 500 0 0 0 CKB
port 6 nsew
<< end >>
