magic
tech sky130A
magscale 1 2
timestamp 1746183165
<< pwell >>
rect -246 -1415 246 1415
<< nmos >>
rect -50 1105 50 1205
rect -50 895 50 995
rect -50 685 50 785
rect -50 475 50 575
rect -50 265 50 365
rect -50 55 50 155
rect -50 -155 50 -55
rect -50 -365 50 -265
rect -50 -575 50 -475
rect -50 -785 50 -685
rect -50 -995 50 -895
rect -50 -1205 50 -1105
<< ndiff >>
rect -108 1193 -50 1205
rect -108 1117 -96 1193
rect -62 1117 -50 1193
rect -108 1105 -50 1117
rect 50 1193 108 1205
rect 50 1117 62 1193
rect 96 1117 108 1193
rect 50 1105 108 1117
rect -108 983 -50 995
rect -108 907 -96 983
rect -62 907 -50 983
rect -108 895 -50 907
rect 50 983 108 995
rect 50 907 62 983
rect 96 907 108 983
rect 50 895 108 907
rect -108 773 -50 785
rect -108 697 -96 773
rect -62 697 -50 773
rect -108 685 -50 697
rect 50 773 108 785
rect 50 697 62 773
rect 96 697 108 773
rect 50 685 108 697
rect -108 563 -50 575
rect -108 487 -96 563
rect -62 487 -50 563
rect -108 475 -50 487
rect 50 563 108 575
rect 50 487 62 563
rect 96 487 108 563
rect 50 475 108 487
rect -108 353 -50 365
rect -108 277 -96 353
rect -62 277 -50 353
rect -108 265 -50 277
rect 50 353 108 365
rect 50 277 62 353
rect 96 277 108 353
rect 50 265 108 277
rect -108 143 -50 155
rect -108 67 -96 143
rect -62 67 -50 143
rect -108 55 -50 67
rect 50 143 108 155
rect 50 67 62 143
rect 96 67 108 143
rect 50 55 108 67
rect -108 -67 -50 -55
rect -108 -143 -96 -67
rect -62 -143 -50 -67
rect -108 -155 -50 -143
rect 50 -67 108 -55
rect 50 -143 62 -67
rect 96 -143 108 -67
rect 50 -155 108 -143
rect -108 -277 -50 -265
rect -108 -353 -96 -277
rect -62 -353 -50 -277
rect -108 -365 -50 -353
rect 50 -277 108 -265
rect 50 -353 62 -277
rect 96 -353 108 -277
rect 50 -365 108 -353
rect -108 -487 -50 -475
rect -108 -563 -96 -487
rect -62 -563 -50 -487
rect -108 -575 -50 -563
rect 50 -487 108 -475
rect 50 -563 62 -487
rect 96 -563 108 -487
rect 50 -575 108 -563
rect -108 -697 -50 -685
rect -108 -773 -96 -697
rect -62 -773 -50 -697
rect -108 -785 -50 -773
rect 50 -697 108 -685
rect 50 -773 62 -697
rect 96 -773 108 -697
rect 50 -785 108 -773
rect -108 -907 -50 -895
rect -108 -983 -96 -907
rect -62 -983 -50 -907
rect -108 -995 -50 -983
rect 50 -907 108 -895
rect 50 -983 62 -907
rect 96 -983 108 -907
rect 50 -995 108 -983
rect -108 -1117 -50 -1105
rect -108 -1193 -96 -1117
rect -62 -1193 -50 -1117
rect -108 -1205 -50 -1193
rect 50 -1117 108 -1105
rect 50 -1193 62 -1117
rect 96 -1193 108 -1117
rect 50 -1205 108 -1193
<< ndiffc >>
rect -96 1117 -62 1193
rect 62 1117 96 1193
rect -96 907 -62 983
rect 62 907 96 983
rect -96 697 -62 773
rect 62 697 96 773
rect -96 487 -62 563
rect 62 487 96 563
rect -96 277 -62 353
rect 62 277 96 353
rect -96 67 -62 143
rect 62 67 96 143
rect -96 -143 -62 -67
rect 62 -143 96 -67
rect -96 -353 -62 -277
rect 62 -353 96 -277
rect -96 -563 -62 -487
rect 62 -563 96 -487
rect -96 -773 -62 -697
rect 62 -773 96 -697
rect -96 -983 -62 -907
rect 62 -983 96 -907
rect -96 -1193 -62 -1117
rect 62 -1193 96 -1117
<< psubdiff >>
rect -210 1345 -114 1379
rect 114 1345 210 1379
rect -210 1283 -176 1345
rect 176 1283 210 1345
rect -210 -1345 -176 -1283
rect 176 -1345 210 -1283
rect -210 -1379 -114 -1345
rect 114 -1379 210 -1345
<< psubdiffcont >>
rect -114 1345 114 1379
rect -210 -1283 -176 1283
rect 176 -1283 210 1283
rect -114 -1379 114 -1345
<< poly >>
rect -50 1277 50 1293
rect -50 1243 -34 1277
rect 34 1243 50 1277
rect -50 1205 50 1243
rect -50 1067 50 1105
rect -50 1033 -34 1067
rect 34 1033 50 1067
rect -50 995 50 1033
rect -50 857 50 895
rect -50 823 -34 857
rect 34 823 50 857
rect -50 785 50 823
rect -50 647 50 685
rect -50 613 -34 647
rect 34 613 50 647
rect -50 575 50 613
rect -50 437 50 475
rect -50 403 -34 437
rect 34 403 50 437
rect -50 365 50 403
rect -50 227 50 265
rect -50 193 -34 227
rect 34 193 50 227
rect -50 155 50 193
rect -50 17 50 55
rect -50 -17 -34 17
rect 34 -17 50 17
rect -50 -55 50 -17
rect -50 -193 50 -155
rect -50 -227 -34 -193
rect 34 -227 50 -193
rect -50 -265 50 -227
rect -50 -403 50 -365
rect -50 -437 -34 -403
rect 34 -437 50 -403
rect -50 -475 50 -437
rect -50 -613 50 -575
rect -50 -647 -34 -613
rect 34 -647 50 -613
rect -50 -685 50 -647
rect -50 -823 50 -785
rect -50 -857 -34 -823
rect 34 -857 50 -823
rect -50 -895 50 -857
rect -50 -1033 50 -995
rect -50 -1067 -34 -1033
rect 34 -1067 50 -1033
rect -50 -1105 50 -1067
rect -50 -1243 50 -1205
rect -50 -1277 -34 -1243
rect 34 -1277 50 -1243
rect -50 -1293 50 -1277
<< polycont >>
rect -34 1243 34 1277
rect -34 1033 34 1067
rect -34 823 34 857
rect -34 613 34 647
rect -34 403 34 437
rect -34 193 34 227
rect -34 -17 34 17
rect -34 -227 34 -193
rect -34 -437 34 -403
rect -34 -647 34 -613
rect -34 -857 34 -823
rect -34 -1067 34 -1033
rect -34 -1277 34 -1243
<< locali >>
rect -210 1345 -114 1379
rect 114 1345 210 1379
rect -210 1283 -176 1345
rect 176 1283 210 1345
rect -50 1243 -34 1277
rect 34 1243 50 1277
rect -96 1193 -62 1209
rect -96 1101 -62 1117
rect 62 1193 96 1209
rect 62 1101 96 1117
rect -50 1033 -34 1067
rect 34 1033 50 1067
rect -96 983 -62 999
rect -96 891 -62 907
rect 62 983 96 999
rect 62 891 96 907
rect -50 823 -34 857
rect 34 823 50 857
rect -96 773 -62 789
rect -96 681 -62 697
rect 62 773 96 789
rect 62 681 96 697
rect -50 613 -34 647
rect 34 613 50 647
rect -96 563 -62 579
rect -96 471 -62 487
rect 62 563 96 579
rect 62 471 96 487
rect -50 403 -34 437
rect 34 403 50 437
rect -96 353 -62 369
rect -96 261 -62 277
rect 62 353 96 369
rect 62 261 96 277
rect -50 193 -34 227
rect 34 193 50 227
rect -96 143 -62 159
rect -96 51 -62 67
rect 62 143 96 159
rect 62 51 96 67
rect -50 -17 -34 17
rect 34 -17 50 17
rect -96 -67 -62 -51
rect -96 -159 -62 -143
rect 62 -67 96 -51
rect 62 -159 96 -143
rect -50 -227 -34 -193
rect 34 -227 50 -193
rect -96 -277 -62 -261
rect -96 -369 -62 -353
rect 62 -277 96 -261
rect 62 -369 96 -353
rect -50 -437 -34 -403
rect 34 -437 50 -403
rect -96 -487 -62 -471
rect -96 -579 -62 -563
rect 62 -487 96 -471
rect 62 -579 96 -563
rect -50 -647 -34 -613
rect 34 -647 50 -613
rect -96 -697 -62 -681
rect -96 -789 -62 -773
rect 62 -697 96 -681
rect 62 -789 96 -773
rect -50 -857 -34 -823
rect 34 -857 50 -823
rect -96 -907 -62 -891
rect -96 -999 -62 -983
rect 62 -907 96 -891
rect 62 -999 96 -983
rect -50 -1067 -34 -1033
rect 34 -1067 50 -1033
rect -96 -1117 -62 -1101
rect -96 -1209 -62 -1193
rect 62 -1117 96 -1101
rect 62 -1209 96 -1193
rect -50 -1277 -34 -1243
rect 34 -1277 50 -1243
rect -210 -1345 -176 -1283
rect 176 -1345 210 -1283
rect -210 -1379 -114 -1345
rect 114 -1379 210 -1345
<< viali >>
rect -34 1243 34 1277
rect -96 1117 -62 1193
rect 62 1117 96 1193
rect -34 1033 34 1067
rect -96 907 -62 983
rect 62 907 96 983
rect -34 823 34 857
rect -96 697 -62 773
rect 62 697 96 773
rect -34 613 34 647
rect -96 487 -62 563
rect 62 487 96 563
rect -34 403 34 437
rect -96 277 -62 353
rect 62 277 96 353
rect -34 193 34 227
rect -96 67 -62 143
rect 62 67 96 143
rect -34 -17 34 17
rect -96 -143 -62 -67
rect 62 -143 96 -67
rect -34 -227 34 -193
rect -96 -353 -62 -277
rect 62 -353 96 -277
rect -34 -437 34 -403
rect -96 -563 -62 -487
rect 62 -563 96 -487
rect -34 -647 34 -613
rect -96 -773 -62 -697
rect 62 -773 96 -697
rect -34 -857 34 -823
rect -96 -983 -62 -907
rect 62 -983 96 -907
rect -34 -1067 34 -1033
rect -96 -1193 -62 -1117
rect 62 -1193 96 -1117
rect -34 -1277 34 -1243
<< metal1 >>
rect -46 1277 46 1283
rect -46 1243 -34 1277
rect 34 1243 46 1277
rect -46 1237 46 1243
rect -102 1193 -56 1205
rect -102 1117 -96 1193
rect -62 1117 -56 1193
rect -102 1105 -56 1117
rect 56 1193 102 1205
rect 56 1117 62 1193
rect 96 1117 102 1193
rect 56 1105 102 1117
rect -46 1067 46 1073
rect -46 1033 -34 1067
rect 34 1033 46 1067
rect -46 1027 46 1033
rect -102 983 -56 995
rect -102 907 -96 983
rect -62 907 -56 983
rect -102 895 -56 907
rect 56 983 102 995
rect 56 907 62 983
rect 96 907 102 983
rect 56 895 102 907
rect -46 857 46 863
rect -46 823 -34 857
rect 34 823 46 857
rect -46 817 46 823
rect -102 773 -56 785
rect -102 697 -96 773
rect -62 697 -56 773
rect -102 685 -56 697
rect 56 773 102 785
rect 56 697 62 773
rect 96 697 102 773
rect 56 685 102 697
rect -46 647 46 653
rect -46 613 -34 647
rect 34 613 46 647
rect -46 607 46 613
rect -102 563 -56 575
rect -102 487 -96 563
rect -62 487 -56 563
rect -102 475 -56 487
rect 56 563 102 575
rect 56 487 62 563
rect 96 487 102 563
rect 56 475 102 487
rect -46 437 46 443
rect -46 403 -34 437
rect 34 403 46 437
rect -46 397 46 403
rect -102 353 -56 365
rect -102 277 -96 353
rect -62 277 -56 353
rect -102 265 -56 277
rect 56 353 102 365
rect 56 277 62 353
rect 96 277 102 353
rect 56 265 102 277
rect -46 227 46 233
rect -46 193 -34 227
rect 34 193 46 227
rect -46 187 46 193
rect -102 143 -56 155
rect -102 67 -96 143
rect -62 67 -56 143
rect -102 55 -56 67
rect 56 143 102 155
rect 56 67 62 143
rect 96 67 102 143
rect 56 55 102 67
rect -46 17 46 23
rect -46 -17 -34 17
rect 34 -17 46 17
rect -46 -23 46 -17
rect -102 -67 -56 -55
rect -102 -143 -96 -67
rect -62 -143 -56 -67
rect -102 -155 -56 -143
rect 56 -67 102 -55
rect 56 -143 62 -67
rect 96 -143 102 -67
rect 56 -155 102 -143
rect -46 -193 46 -187
rect -46 -227 -34 -193
rect 34 -227 46 -193
rect -46 -233 46 -227
rect -102 -277 -56 -265
rect -102 -353 -96 -277
rect -62 -353 -56 -277
rect -102 -365 -56 -353
rect 56 -277 102 -265
rect 56 -353 62 -277
rect 96 -353 102 -277
rect 56 -365 102 -353
rect -46 -403 46 -397
rect -46 -437 -34 -403
rect 34 -437 46 -403
rect -46 -443 46 -437
rect -102 -487 -56 -475
rect -102 -563 -96 -487
rect -62 -563 -56 -487
rect -102 -575 -56 -563
rect 56 -487 102 -475
rect 56 -563 62 -487
rect 96 -563 102 -487
rect 56 -575 102 -563
rect -46 -613 46 -607
rect -46 -647 -34 -613
rect 34 -647 46 -613
rect -46 -653 46 -647
rect -102 -697 -56 -685
rect -102 -773 -96 -697
rect -62 -773 -56 -697
rect -102 -785 -56 -773
rect 56 -697 102 -685
rect 56 -773 62 -697
rect 96 -773 102 -697
rect 56 -785 102 -773
rect -46 -823 46 -817
rect -46 -857 -34 -823
rect 34 -857 46 -823
rect -46 -863 46 -857
rect -102 -907 -56 -895
rect -102 -983 -96 -907
rect -62 -983 -56 -907
rect -102 -995 -56 -983
rect 56 -907 102 -895
rect 56 -983 62 -907
rect 96 -983 102 -907
rect 56 -995 102 -983
rect -46 -1033 46 -1027
rect -46 -1067 -34 -1033
rect 34 -1067 46 -1033
rect -46 -1073 46 -1067
rect -102 -1117 -56 -1105
rect -102 -1193 -96 -1117
rect -62 -1193 -56 -1117
rect -102 -1205 -56 -1193
rect 56 -1117 102 -1105
rect 56 -1193 62 -1117
rect 96 -1193 102 -1117
rect 56 -1205 102 -1193
rect -46 -1243 46 -1237
rect -46 -1277 -34 -1243
rect 34 -1277 46 -1243
rect -46 -1283 46 -1277
<< properties >>
string FIXED_BBOX -193 -1362 193 1362
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 0.5 m 12 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
