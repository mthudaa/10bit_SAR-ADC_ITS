magic
tech sky130A
magscale 1 2
timestamp 1750100919
<< locali >>
rect 238 1527 264 1561
rect 298 1527 336 1561
rect 370 1527 408 1561
rect 442 1527 480 1561
rect 514 1527 552 1561
rect 586 1527 624 1561
rect 658 1527 696 1561
rect 730 1527 768 1561
rect 802 1527 840 1561
rect 874 1527 912 1561
rect 946 1527 984 1561
rect 1018 1527 1056 1561
rect 1090 1527 1128 1561
rect 1162 1527 1200 1561
rect 1234 1527 1272 1561
rect 1306 1527 1344 1561
rect 1378 1527 1416 1561
rect 1450 1527 1488 1561
rect 1522 1527 1560 1561
rect 1594 1527 1632 1561
rect 1666 1527 1704 1561
rect 1738 1527 1776 1561
rect 1810 1527 1848 1561
rect 1882 1527 1920 1561
rect 1954 1527 1992 1561
rect 2026 1527 2064 1561
rect 2098 1527 2136 1561
rect 2170 1527 2208 1561
rect 2242 1527 2280 1561
rect 2314 1527 2352 1561
rect 2386 1527 2424 1561
rect 2458 1527 2496 1561
rect 2530 1527 2568 1561
rect 2602 1527 2640 1561
rect 2674 1527 2712 1561
rect 2746 1527 2784 1561
rect 2818 1527 2856 1561
rect 2890 1527 2928 1561
rect 2962 1527 3000 1561
rect 3034 1527 3072 1561
rect 3106 1527 3144 1561
rect 3178 1527 3216 1561
rect 3250 1527 3288 1561
rect 3322 1527 3360 1561
rect 3394 1527 3432 1561
rect 3466 1527 3504 1561
rect 3538 1527 3576 1561
rect 3610 1527 3648 1561
rect 3682 1527 3708 1561
rect 238 -123 256 -89
rect 290 -123 328 -89
rect 362 -123 400 -89
rect 434 -123 472 -89
rect 506 -123 544 -89
rect 578 -123 616 -89
rect 650 -123 688 -89
rect 722 -123 760 -89
rect 794 -123 832 -89
rect 866 -123 904 -89
rect 938 -123 976 -89
rect 1010 -123 1048 -89
rect 1082 -123 1120 -89
rect 1154 -123 1192 -89
rect 1226 -123 1264 -89
rect 1298 -123 1336 -89
rect 1370 -123 1408 -89
rect 1442 -123 1480 -89
rect 1514 -123 1552 -89
rect 1586 -123 1624 -89
rect 1658 -123 1696 -89
rect 1730 -123 1768 -89
rect 1802 -123 1840 -89
rect 1874 -123 1912 -89
rect 1946 -123 1964 -89
<< viali >>
rect 264 1527 298 1561
rect 336 1527 370 1561
rect 408 1527 442 1561
rect 480 1527 514 1561
rect 552 1527 586 1561
rect 624 1527 658 1561
rect 696 1527 730 1561
rect 768 1527 802 1561
rect 840 1527 874 1561
rect 912 1527 946 1561
rect 984 1527 1018 1561
rect 1056 1527 1090 1561
rect 1128 1527 1162 1561
rect 1200 1527 1234 1561
rect 1272 1527 1306 1561
rect 1344 1527 1378 1561
rect 1416 1527 1450 1561
rect 1488 1527 1522 1561
rect 1560 1527 1594 1561
rect 1632 1527 1666 1561
rect 1704 1527 1738 1561
rect 1776 1527 1810 1561
rect 1848 1527 1882 1561
rect 1920 1527 1954 1561
rect 1992 1527 2026 1561
rect 2064 1527 2098 1561
rect 2136 1527 2170 1561
rect 2208 1527 2242 1561
rect 2280 1527 2314 1561
rect 2352 1527 2386 1561
rect 2424 1527 2458 1561
rect 2496 1527 2530 1561
rect 2568 1527 2602 1561
rect 2640 1527 2674 1561
rect 2712 1527 2746 1561
rect 2784 1527 2818 1561
rect 2856 1527 2890 1561
rect 2928 1527 2962 1561
rect 3000 1527 3034 1561
rect 3072 1527 3106 1561
rect 3144 1527 3178 1561
rect 3216 1527 3250 1561
rect 3288 1527 3322 1561
rect 3360 1527 3394 1561
rect 3432 1527 3466 1561
rect 3504 1527 3538 1561
rect 3576 1527 3610 1561
rect 3648 1527 3682 1561
rect 256 -123 290 -89
rect 328 -123 362 -89
rect 400 -123 434 -89
rect 472 -123 506 -89
rect 544 -123 578 -89
rect 616 -123 650 -89
rect 688 -123 722 -89
rect 760 -123 794 -89
rect 832 -123 866 -89
rect 904 -123 938 -89
rect 976 -123 1010 -89
rect 1048 -123 1082 -89
rect 1120 -123 1154 -89
rect 1192 -123 1226 -89
rect 1264 -123 1298 -89
rect 1336 -123 1370 -89
rect 1408 -123 1442 -89
rect 1480 -123 1514 -89
rect 1552 -123 1586 -89
rect 1624 -123 1658 -89
rect 1696 -123 1730 -89
rect 1768 -123 1802 -89
rect 1840 -123 1874 -89
rect 1912 -123 1946 -89
<< metal1 >>
rect 106 1561 3840 1597
rect 106 1527 264 1561
rect 298 1527 336 1561
rect 370 1527 408 1561
rect 442 1527 480 1561
rect 514 1527 552 1561
rect 586 1527 624 1561
rect 658 1527 696 1561
rect 730 1527 768 1561
rect 802 1527 840 1561
rect 874 1527 912 1561
rect 946 1527 984 1561
rect 1018 1527 1056 1561
rect 1090 1527 1128 1561
rect 1162 1527 1200 1561
rect 1234 1527 1272 1561
rect 1306 1527 1344 1561
rect 1378 1527 1416 1561
rect 1450 1527 1488 1561
rect 1522 1527 1560 1561
rect 1594 1527 1632 1561
rect 1666 1527 1704 1561
rect 1738 1527 1776 1561
rect 1810 1527 1848 1561
rect 1882 1527 1920 1561
rect 1954 1527 1992 1561
rect 2026 1527 2064 1561
rect 2098 1527 2136 1561
rect 2170 1527 2208 1561
rect 2242 1527 2280 1561
rect 2314 1527 2352 1561
rect 2386 1527 2424 1561
rect 2458 1527 2496 1561
rect 2530 1527 2568 1561
rect 2602 1527 2640 1561
rect 2674 1527 2712 1561
rect 2746 1527 2784 1561
rect 2818 1527 2856 1561
rect 2890 1527 2928 1561
rect 2962 1527 3000 1561
rect 3034 1527 3072 1561
rect 3106 1527 3144 1561
rect 3178 1527 3216 1561
rect 3250 1527 3288 1561
rect 3322 1527 3360 1561
rect 3394 1527 3432 1561
rect 3466 1527 3504 1561
rect 3538 1527 3576 1561
rect 3610 1527 3648 1561
rect 3682 1527 3840 1561
rect 106 1521 3840 1527
rect 325 1447 3621 1521
rect 106 1377 284 1401
rect 106 1325 176 1377
rect 228 1325 284 1377
rect 106 1301 284 1325
rect 325 1061 3621 1255
rect 106 915 284 1015
rect 106 569 3840 868
rect 106 423 284 523
rect 316 183 1886 377
rect 166 113 280 137
rect 166 61 176 113
rect 228 61 280 113
rect 166 37 280 61
rect 316 -83 1886 -9
rect 106 -89 3840 -83
rect 106 -123 256 -89
rect 290 -123 328 -89
rect 362 -123 400 -89
rect 434 -123 472 -89
rect 506 -123 544 -89
rect 578 -123 616 -89
rect 650 -123 688 -89
rect 722 -123 760 -89
rect 794 -123 832 -89
rect 866 -123 904 -89
rect 938 -123 976 -89
rect 1010 -123 1048 -89
rect 1082 -123 1120 -89
rect 1154 -123 1192 -89
rect 1226 -123 1264 -89
rect 1298 -123 1336 -89
rect 1370 -123 1408 -89
rect 1442 -123 1480 -89
rect 1514 -123 1552 -89
rect 1586 -123 1624 -89
rect 1658 -123 1696 -89
rect 1730 -123 1768 -89
rect 1802 -123 1840 -89
rect 1874 -123 1912 -89
rect 1946 -123 3840 -89
rect 106 -159 3840 -123
<< via1 >>
rect 176 1325 228 1377
rect 176 61 228 113
<< metal2 >>
rect 176 1377 228 1411
rect 176 113 228 1325
rect 176 27 228 61
use sky130_fd_pr__nfet_01v8_X73VMN  sky130_fd_pr__nfet_01v8_X73VMN_0
timestamp 1750100919
transform 0 1 1101 -1 0 87
box -236 -985 236 985
use sky130_fd_pr__pfet_01v8_NMYLRJ  sky130_fd_pr__pfet_01v8_NMYLRJ_0
timestamp 1750100919
transform 0 1 1973 -1 0 965
box -246 -1867 246 1867
use sky130_fd_pr__pfet_01v8_NMYLRJ  XM1
timestamp 1750100919
transform 0 1 1973 -1 0 1351
box -246 -1867 246 1867
use sky130_fd_pr__nfet_01v8_X73VMN  XM3
timestamp 1750100919
transform 0 1 1101 -1 0 473
box -236 -985 236 985
<< labels >>
flabel metal1 s 106 1521 238 1597 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 106 1301 176 1401 0 FreeSans 500 0 0 0 IN
port 2 nsew
flabel metal1 s 106 915 284 1015 0 FreeSans 500 0 0 0 CKB
port 3 nsew
flabel metal1 s 106 423 284 523 0 FreeSans 500 0 0 0 CK
port 4 nsew
flabel metal1 s 106 -159 238 -83 0 FreeSans 500 0 0 0 VSS
port 5 nsew
flabel metal1 s 3667 678 3799 754 0 FreeSans 500 0 0 0 OUT
port 6 nsew
<< end >>
