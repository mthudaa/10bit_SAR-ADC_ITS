../mag/tdc.pex.spice