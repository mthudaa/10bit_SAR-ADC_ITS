* NGSPICE file created from sar8b.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

.subckt sar8b CF[0] CF[1] CF[2] CF[3] CF[4] CF[5] CF[6] CF[7] CKO CKS CKSB CLK CMP_N
+ CMP_P DATA[0] DATA[1] DATA[2] DATA[3] DATA[4] DATA[5] DATA[6] DATA[7] EN RDY SWN[0]
+ SWN[1] SWN[2] SWN[3] SWN[4] SWN[5] SWN[6] SWN[7] SWP[0] SWP[1] SWP[2] SWP[3] SWP[4]
+ SWP[5] SWP[6] SWP[7] VGND VPWR
X_66_ cyclic_flag_0.FINAL net39 net3 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfrtp_1
X_49_ clknet_1_1__leaf_CLK _05_ VGND VGND VPWR VPWR clk_div_0.COUNT\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_5_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput7 net7 VGND VGND VPWR VPWR CF[2] sky130_fd_sc_hd__buf_1
Xoutput20 net20 VGND VGND VPWR VPWR DATA[4] sky130_fd_sc_hd__buf_1
Xoutput31 net31 VGND VGND VPWR VPWR SWN[7] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_65_ net5 net1 net14 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_48_ clknet_1_0__leaf_CLK _04_ VGND VGND VPWR VPWR clk_div_0.COUNT\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput10 net10 VGND VGND VPWR VPWR CF[5] sky130_fd_sc_hd__buf_1
Xoutput8 net8 VGND VGND VPWR VPWR CF[3] sky130_fd_sc_hd__buf_1
Xoutput32 net32 VGND VGND VPWR VPWR SWP[0] sky130_fd_sc_hd__clkbuf_1
Xoutput21 net21 VGND VGND VPWR VPWR DATA[5] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_47_ clknet_1_0__leaf_CLK _03_ VGND VGND VPWR VPWR clk_div_0.COUNT\[1\] sky130_fd_sc_hd__dfxtp_1
X_64_ net6 net1 net14 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput9 net9 VGND VGND VPWR VPWR CF[4] sky130_fd_sc_hd__buf_1
Xoutput11 net11 VGND VGND VPWR VPWR CF[6] sky130_fd_sc_hd__buf_1
Xoutput33 net33 VGND VGND VPWR VPWR SWP[1] sky130_fd_sc_hd__buf_1
Xoutput22 net22 VGND VGND VPWR VPWR DATA[6] sky130_fd_sc_hd__buf_1
XFILLER_0_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_63_ net7 net1 net14 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_46_ clknet_1_0__leaf_CLK _02_ VGND VGND VPWR VPWR clk_div_0.COUNT\[0\] sky130_fd_sc_hd__dfxtp_1
Xoutput23 net23 VGND VGND VPWR VPWR DATA[7] sky130_fd_sc_hd__buf_1
Xoutput12 net12 VGND VGND VPWR VPWR CF[7] sky130_fd_sc_hd__buf_1
Xoutput34 net34 VGND VGND VPWR VPWR SWP[2] sky130_fd_sc_hd__buf_1
X_29_ clk_div_0.COUNT\[0\] clk_div_0.COUNT\[1\] clk_div_0.COUNT\[2\] VGND VGND VPWR
+ VPWR _13_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_62_ net8 net1 net14 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_28_ clk_div_0.COUNT\[0\] clk_div_0.COUNT\[1\] clk_div_0.COUNT\[2\] VGND VGND VPWR
+ VPWR _12_ sky130_fd_sc_hd__nand3_1
X_45_ net4 net12 net14 VGND VGND VPWR VPWR cyclic_flag_0.FINAL sky130_fd_sc_hd__dfrtp_2
Xclkload0 clknet_1_0__leaf_CLK VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput13 net13 VGND VGND VPWR VPWR CKO sky130_fd_sc_hd__buf_1
Xoutput35 net35 VGND VGND VPWR VPWR SWP[3] sky130_fd_sc_hd__buf_1
XFILLER_0_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput24 net24 VGND VGND VPWR VPWR SWN[0] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_8_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_61_ net9 net1 net14 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_1_1__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_1_1__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_44_ net4 net11 net14 VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfrtp_1
X_27_ clk_div_0.COUNT\[0\] clk_div_0.COUNT\[1\] _11_ VGND VGND VPWR VPWR _03_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput36 net36 VGND VGND VPWR VPWR SWP[4] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_15_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput14 net14 VGND VGND VPWR VPWR CKS sky130_fd_sc_hd__buf_1
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput25 net25 VGND VGND VPWR VPWR SWN[1] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_60_ net10 net1 net14 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_26_ clk_div_0.COUNT\[0\] clk_div_0.COUNT\[1\] net3 VGND VGND VPWR VPWR _11_ sky130_fd_sc_hd__o21ai_1
X_43_ net4 net10 net14 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput37 net37 VGND VGND VPWR VPWR SWP[5] sky130_fd_sc_hd__buf_1
Xoutput15 net15 VGND VGND VPWR VPWR CKSB sky130_fd_sc_hd__buf_1
Xoutput26 net26 VGND VGND VPWR VPWR SWN[2] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_42_ net4 net9 net14 VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25_ _10_ VGND VGND VPWR VPWR _02_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput38 net38 VGND VGND VPWR VPWR SWP[6] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput27 net27 VGND VGND VPWR VPWR SWN[3] sky130_fd_sc_hd__buf_1
Xoutput16 net16 VGND VGND VPWR VPWR DATA[0] sky130_fd_sc_hd__buf_1
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_24_ clk_div_0.COUNT\[0\] net3 VGND VGND VPWR VPWR _10_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_9_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_41_ net4 net8 net14 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfrtp_1
Xoutput39 net39 VGND VGND VPWR VPWR SWP[7] sky130_fd_sc_hd__buf_1
XFILLER_0_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput28 net28 VGND VGND VPWR VPWR SWN[4] sky130_fd_sc_hd__buf_1
Xoutput17 net17 VGND VGND VPWR VPWR DATA[1] sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_16_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_40_ net4 net7 net14 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfrtp_1
X_23_ net14 _07_ _09_ VGND VGND VPWR VPWR _01_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_10_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput29 net29 VGND VGND VPWR VPWR SWN[5] sky130_fd_sc_hd__buf_1
Xoutput18 net18 VGND VGND VPWR VPWR DATA[2] sky130_fd_sc_hd__buf_1
X_22_ net14 _07_ net3 VGND VGND VPWR VPWR _09_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_10_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput19 net19 VGND VGND VPWR VPWR DATA[3] sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_21_ net3 _08_ VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20_ net15 _07_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hd__xnor2_1
Xinput1 CMP_N VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_17 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 CMP_P VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 EN VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_2_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 RDY VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_59_ net11 net1 net14 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_58_ net12 net1 net14 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_57_ net5 net2 net14 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_73_ cyclic_flag_0.FINAL net32 net3 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_1
X_56_ net6 net2 net14 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dfrtp_1
X_39_ net4 net6 net14 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_72_ cyclic_flag_0.FINAL net33 net3 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_55_ net7 net2 net14 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfrtp_1
X_38_ net4 net5 net14 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_54_ net8 net2 net14 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfrtp_1
X_71_ cyclic_flag_0.FINAL net34 net3 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_37_ net4 net14 net14 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_13_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_70_ cyclic_flag_0.FINAL net35 net3 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_1
Xclkbuf_0_CLK CLK VGND VGND VPWR VPWR clknet_0_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_53_ net9 net2 net14 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_36_ clknet_1_1__leaf_CLK _01_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dfxtp_4
X_19_ clk_div_0.COUNT\[0\] clk_div_0.COUNT\[1\] clk_div_0.COUNT\[2\] clk_div_0.COUNT\[3\]
+ VGND VGND VPWR VPWR _07_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_52_ net10 net2 net14 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_35_ clknet_1_1__leaf_CLK _00_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18_ _06_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_17_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_51_ net11 net2 net14 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17_ net14 cyclic_flag_0.FINAL VGND VGND VPWR VPWR _06_ sky130_fd_sc_hd__and2_1
X_34_ _16_ VGND VGND VPWR VPWR _05_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_17_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_50_ net12 net2 net14 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_33_ _07_ _15_ net3 VGND VGND VPWR VPWR _16_ sky130_fd_sc_hd__and3b_1
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_32_ clk_div_0.COUNT\[0\] clk_div_0.COUNT\[1\] clk_div_0.COUNT\[2\] clk_div_0.COUNT\[3\]
+ VGND VGND VPWR VPWR _15_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_31_ _14_ VGND VGND VPWR VPWR _04_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30_ net3 _12_ _13_ VGND VGND VPWR VPWR _14_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_69_ cyclic_flag_0.FINAL net36 net3 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_68_ cyclic_flag_0.FINAL net37 net3 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_4_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput5 net5 VGND VGND VPWR VPWR CF[0] sky130_fd_sc_hd__buf_1
XFILLER_0_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f_CLK clknet_0_CLK VGND VGND VPWR VPWR clknet_1_0__leaf_CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_67_ cyclic_flag_0.FINAL net38 net3 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput6 net6 VGND VGND VPWR VPWR CF[1] sky130_fd_sc_hd__buf_1
XFILLER_0_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput30 net30 VGND VGND VPWR VPWR SWN[6] sky130_fd_sc_hd__buf_1
.ends

