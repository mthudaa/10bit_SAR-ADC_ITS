magic
tech sky130A
magscale 1 2
timestamp 1748789218
<< viali >>
rect 142 1527 8084 1561
rect 142 -123 4160 -89
<< metal1 >>
rect 106 1561 8120 1597
rect 106 1527 142 1561
rect 8084 1527 8120 1561
rect 106 1521 8120 1527
rect 325 1447 7901 1521
rect 106 1301 176 1401
rect 228 1301 284 1401
rect 325 1061 7901 1255
rect 106 915 284 1015
rect 106 569 8120 868
rect 106 423 284 523
rect 316 183 3986 377
rect 166 37 176 137
rect 228 37 284 137
rect 316 -83 3986 -9
rect 106 -89 8120 -83
rect 106 -123 142 -89
rect 4160 -123 8120 -89
rect 106 -159 8120 -123
<< via1 >>
rect 176 1301 228 1401
rect 176 37 228 137
<< metal2 >>
rect 176 1401 228 1411
rect 176 137 228 1301
rect 176 27 228 37
use sky130_fd_pr__nfet_01v8_DPTN2D  sky130_fd_pr__nfet_01v8_DPTN2D_0
timestamp 1746262467
transform 0 1 2151 -1 0 87
box -246 -2045 246 2045
use sky130_fd_pr__pfet_01v8_D9QHA6  sky130_fd_pr__pfet_01v8_D9QHA6_0
timestamp 1746262467
transform 0 1 4113 -1 0 965
box -246 -4007 246 4007
use sky130_fd_pr__pfet_01v8_D9QHA6  XM1
timestamp 1746262467
transform 0 1 4113 -1 0 1351
box -246 -4007 246 4007
use sky130_fd_pr__nfet_01v8_DPTN2D  XM3
timestamp 1746262467
transform 0 1 2151 -1 0 473
box -246 -2045 246 2045
<< labels >>
flabel metal1 117 1553 126 1563 0 FreeSans 400 0 0 0 VDD
port 0 nsew
flabel metal1 118 1345 127 1355 0 FreeSans 400 0 0 0 IN
port 1 nsew
flabel metal1 123 958 132 968 0 FreeSans 400 0 0 0 CKB
port 2 nsew
flabel metal1 120 467 129 477 0 FreeSans 400 0 0 0 CK
port 3 nsew
flabel metal1 121 -124 130 -114 0 FreeSans 400 0 0 0 VSS
port 4 nsew
flabel metal1 8079 708 8088 718 0 FreeSans 400 0 0 0 OUT
port 6 nsew
<< end >>
