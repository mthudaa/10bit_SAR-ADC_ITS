magic
tech sky130A
magscale 1 2
timestamp 1749043030
<< nwell >>
rect 213 707 713 827
rect 213 5 319 707
<< pwell >>
rect 344 -441 677 -69
<< psubdiff >>
rect 353 -127 387 -103
rect 353 -259 387 -235
<< nsubdiff >>
rect 265 621 299 645
rect 265 89 299 113
<< psubdiffcont >>
rect 353 -235 387 -127
<< nsubdiffcont >>
rect 265 113 299 621
<< poly >>
rect 163 54 229 70
rect 163 20 179 54
rect 213 52 229 54
rect 413 52 443 58
rect 213 22 443 52
rect 213 20 229 22
rect 163 4 229 20
rect 501 -34 531 76
rect 295 -64 531 -34
rect 589 34 619 90
rect 713 54 779 70
rect 713 34 729 54
rect 589 20 729 34
rect 763 20 779 54
rect 589 4 779 20
rect 589 -55 619 4
rect 163 -95 229 -79
rect 163 -129 179 -95
rect 213 -97 229 -95
rect 295 -97 325 -64
rect 501 -77 531 -64
rect 213 -127 325 -97
rect 213 -129 229 -127
rect 163 -145 229 -129
<< polycont >>
rect 179 20 213 54
rect 729 20 763 54
rect 179 -129 213 -95
<< locali >>
rect 96 761 158 795
rect 192 761 254 795
rect 288 761 350 795
rect 384 761 446 795
rect 480 761 542 795
rect 576 761 638 795
rect 672 761 734 795
rect 768 761 830 795
rect 265 621 299 761
rect 367 636 401 761
rect 631 671 665 761
rect 265 97 299 113
rect 163 54 229 70
rect 163 20 179 54
rect 213 20 229 54
rect 163 4 229 20
rect 543 4 577 67
rect 713 54 779 70
rect 713 20 729 54
rect 763 20 779 54
rect 713 4 779 20
rect 543 -30 665 4
rect 631 -35 665 -30
rect 631 -51 779 -35
rect 631 -69 729 -51
rect 163 -95 229 -79
rect 631 -81 665 -69
rect 163 -129 179 -95
rect 213 -129 229 -95
rect 713 -85 729 -69
rect 763 -85 779 -51
rect 713 -101 779 -85
rect 163 -145 229 -129
rect 353 -127 387 -111
rect 353 -375 387 -235
rect 455 -375 489 -285
rect 96 -409 158 -375
rect 192 -409 254 -375
rect 288 -409 350 -375
rect 384 -409 446 -375
rect 480 -409 542 -375
rect 576 -409 638 -375
rect 672 -409 734 -375
rect 768 -409 830 -375
<< viali >>
rect 158 761 192 795
rect 254 761 288 795
rect 350 761 384 795
rect 446 761 480 795
rect 542 761 576 795
rect 638 761 672 795
rect 734 761 768 795
rect 179 20 213 54
rect 729 20 763 54
rect 179 -129 213 -95
rect 729 -85 763 -51
rect 158 -409 192 -375
rect 254 -409 288 -375
rect 350 -409 384 -375
rect 446 -409 480 -375
rect 542 -409 576 -375
rect 638 -409 672 -375
rect 734 -409 768 -375
<< metal1 >>
rect 96 795 830 827
rect 96 761 158 795
rect 192 761 254 795
rect 288 761 350 795
rect 384 761 446 795
rect 480 761 542 795
rect 576 761 638 795
rect 672 761 734 795
rect 768 761 830 795
rect 96 729 830 761
rect 163 54 229 70
rect 163 20 179 54
rect 213 20 229 54
rect 163 4 229 20
rect 713 54 779 70
rect 713 20 729 54
rect 763 20 779 54
rect 713 4 779 20
rect 713 -51 779 -35
rect 163 -95 229 -79
rect 163 -129 179 -95
rect 213 -129 229 -95
rect 713 -85 729 -51
rect 763 -85 779 -51
rect 713 -101 779 -85
rect 163 -145 229 -129
rect 96 -375 830 -343
rect 96 -409 158 -375
rect 192 -409 254 -375
rect 288 -409 350 -375
rect 384 -409 446 -375
rect 480 -409 542 -375
rect 576 -409 638 -375
rect 672 -409 734 -375
rect 768 -409 830 -375
rect 96 -441 830 -409
use sky130_fd_pr__nfet_01v8_QQ7V57  sky130_fd_pr__nfet_01v8_QQ7V57_0
timestamp 1749010377
transform 1 0 516 0 1 -181
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_QQ7V57  sky130_fd_pr__nfet_01v8_QQ7V57_1
timestamp 1749010377
transform 1 0 604 0 1 -181
box -73 -126 73 126
use sky130_fd_pr__pfet_01v8_5EUKDE  sky130_fd_pr__pfet_01v8_5EUKDE_0
timestamp 1749010377
transform 1 0 604 0 1 367
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_5EUKDE  sky130_fd_pr__pfet_01v8_5EUKDE_1
timestamp 1749010377
transform 1 0 516 0 1 367
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_5EUKDE  sky130_fd_pr__pfet_01v8_5EUKDE_2
timestamp 1749010377
transform 1 0 428 0 1 367
box -109 -362 109 362
<< labels >>
flabel metal1 96 729 158 827 0 FreeSans 400 0 0 0 VDD
port 4 nsew
flabel metal1 96 -441 158 -343 0 FreeSans 400 0 0 0 VSS
port 5 nsew
flabel metal1 179 20 213 54 0 FreeSans 400 0 0 0 INB
port 8 nsew
flabel metal1 179 -129 213 -95 0 FreeSans 400 0 0 0 IN
port 9 nsew
flabel metal1 729 20 763 54 0 FreeSans 400 0 0 0 OUTB
port 10 nsew
flabel viali 729 -85 763 -51 0 FreeSans 400 0 0 0 OUT
port 3 nsew
<< end >>
