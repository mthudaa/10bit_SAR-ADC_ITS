magic
tech sky130A
magscale 1 2
timestamp 1749411235
<< viali >>
rect 1567 25846 1601 25880
rect 2143 25846 2177 25880
rect 2719 25846 2753 25880
rect 3295 25846 3329 25880
rect 3871 25846 3905 25880
rect 4447 25846 4481 25880
rect 5023 25846 5057 25880
rect 5599 25846 5633 25880
rect 6271 25846 6305 25880
rect 6751 25846 6785 25880
rect 7327 25846 7361 25880
rect 7903 25846 7937 25880
rect 8479 25846 8513 25880
rect 9055 25846 9089 25880
rect 9631 25846 9665 25880
rect 1759 25624 1793 25658
rect 2431 25624 2465 25658
rect 3007 25624 3041 25658
rect 3583 25624 3617 25658
rect 4159 25624 4193 25658
rect 4735 25624 4769 25658
rect 5311 25624 5345 25658
rect 5887 25624 5921 25658
rect 5983 25624 6017 25658
rect 6943 25624 6977 25658
rect 7519 25624 7553 25658
rect 8095 25624 8129 25658
rect 8671 25624 8705 25658
rect 9247 25624 9281 25658
rect 9823 25624 9857 25658
rect 1567 25180 1601 25214
rect 9343 25180 9377 25214
rect 10111 25180 10145 25214
rect 1951 25106 1985 25140
rect 9727 25106 9761 25140
rect 1855 24958 1889 24992
rect 2239 24958 2273 24992
rect 9151 24958 9185 24992
rect 9439 24958 9473 24992
rect 9823 24958 9857 24992
rect 1567 24440 1601 24474
rect 6751 24440 6785 24474
rect 10111 24440 10145 24474
rect 1759 24292 1793 24326
rect 5215 24292 5249 24326
rect 9823 24292 9857 24326
rect 4831 24218 4865 24252
rect 6175 23848 6209 23882
rect 7711 23700 7745 23734
rect 4543 23626 4577 23660
rect 8095 23626 8129 23660
rect 4159 23552 4193 23586
rect 9727 23404 9761 23438
rect 3295 22960 3329 22994
rect 5503 22960 5537 22994
rect 7135 22960 7169 22994
rect 9055 22960 9089 22994
rect 9343 22960 9377 22994
rect 9823 22960 9857 22994
rect 3679 22886 3713 22920
rect 5119 22886 5153 22920
rect 8287 22886 8321 22920
rect 8479 22812 8513 22846
rect 1663 22738 1697 22772
rect 8095 22738 8129 22772
rect 10111 22738 10145 22772
rect 1567 22516 1601 22550
rect 4255 22516 4289 22550
rect 2239 22368 2273 22402
rect 7711 22368 7745 22402
rect 1855 22294 1889 22328
rect 2623 22294 2657 22328
rect 8095 22294 8129 22328
rect 9727 22072 9761 22106
rect 6943 21850 6977 21884
rect 1759 21702 1793 21736
rect 3295 21628 3329 21662
rect 3679 21628 3713 21662
rect 4927 21628 4961 21662
rect 5311 21628 5345 21662
rect 4255 21184 4289 21218
rect 2239 21036 2273 21070
rect 2623 20962 2657 20996
rect 6943 20962 6977 20996
rect 7327 20962 7361 20996
rect 8959 20740 8993 20774
rect 6751 20370 6785 20404
rect 7135 20296 7169 20330
rect 9823 20296 9857 20330
rect 8767 20148 8801 20182
rect 10111 20148 10145 20182
rect 6943 19704 6977 19738
rect 7327 19630 7361 19664
rect 8959 19408 8993 19442
rect 1663 18890 1697 18924
rect 1759 18742 1793 18776
rect 2815 18520 2849 18554
rect 4831 18372 4865 18406
rect 7519 18372 7553 18406
rect 4447 18298 4481 18332
rect 7903 18298 7937 18332
rect 9535 18298 9569 18332
rect 9823 18298 9857 18332
rect 10111 18076 10145 18110
rect 3583 17854 3617 17888
rect 5791 17854 5825 17888
rect 3871 17706 3905 17740
rect 1951 17632 1985 17666
rect 4255 17632 4289 17666
rect 1567 17558 1601 17592
rect 5791 17188 5825 17222
rect 7423 17040 7457 17074
rect 4159 16966 4193 17000
rect 7807 16966 7841 17000
rect 3775 16892 3809 16926
rect 9439 16744 9473 16778
rect 8191 16522 8225 16556
rect 3679 16374 3713 16408
rect 3295 16300 3329 16334
rect 4255 16300 4289 16334
rect 6463 16300 6497 16334
rect 3871 16226 3905 16260
rect 6079 16226 6113 16260
rect 1663 16078 1697 16112
rect 5887 16078 5921 16112
rect 3775 15708 3809 15742
rect 7519 15708 7553 15742
rect 3391 15634 3425 15668
rect 7903 15634 7937 15668
rect 9535 15634 9569 15668
rect 9823 15634 9857 15668
rect 1759 15412 1793 15446
rect 10111 15412 10145 15446
rect 6751 15042 6785 15076
rect 7135 14968 7169 15002
rect 8767 14746 8801 14780
rect 7423 14376 7457 14410
rect 7807 14302 7841 14336
rect 1663 14228 1697 14262
rect 1759 14228 1793 14262
rect 9439 14080 9473 14114
rect 9823 13636 9857 13670
rect 10111 13414 10145 13448
rect 4735 13192 4769 13226
rect 2719 13044 2753 13078
rect 3103 12970 3137 13004
rect 7039 12526 7073 12560
rect 5119 12378 5153 12412
rect 1951 12304 1985 12338
rect 5503 12304 5537 12338
rect 1567 12230 1601 12264
rect 3583 12082 3617 12116
rect 2623 11860 2657 11894
rect 8479 11860 8513 11894
rect 4639 11712 4673 11746
rect 6463 11712 6497 11746
rect 4255 11638 4289 11672
rect 6847 11638 6881 11672
rect 8671 11194 8705 11228
rect 4543 11046 4577 11080
rect 6751 11046 6785 11080
rect 1951 10972 1985 11006
rect 4927 10972 4961 11006
rect 7135 10972 7169 11006
rect 9823 10972 9857 11006
rect 1567 10898 1601 10932
rect 3583 10750 3617 10784
rect 6559 10750 6593 10784
rect 10111 10750 10145 10784
rect 1951 10528 1985 10562
rect 8671 10528 8705 10562
rect 1663 10380 1697 10414
rect 3391 10380 3425 10414
rect 6655 10380 6689 10414
rect 3775 10306 3809 10340
rect 7039 10306 7073 10340
rect 5407 10084 5441 10118
rect 8479 9862 8513 9896
rect 6943 9640 6977 9674
rect 6559 9566 6593 9600
rect 8191 8974 8225 9008
rect 7807 8900 7841 8934
rect 9727 8752 9761 8786
rect 6751 8382 6785 8416
rect 3679 8308 3713 8342
rect 7135 8308 7169 8342
rect 9823 8308 9857 8342
rect 10111 8308 10145 8342
rect 8767 8086 8801 8120
rect 3679 7864 3713 7898
rect 3199 7716 3233 7750
rect 4447 7716 4481 7750
rect 7423 7716 7457 7750
rect 2623 7642 2657 7676
rect 2815 7642 2849 7676
rect 2911 7642 2945 7676
rect 3583 7642 3617 7676
rect 3967 7642 4001 7676
rect 7807 7642 7841 7676
rect 3775 7568 3809 7602
rect 2431 7420 2465 7454
rect 3007 7420 3041 7454
rect 4063 7420 4097 7454
rect 9439 7420 9473 7454
rect 3487 7198 3521 7232
rect 2335 7050 2369 7084
rect 1663 6976 1697 7010
rect 1951 6976 1985 7010
rect 4063 6976 4097 7010
rect 4159 6976 4193 7010
rect 4735 6976 4769 7010
rect 5023 6976 5057 7010
rect 5215 6976 5249 7010
rect 5407 6976 5441 7010
rect 6367 6976 6401 7010
rect 4543 6902 4577 6936
rect 5983 6902 6017 6936
rect 1855 6754 1889 6788
rect 3871 6754 3905 6788
rect 4831 6754 4865 6788
rect 5311 6754 5345 6788
rect 7999 6754 8033 6788
rect 1951 6532 1985 6566
rect 2335 6532 2369 6566
rect 2527 6532 2561 6566
rect 4639 6532 4673 6566
rect 2815 6458 2849 6492
rect 5311 6458 5345 6492
rect 5695 6458 5729 6492
rect 1567 6384 1601 6418
rect 2143 6384 2177 6418
rect 2623 6384 2657 6418
rect 3295 6384 3329 6418
rect 4831 6384 4865 6418
rect 5599 6384 5633 6418
rect 5791 6384 5825 6418
rect 1759 6310 1793 6344
rect 1855 6310 1889 6344
rect 2911 6310 2945 6344
rect 5119 6310 5153 6344
rect 9823 6310 9857 6344
rect 1855 6162 1889 6196
rect 10111 6088 10145 6122
rect 5791 5866 5825 5900
rect 2527 5718 2561 5752
rect 1759 5644 1793 5678
rect 2143 5644 2177 5678
rect 3871 5644 3905 5678
rect 5983 5644 6017 5678
rect 6559 5644 6593 5678
rect 6079 5570 6113 5604
rect 6367 5570 6401 5604
rect 6655 5570 6689 5604
rect 6463 5496 6497 5530
rect 2047 5422 2081 5456
rect 3679 5422 3713 5456
rect 6079 5422 6113 5456
rect 5407 5200 5441 5234
rect 6751 5200 6785 5234
rect 2239 5126 2273 5160
rect 5983 5126 6017 5160
rect 4255 5052 4289 5086
rect 5503 5052 5537 5086
rect 6655 5052 6689 5086
rect 3775 4978 3809 5012
rect 3871 4978 3905 5012
rect 5791 4978 5825 5012
rect 3391 4904 3425 4938
rect 6463 4830 6497 4864
rect 1759 4312 1793 4346
rect 4543 4312 4577 4346
rect 1567 4090 1601 4124
rect 5407 3868 5441 3902
rect 4255 3720 4289 3754
rect 2143 3646 2177 3680
rect 3871 3646 3905 3680
rect 9535 3646 9569 3680
rect 9919 3646 9953 3680
rect 10111 3572 10145 3606
rect 1855 3424 1889 3458
rect 9727 3424 9761 3458
rect 1951 3202 1985 3236
rect 1567 2980 1601 3014
rect 3199 2980 3233 3014
rect 4447 2980 4481 3014
rect 5599 2980 5633 3014
rect 6655 2980 6689 3014
rect 7903 2980 7937 3014
rect 9247 2980 9281 3014
rect 9439 2980 9473 3014
rect 10015 2980 10049 3014
rect 3007 2906 3041 2940
rect 4159 2906 4193 2940
rect 5311 2906 5345 2940
rect 6463 2906 6497 2940
rect 7615 2906 7649 2940
rect 9055 2906 9089 2940
rect 9727 2906 9761 2940
rect 9823 2906 9857 2940
<< metal1 >>
rect 1152 26000 10560 26022
rect 1152 25948 1966 26000
rect 2018 25948 2030 26000
rect 2082 25948 2094 26000
rect 2146 25948 2158 26000
rect 2210 25948 2222 26000
rect 2274 25948 2286 26000
rect 2338 25948 7966 26000
rect 8018 25948 8030 26000
rect 8082 25948 8094 26000
rect 8146 25948 8158 26000
rect 8210 25948 8222 26000
rect 8274 25948 8286 26000
rect 8338 25948 10560 26000
rect 1152 25926 10560 25948
rect 1552 25837 1558 25889
rect 1610 25837 1616 25889
rect 1840 25837 1846 25889
rect 1898 25877 1904 25889
rect 2131 25880 2189 25886
rect 2131 25877 2143 25880
rect 1898 25849 2143 25877
rect 1898 25837 1904 25849
rect 2131 25846 2143 25849
rect 2177 25846 2189 25880
rect 2131 25840 2189 25846
rect 2608 25837 2614 25889
rect 2666 25877 2672 25889
rect 2707 25880 2765 25886
rect 2707 25877 2719 25880
rect 2666 25849 2719 25877
rect 2666 25837 2672 25849
rect 2707 25846 2719 25849
rect 2753 25846 2765 25880
rect 2707 25840 2765 25846
rect 3280 25837 3286 25889
rect 3338 25837 3344 25889
rect 3856 25837 3862 25889
rect 3914 25837 3920 25889
rect 4432 25837 4438 25889
rect 4490 25837 4496 25889
rect 5008 25837 5014 25889
rect 5066 25837 5072 25889
rect 5488 25837 5494 25889
rect 5546 25877 5552 25889
rect 5587 25880 5645 25886
rect 5587 25877 5599 25880
rect 5546 25849 5599 25877
rect 5546 25837 5552 25849
rect 5587 25846 5599 25849
rect 5633 25846 5645 25880
rect 5587 25840 5645 25846
rect 6256 25837 6262 25889
rect 6314 25837 6320 25889
rect 6736 25837 6742 25889
rect 6794 25837 6800 25889
rect 7312 25837 7318 25889
rect 7370 25837 7376 25889
rect 7888 25837 7894 25889
rect 7946 25837 7952 25889
rect 8464 25837 8470 25889
rect 8522 25837 8528 25889
rect 9040 25837 9046 25889
rect 9098 25837 9104 25889
rect 9616 25837 9622 25889
rect 9674 25837 9680 25889
rect 5968 25803 5974 25815
rect 3586 25775 5974 25803
rect 1648 25615 1654 25667
rect 1706 25655 1712 25667
rect 1747 25658 1805 25664
rect 1747 25655 1759 25658
rect 1706 25627 1759 25655
rect 1706 25615 1712 25627
rect 1747 25624 1759 25627
rect 1793 25624 1805 25658
rect 1747 25618 1805 25624
rect 2419 25658 2477 25664
rect 2419 25624 2431 25658
rect 2465 25655 2477 25658
rect 2896 25655 2902 25667
rect 2465 25627 2902 25655
rect 2465 25624 2477 25627
rect 2419 25618 2477 25624
rect 2896 25615 2902 25627
rect 2954 25615 2960 25667
rect 2992 25615 2998 25667
rect 3050 25615 3056 25667
rect 3586 25664 3614 25775
rect 5968 25763 5974 25775
rect 6026 25763 6032 25815
rect 3664 25689 3670 25741
rect 3722 25729 3728 25741
rect 3722 25701 6014 25729
rect 3722 25689 3728 25701
rect 3571 25658 3629 25664
rect 3571 25624 3583 25658
rect 3617 25624 3629 25658
rect 3571 25618 3629 25624
rect 4147 25658 4205 25664
rect 4147 25624 4159 25658
rect 4193 25624 4205 25658
rect 4147 25618 4205 25624
rect 4723 25658 4781 25664
rect 4723 25624 4735 25658
rect 4769 25624 4781 25658
rect 4723 25618 4781 25624
rect 5299 25658 5357 25664
rect 5299 25624 5311 25658
rect 5345 25655 5357 25658
rect 5776 25655 5782 25667
rect 5345 25627 5782 25655
rect 5345 25624 5357 25627
rect 5299 25618 5357 25624
rect 4162 25507 4190 25618
rect 4738 25581 4766 25618
rect 5776 25615 5782 25627
rect 5834 25615 5840 25667
rect 5872 25615 5878 25667
rect 5930 25615 5936 25667
rect 5986 25664 6014 25701
rect 5971 25658 6029 25664
rect 5971 25624 5983 25658
rect 6017 25624 6029 25658
rect 5971 25618 6029 25624
rect 6928 25615 6934 25667
rect 6986 25615 6992 25667
rect 7504 25615 7510 25667
rect 7562 25615 7568 25667
rect 8080 25615 8086 25667
rect 8138 25615 8144 25667
rect 8659 25658 8717 25664
rect 8659 25624 8671 25658
rect 8705 25624 8717 25658
rect 8659 25618 8717 25624
rect 7216 25581 7222 25593
rect 4738 25553 7222 25581
rect 7216 25541 7222 25553
rect 7274 25541 7280 25593
rect 6736 25507 6742 25519
rect 4162 25479 6742 25507
rect 6736 25467 6742 25479
rect 6794 25467 6800 25519
rect 5392 25393 5398 25445
rect 5450 25433 5456 25445
rect 8674 25433 8702 25618
rect 9232 25615 9238 25667
rect 9290 25615 9296 25667
rect 9712 25615 9718 25667
rect 9770 25655 9776 25667
rect 9811 25658 9869 25664
rect 9811 25655 9823 25658
rect 9770 25627 9823 25655
rect 9770 25615 9776 25627
rect 9811 25624 9823 25627
rect 9857 25624 9869 25658
rect 9811 25618 9869 25624
rect 5450 25405 8702 25433
rect 5450 25393 5456 25405
rect 1152 25334 10560 25356
rect 1152 25282 4966 25334
rect 5018 25282 5030 25334
rect 5082 25282 5094 25334
rect 5146 25282 5158 25334
rect 5210 25282 5222 25334
rect 5274 25282 5286 25334
rect 5338 25282 10560 25334
rect 1152 25260 10560 25282
rect 1456 25171 1462 25223
rect 1514 25211 1520 25223
rect 1555 25214 1613 25220
rect 1555 25211 1567 25214
rect 1514 25183 1567 25211
rect 1514 25171 1520 25183
rect 1555 25180 1567 25183
rect 1601 25180 1613 25214
rect 1555 25174 1613 25180
rect 3280 25171 3286 25223
rect 3338 25211 3344 25223
rect 6928 25211 6934 25223
rect 3338 25183 6934 25211
rect 3338 25171 3344 25183
rect 6928 25171 6934 25183
rect 6986 25171 6992 25223
rect 9328 25171 9334 25223
rect 9386 25171 9392 25223
rect 10096 25171 10102 25223
rect 10154 25171 10160 25223
rect 304 25097 310 25149
rect 362 25137 368 25149
rect 1939 25140 1997 25146
rect 1939 25137 1951 25140
rect 362 25109 1951 25137
rect 362 25097 368 25109
rect 1939 25106 1951 25109
rect 1985 25106 1997 25140
rect 1939 25100 1997 25106
rect 3376 25097 3382 25149
rect 3434 25137 3440 25149
rect 7504 25137 7510 25149
rect 3434 25109 7510 25137
rect 3434 25097 3440 25109
rect 7504 25097 7510 25109
rect 7562 25097 7568 25149
rect 9715 25140 9773 25146
rect 9715 25106 9727 25140
rect 9761 25137 9773 25140
rect 10672 25137 10678 25149
rect 9761 25109 10678 25137
rect 9761 25106 9773 25109
rect 9715 25100 9773 25106
rect 10672 25097 10678 25109
rect 10730 25097 10736 25149
rect 2608 25023 2614 25075
rect 2666 25063 2672 25075
rect 8080 25063 8086 25075
rect 2666 25035 8086 25063
rect 2666 25023 2672 25035
rect 8080 25023 8086 25035
rect 8138 25023 8144 25075
rect 1840 24949 1846 25001
rect 1898 24949 1904 25001
rect 2227 24992 2285 24998
rect 2227 24958 2239 24992
rect 2273 24989 2285 24992
rect 4240 24989 4246 25001
rect 2273 24961 4246 24989
rect 2273 24958 2285 24961
rect 2227 24952 2285 24958
rect 4240 24949 4246 24961
rect 4298 24949 4304 25001
rect 9139 24992 9197 24998
rect 9139 24958 9151 24992
rect 9185 24989 9197 24992
rect 9328 24989 9334 25001
rect 9185 24961 9334 24989
rect 9185 24958 9197 24961
rect 9139 24952 9197 24958
rect 9328 24949 9334 24961
rect 9386 24949 9392 25001
rect 9424 24949 9430 25001
rect 9482 24949 9488 25001
rect 9811 24992 9869 24998
rect 9811 24958 9823 24992
rect 9857 24958 9869 24992
rect 9811 24952 9869 24958
rect 6832 24875 6838 24927
rect 6890 24915 6896 24927
rect 9826 24915 9854 24952
rect 6890 24887 9854 24915
rect 6890 24875 6896 24887
rect 1152 24668 10560 24690
rect 1152 24616 1966 24668
rect 2018 24616 2030 24668
rect 2082 24616 2094 24668
rect 2146 24616 2158 24668
rect 2210 24616 2222 24668
rect 2274 24616 2286 24668
rect 2338 24616 7966 24668
rect 8018 24616 8030 24668
rect 8082 24616 8094 24668
rect 8146 24616 8158 24668
rect 8210 24616 8222 24668
rect 8274 24616 8286 24668
rect 8338 24616 10560 24668
rect 1152 24594 10560 24616
rect 880 24431 886 24483
rect 938 24471 944 24483
rect 1555 24474 1613 24480
rect 1555 24471 1567 24474
rect 938 24443 1567 24471
rect 938 24431 944 24443
rect 1555 24440 1567 24443
rect 1601 24440 1613 24474
rect 1555 24434 1613 24440
rect 6736 24431 6742 24483
rect 6794 24431 6800 24483
rect 10099 24474 10157 24480
rect 10099 24440 10111 24474
rect 10145 24471 10157 24474
rect 11248 24471 11254 24483
rect 10145 24443 11254 24471
rect 10145 24440 10157 24443
rect 10099 24434 10157 24440
rect 11248 24431 11254 24443
rect 11306 24431 11312 24483
rect 6064 24357 6070 24409
rect 6122 24357 6128 24409
rect 9712 24397 9718 24409
rect 7810 24369 9718 24397
rect 7810 24335 7838 24369
rect 9712 24357 9718 24369
rect 9770 24357 9776 24409
rect 1744 24283 1750 24335
rect 1802 24283 1808 24335
rect 5203 24326 5261 24332
rect 5203 24292 5215 24326
rect 5249 24323 5261 24326
rect 7792 24323 7798 24335
rect 5249 24295 7798 24323
rect 5249 24292 5261 24295
rect 5203 24286 5261 24292
rect 7792 24283 7798 24295
rect 7850 24283 7856 24335
rect 8464 24283 8470 24335
rect 8522 24323 8528 24335
rect 9811 24326 9869 24332
rect 9811 24323 9823 24326
rect 8522 24295 9823 24323
rect 8522 24283 8528 24295
rect 9811 24292 9823 24295
rect 9857 24292 9869 24326
rect 9811 24286 9869 24292
rect 4144 24209 4150 24261
rect 4202 24249 4208 24261
rect 4819 24252 4877 24258
rect 4819 24249 4831 24252
rect 4202 24221 4831 24249
rect 4202 24209 4208 24221
rect 4819 24218 4831 24221
rect 4865 24218 4877 24252
rect 4819 24212 4877 24218
rect 6736 24061 6742 24113
rect 6794 24101 6800 24113
rect 8560 24101 8566 24113
rect 6794 24073 8566 24101
rect 6794 24061 6800 24073
rect 8560 24061 8566 24073
rect 8618 24061 8624 24113
rect 1152 24002 10560 24024
rect 1152 23950 4966 24002
rect 5018 23950 5030 24002
rect 5082 23950 5094 24002
rect 5146 23950 5158 24002
rect 5210 23950 5222 24002
rect 5274 23950 5286 24002
rect 5338 23950 10560 24002
rect 1152 23928 10560 23950
rect 5872 23839 5878 23891
rect 5930 23879 5936 23891
rect 6163 23882 6221 23888
rect 6163 23879 6175 23882
rect 5930 23851 6175 23879
rect 5930 23839 5936 23851
rect 6163 23848 6175 23851
rect 6209 23879 6221 23882
rect 6209 23851 7742 23879
rect 6209 23848 6221 23851
rect 6163 23842 6221 23848
rect 7714 23740 7742 23851
rect 7699 23734 7757 23740
rect 7699 23700 7711 23734
rect 7745 23700 7757 23734
rect 7699 23694 7757 23700
rect 4531 23660 4589 23666
rect 4531 23626 4543 23660
rect 4577 23657 4589 23660
rect 8083 23660 8141 23666
rect 4577 23629 7214 23657
rect 4577 23626 4589 23629
rect 4531 23620 4589 23626
rect 4144 23543 4150 23595
rect 4202 23543 4208 23595
rect 6064 23583 6070 23595
rect 5712 23555 6070 23583
rect 6064 23543 6070 23555
rect 6122 23543 6128 23595
rect 7186 23509 7214 23629
rect 8083 23626 8095 23660
rect 8129 23657 8141 23660
rect 8368 23657 8374 23669
rect 8129 23629 8374 23657
rect 8129 23626 8141 23629
rect 8083 23620 8141 23626
rect 8368 23617 8374 23629
rect 8426 23617 8432 23669
rect 7894 23595 7946 23601
rect 7894 23537 7946 23543
rect 8464 23509 8470 23521
rect 7186 23481 8470 23509
rect 8464 23469 8470 23481
rect 8522 23469 8528 23521
rect 9715 23438 9773 23444
rect 9715 23404 9727 23438
rect 9761 23435 9773 23438
rect 9808 23435 9814 23447
rect 9761 23407 9814 23435
rect 9761 23404 9773 23407
rect 9715 23398 9773 23404
rect 9808 23395 9814 23407
rect 9866 23395 9872 23447
rect 1152 23336 10560 23358
rect 1152 23284 1966 23336
rect 2018 23284 2030 23336
rect 2082 23284 2094 23336
rect 2146 23284 2158 23336
rect 2210 23284 2222 23336
rect 2274 23284 2286 23336
rect 2338 23284 7966 23336
rect 8018 23284 8030 23336
rect 8082 23284 8094 23336
rect 8146 23284 8158 23336
rect 8210 23284 8222 23336
rect 8274 23284 8286 23336
rect 8338 23284 10560 23336
rect 1152 23262 10560 23284
rect 3490 23111 6110 23139
rect 3490 23083 3518 23111
rect 6082 23083 6110 23111
rect 3478 23077 3530 23083
rect 3478 23019 3530 23025
rect 6070 23077 6122 23083
rect 6070 23019 6122 23025
rect 3283 22994 3341 23000
rect 3283 22960 3295 22994
rect 3329 22991 3341 22994
rect 3376 22991 3382 23003
rect 3329 22963 3382 22991
rect 3329 22960 3341 22963
rect 3283 22954 3341 22960
rect 3376 22951 3382 22963
rect 3434 22951 3440 23003
rect 5491 22994 5549 23000
rect 5491 22960 5503 22994
rect 5537 22960 5549 22994
rect 5491 22954 5549 22960
rect 3667 22920 3725 22926
rect 3667 22886 3679 22920
rect 3713 22917 3725 22920
rect 3760 22917 3766 22929
rect 3713 22889 3766 22917
rect 3713 22886 3725 22889
rect 3667 22880 3725 22886
rect 3760 22877 3766 22889
rect 3818 22917 3824 22929
rect 4144 22917 4150 22929
rect 3818 22889 4150 22917
rect 3818 22877 3824 22889
rect 4144 22877 4150 22889
rect 4202 22917 4208 22929
rect 5107 22920 5165 22926
rect 5107 22917 5119 22920
rect 4202 22889 5119 22917
rect 4202 22877 4208 22889
rect 5107 22886 5119 22889
rect 5153 22886 5165 22920
rect 5506 22917 5534 22954
rect 5776 22951 5782 23003
rect 5834 22991 5840 23003
rect 7120 22991 7126 23003
rect 5834 22963 7126 22991
rect 5834 22951 5840 22963
rect 7120 22951 7126 22963
rect 7178 22951 7184 23003
rect 9043 22994 9101 23000
rect 9043 22991 9055 22994
rect 8482 22963 9055 22991
rect 6832 22917 6838 22929
rect 5506 22889 6838 22917
rect 5107 22880 5165 22886
rect 6832 22877 6838 22889
rect 6890 22917 6896 22929
rect 6890 22889 8222 22917
rect 6890 22877 6896 22889
rect 1648 22729 1654 22781
rect 1706 22769 1712 22781
rect 2704 22769 2710 22781
rect 1706 22741 2710 22769
rect 1706 22729 1712 22741
rect 2704 22729 2710 22741
rect 2762 22729 2768 22781
rect 6064 22729 6070 22781
rect 6122 22769 6128 22781
rect 8083 22772 8141 22778
rect 8083 22769 8095 22772
rect 6122 22741 8095 22769
rect 6122 22729 6128 22741
rect 8083 22738 8095 22741
rect 8129 22738 8141 22772
rect 8194 22769 8222 22889
rect 8272 22877 8278 22929
rect 8330 22877 8336 22929
rect 8482 22852 8510 22963
rect 9043 22960 9055 22963
rect 9089 22960 9101 22994
rect 9043 22954 9101 22960
rect 9328 22951 9334 23003
rect 9386 22951 9392 23003
rect 9808 22951 9814 23003
rect 9866 22951 9872 23003
rect 8467 22846 8525 22852
rect 8467 22812 8479 22846
rect 8513 22812 8525 22846
rect 8467 22806 8525 22812
rect 9424 22769 9430 22781
rect 8194 22741 9430 22769
rect 8083 22732 8141 22738
rect 9424 22729 9430 22741
rect 9482 22729 9488 22781
rect 10096 22729 10102 22781
rect 10154 22729 10160 22781
rect 1152 22670 10560 22692
rect 1152 22618 4966 22670
rect 5018 22618 5030 22670
rect 5082 22618 5094 22670
rect 5146 22618 5158 22670
rect 5210 22618 5222 22670
rect 5274 22618 5286 22670
rect 5338 22618 10560 22670
rect 1152 22596 10560 22618
rect 1264 22507 1270 22559
rect 1322 22547 1328 22559
rect 1555 22550 1613 22556
rect 1555 22547 1567 22550
rect 1322 22519 1567 22547
rect 1322 22507 1328 22519
rect 1555 22516 1567 22519
rect 1601 22516 1613 22550
rect 1555 22510 1613 22516
rect 4240 22507 4246 22559
rect 4298 22507 4304 22559
rect 7792 22507 7798 22559
rect 7850 22547 7856 22559
rect 8464 22547 8470 22559
rect 7850 22519 8470 22547
rect 7850 22507 7856 22519
rect 8464 22507 8470 22519
rect 8522 22507 8528 22559
rect 2227 22402 2285 22408
rect 2227 22368 2239 22402
rect 2273 22399 2285 22402
rect 3760 22399 3766 22411
rect 2273 22371 3766 22399
rect 2273 22368 2285 22371
rect 2227 22362 2285 22368
rect 3760 22359 3766 22371
rect 3818 22359 3824 22411
rect 7120 22359 7126 22411
rect 7178 22399 7184 22411
rect 7699 22402 7757 22408
rect 7699 22399 7711 22402
rect 7178 22371 7711 22399
rect 7178 22359 7184 22371
rect 7699 22368 7711 22371
rect 7745 22368 7757 22402
rect 7699 22362 7757 22368
rect 1843 22328 1901 22334
rect 1843 22294 1855 22328
rect 1889 22294 1901 22328
rect 1843 22288 1901 22294
rect 2611 22328 2669 22334
rect 2611 22294 2623 22328
rect 2657 22325 2669 22328
rect 3664 22325 3670 22337
rect 2657 22297 3670 22325
rect 2657 22294 2669 22297
rect 2611 22288 2669 22294
rect 1858 22177 1886 22288
rect 3664 22285 3670 22297
rect 3722 22285 3728 22337
rect 7312 22285 7318 22337
rect 7370 22325 7376 22337
rect 8083 22328 8141 22334
rect 8083 22325 8095 22328
rect 7370 22297 8095 22325
rect 7370 22285 7376 22297
rect 8083 22294 8095 22297
rect 8129 22325 8141 22328
rect 8272 22325 8278 22337
rect 8129 22297 8278 22325
rect 8129 22294 8141 22297
rect 8083 22288 8141 22294
rect 8272 22285 8278 22297
rect 8330 22285 8336 22337
rect 7894 22263 7946 22269
rect 3472 22211 3478 22263
rect 3530 22211 3536 22263
rect 3490 22177 3518 22211
rect 7894 22205 7946 22211
rect 1858 22149 3518 22177
rect 9715 22106 9773 22112
rect 9715 22072 9727 22106
rect 9761 22103 9773 22106
rect 9808 22103 9814 22115
rect 9761 22075 9814 22103
rect 9761 22072 9773 22075
rect 9715 22066 9773 22072
rect 9808 22063 9814 22075
rect 9866 22063 9872 22115
rect 1152 22004 10560 22026
rect 1152 21952 1966 22004
rect 2018 21952 2030 22004
rect 2082 21952 2094 22004
rect 2146 21952 2158 22004
rect 2210 21952 2222 22004
rect 2274 21952 2286 22004
rect 2338 21952 7966 22004
rect 8018 21952 8030 22004
rect 8082 21952 8094 22004
rect 8146 21952 8158 22004
rect 8210 21952 8222 22004
rect 8274 21952 8286 22004
rect 8338 21952 10560 22004
rect 1152 21930 10560 21952
rect 6931 21884 6989 21890
rect 6931 21850 6943 21884
rect 6977 21881 6989 21884
rect 7216 21881 7222 21893
rect 6977 21853 7222 21881
rect 6977 21850 6989 21853
rect 6931 21844 6989 21850
rect 7216 21841 7222 21853
rect 7274 21881 7280 21893
rect 7504 21881 7510 21893
rect 7274 21853 7510 21881
rect 7274 21841 7280 21853
rect 7504 21841 7510 21853
rect 7562 21841 7568 21893
rect 3478 21745 3530 21751
rect 1744 21693 1750 21745
rect 1802 21693 1808 21745
rect 6064 21693 6070 21745
rect 6122 21693 6128 21745
rect 3478 21687 3530 21693
rect 3280 21619 3286 21671
rect 3338 21619 3344 21671
rect 3667 21662 3725 21668
rect 3667 21628 3679 21662
rect 3713 21659 3725 21662
rect 3760 21659 3766 21671
rect 3713 21631 3766 21659
rect 3713 21628 3725 21631
rect 3667 21622 3725 21628
rect 3760 21619 3766 21631
rect 3818 21659 3824 21671
rect 4915 21662 4973 21668
rect 4915 21659 4927 21662
rect 3818 21631 4927 21659
rect 3818 21619 3824 21631
rect 4915 21628 4927 21631
rect 4961 21628 4973 21662
rect 4915 21622 4973 21628
rect 5299 21662 5357 21668
rect 5299 21628 5311 21662
rect 5345 21659 5357 21662
rect 6736 21659 6742 21671
rect 5345 21631 6742 21659
rect 5345 21628 5357 21631
rect 5299 21622 5357 21628
rect 6736 21619 6742 21631
rect 6794 21619 6800 21671
rect 1152 21338 10560 21360
rect 1152 21286 4966 21338
rect 5018 21286 5030 21338
rect 5082 21286 5094 21338
rect 5146 21286 5158 21338
rect 5210 21286 5222 21338
rect 5274 21286 5286 21338
rect 5338 21286 10560 21338
rect 1152 21264 10560 21286
rect 2896 21175 2902 21227
rect 2954 21215 2960 21227
rect 4243 21218 4301 21224
rect 4243 21215 4255 21218
rect 2954 21187 4255 21215
rect 2954 21175 2960 21187
rect 4243 21184 4255 21187
rect 4289 21215 4301 21218
rect 7408 21215 7414 21227
rect 4289 21187 7414 21215
rect 4289 21184 4301 21187
rect 4243 21178 4301 21184
rect 7408 21175 7414 21187
rect 7466 21175 7472 21227
rect 2227 21070 2285 21076
rect 2227 21036 2239 21070
rect 2273 21067 2285 21070
rect 3760 21067 3766 21079
rect 2273 21039 3766 21067
rect 2273 21036 2285 21039
rect 2227 21030 2285 21036
rect 3760 21027 3766 21039
rect 3818 21027 3824 21079
rect 2608 20953 2614 21005
rect 2666 20953 2672 21005
rect 2704 20953 2710 21005
rect 2762 20993 2768 21005
rect 6931 20996 6989 21002
rect 6931 20993 6943 20996
rect 2762 20965 6943 20993
rect 2762 20953 2768 20965
rect 6931 20962 6943 20965
rect 6977 20962 6989 20996
rect 6931 20956 6989 20962
rect 7312 20953 7318 21005
rect 7370 20953 7376 21005
rect 7894 20931 7946 20937
rect 3472 20879 3478 20931
rect 3530 20879 3536 20931
rect 7894 20873 7946 20879
rect 8947 20774 9005 20780
rect 8947 20740 8959 20774
rect 8993 20771 9005 20774
rect 9712 20771 9718 20783
rect 8993 20743 9718 20771
rect 8993 20740 9005 20743
rect 8947 20734 9005 20740
rect 9712 20731 9718 20743
rect 9770 20731 9776 20783
rect 1152 20672 10560 20694
rect 1152 20620 1966 20672
rect 2018 20620 2030 20672
rect 2082 20620 2094 20672
rect 2146 20620 2158 20672
rect 2210 20620 2222 20672
rect 2274 20620 2286 20672
rect 2338 20620 7966 20672
rect 8018 20620 8030 20672
rect 8082 20620 8094 20672
rect 8146 20620 8158 20672
rect 8210 20620 8222 20672
rect 8274 20620 8286 20672
rect 8338 20620 10560 20672
rect 1152 20598 10560 20620
rect 4240 20361 4246 20413
rect 4298 20401 4304 20413
rect 6739 20404 6797 20410
rect 6739 20401 6751 20404
rect 4298 20373 6751 20401
rect 4298 20361 4304 20373
rect 6739 20370 6751 20373
rect 6785 20370 6797 20404
rect 6739 20364 6797 20370
rect 7888 20361 7894 20413
rect 7946 20361 7952 20413
rect 7123 20330 7181 20336
rect 7123 20296 7135 20330
rect 7169 20296 7181 20330
rect 7123 20290 7181 20296
rect 7138 20253 7166 20290
rect 9808 20287 9814 20339
rect 9866 20287 9872 20339
rect 7312 20253 7318 20265
rect 7138 20225 7318 20253
rect 7312 20213 7318 20225
rect 7370 20213 7376 20265
rect 8755 20182 8813 20188
rect 8755 20148 8767 20182
rect 8801 20179 8813 20182
rect 9328 20179 9334 20191
rect 8801 20151 9334 20179
rect 8801 20148 8813 20151
rect 8755 20142 8813 20148
rect 9328 20139 9334 20151
rect 9386 20139 9392 20191
rect 10096 20139 10102 20191
rect 10154 20139 10160 20191
rect 1152 20006 10560 20028
rect 1152 19954 4966 20006
rect 5018 19954 5030 20006
rect 5082 19954 5094 20006
rect 5146 19954 5158 20006
rect 5210 19954 5222 20006
rect 5274 19954 5286 20006
rect 5338 19954 10560 20006
rect 1152 19932 10560 19954
rect 1744 19695 1750 19747
rect 1802 19735 1808 19747
rect 6931 19738 6989 19744
rect 6931 19735 6943 19738
rect 1802 19707 6943 19735
rect 1802 19695 1808 19707
rect 6931 19704 6943 19707
rect 6977 19704 6989 19738
rect 6931 19698 6989 19704
rect 7312 19621 7318 19673
rect 7370 19621 7376 19673
rect 7894 19599 7946 19605
rect 7894 19541 7946 19547
rect 8947 19442 9005 19448
rect 8947 19408 8959 19442
rect 8993 19439 9005 19442
rect 9904 19439 9910 19451
rect 8993 19411 9910 19439
rect 8993 19408 9005 19411
rect 8947 19402 9005 19408
rect 9904 19399 9910 19411
rect 9962 19399 9968 19451
rect 1152 19340 10560 19362
rect 1152 19288 1966 19340
rect 2018 19288 2030 19340
rect 2082 19288 2094 19340
rect 2146 19288 2158 19340
rect 2210 19288 2222 19340
rect 2274 19288 2286 19340
rect 2338 19288 7966 19340
rect 8018 19288 8030 19340
rect 8082 19288 8094 19340
rect 8146 19288 8158 19340
rect 8210 19288 8222 19340
rect 8274 19288 8286 19340
rect 8338 19288 10560 19340
rect 1152 19266 10560 19288
rect 1648 18881 1654 18933
rect 1706 18881 1712 18933
rect 1747 18776 1805 18782
rect 1747 18742 1759 18776
rect 1793 18773 1805 18776
rect 3664 18773 3670 18785
rect 1793 18745 3670 18773
rect 1793 18742 1805 18745
rect 1747 18736 1805 18742
rect 3664 18733 3670 18745
rect 3722 18733 3728 18785
rect 1152 18674 10560 18696
rect 1152 18622 4966 18674
rect 5018 18622 5030 18674
rect 5082 18622 5094 18674
rect 5146 18622 5158 18674
rect 5210 18622 5222 18674
rect 5274 18622 5286 18674
rect 5338 18622 10560 18674
rect 1152 18600 10560 18622
rect 2803 18554 2861 18560
rect 2803 18520 2815 18554
rect 2849 18551 2861 18554
rect 2896 18551 2902 18563
rect 2849 18523 2902 18551
rect 2849 18520 2861 18523
rect 2803 18514 2861 18520
rect 2896 18511 2902 18523
rect 2954 18551 2960 18563
rect 3376 18551 3382 18563
rect 2954 18523 3382 18551
rect 2954 18511 2960 18523
rect 3376 18511 3382 18523
rect 3434 18511 3440 18563
rect 3280 18363 3286 18415
rect 3338 18403 3344 18415
rect 4240 18403 4246 18415
rect 3338 18375 4246 18403
rect 3338 18363 3344 18375
rect 4240 18363 4246 18375
rect 4298 18403 4304 18415
rect 4819 18406 4877 18412
rect 4819 18403 4831 18406
rect 4298 18375 4831 18403
rect 4298 18363 4304 18375
rect 4819 18372 4831 18375
rect 4865 18372 4877 18406
rect 4819 18366 4877 18372
rect 7504 18363 7510 18415
rect 7562 18363 7568 18415
rect 4144 18289 4150 18341
rect 4202 18329 4208 18341
rect 4435 18332 4493 18338
rect 4435 18329 4447 18332
rect 4202 18301 4447 18329
rect 4202 18289 4208 18301
rect 4435 18298 4447 18301
rect 4481 18298 4493 18332
rect 4435 18292 4493 18298
rect 7312 18289 7318 18341
rect 7370 18329 7376 18341
rect 7888 18329 7894 18341
rect 7370 18301 7894 18329
rect 7370 18289 7376 18301
rect 7888 18289 7894 18301
rect 7946 18289 7952 18341
rect 9523 18332 9581 18338
rect 9523 18298 9535 18332
rect 9569 18329 9581 18332
rect 9811 18332 9869 18338
rect 9811 18329 9823 18332
rect 9569 18301 9823 18329
rect 9569 18298 9581 18301
rect 9523 18292 9581 18298
rect 9811 18298 9823 18301
rect 9857 18298 9869 18332
rect 9811 18292 9869 18298
rect 3472 18215 3478 18267
rect 3530 18215 3536 18267
rect 7792 18215 7798 18267
rect 7850 18215 7856 18267
rect 3490 18181 3518 18215
rect 4048 18181 4054 18193
rect 3490 18153 4054 18181
rect 4048 18141 4054 18153
rect 4106 18141 4112 18193
rect 10096 18067 10102 18119
rect 10154 18067 10160 18119
rect 1152 18008 10560 18030
rect 1152 17956 1966 18008
rect 2018 17956 2030 18008
rect 2082 17956 2094 18008
rect 2146 17956 2158 18008
rect 2210 17956 2222 18008
rect 2274 17956 2286 18008
rect 2338 17956 7966 18008
rect 8018 17956 8030 18008
rect 8082 17956 8094 18008
rect 8146 17956 8158 18008
rect 8210 17956 8222 18008
rect 8274 17956 8286 18008
rect 8338 17956 10560 18008
rect 1152 17934 10560 17956
rect 3568 17845 3574 17897
rect 3626 17845 3632 17897
rect 4240 17845 4246 17897
rect 4298 17885 4304 17897
rect 5779 17888 5837 17894
rect 5779 17885 5791 17888
rect 4298 17857 5791 17885
rect 4298 17845 4304 17857
rect 5779 17854 5791 17857
rect 5825 17854 5837 17888
rect 5779 17848 5837 17854
rect 3094 17749 3146 17755
rect 3586 17737 3614 17845
rect 4054 17749 4106 17755
rect 3856 17737 3862 17749
rect 3586 17709 3862 17737
rect 3856 17697 3862 17709
rect 3914 17697 3920 17749
rect 3094 17691 3146 17697
rect 4054 17691 4106 17697
rect 1939 17666 1997 17672
rect 1939 17632 1951 17666
rect 1985 17663 1997 17666
rect 4144 17663 4150 17675
rect 1985 17635 4150 17663
rect 1985 17632 1997 17635
rect 1939 17626 1997 17632
rect 4144 17623 4150 17635
rect 4202 17663 4208 17675
rect 4243 17666 4301 17672
rect 4243 17663 4255 17666
rect 4202 17635 4255 17663
rect 4202 17623 4208 17635
rect 4243 17632 4255 17635
rect 4289 17632 4301 17666
rect 4243 17626 4301 17632
rect 1555 17592 1613 17598
rect 1555 17558 1567 17592
rect 1601 17589 1613 17592
rect 3088 17589 3094 17601
rect 1601 17561 3094 17589
rect 1601 17558 1613 17561
rect 1555 17552 1613 17558
rect 3088 17549 3094 17561
rect 3146 17549 3152 17601
rect 1152 17342 10560 17364
rect 1152 17290 4966 17342
rect 5018 17290 5030 17342
rect 5082 17290 5094 17342
rect 5146 17290 5158 17342
rect 5210 17290 5222 17342
rect 5274 17290 5286 17342
rect 5338 17290 10560 17342
rect 1152 17268 10560 17290
rect 2992 17179 2998 17231
rect 3050 17219 3056 17231
rect 5779 17222 5837 17228
rect 5779 17219 5791 17222
rect 3050 17191 5791 17219
rect 3050 17179 3056 17191
rect 5779 17188 5791 17191
rect 5825 17219 5837 17222
rect 5825 17191 7454 17219
rect 5825 17188 5837 17191
rect 5779 17182 5837 17188
rect 7426 17080 7454 17191
rect 7411 17074 7469 17080
rect 7411 17040 7423 17074
rect 7457 17040 7469 17074
rect 7411 17034 7469 17040
rect 4147 17000 4205 17006
rect 4147 16966 4159 17000
rect 4193 16997 4205 17000
rect 4624 16997 4630 17009
rect 4193 16969 4630 16997
rect 4193 16966 4205 16969
rect 4147 16960 4205 16966
rect 4624 16957 4630 16969
rect 4682 16997 4688 17009
rect 5392 16997 5398 17009
rect 4682 16969 5398 16997
rect 4682 16957 4688 16969
rect 5392 16957 5398 16969
rect 5450 16957 5456 17009
rect 7795 17000 7853 17006
rect 7795 16966 7807 17000
rect 7841 16997 7853 17000
rect 7888 16997 7894 17009
rect 7841 16969 7894 16997
rect 7841 16966 7853 16969
rect 7795 16960 7853 16966
rect 7888 16957 7894 16969
rect 7946 16957 7952 17009
rect 3958 16935 4010 16941
rect 3760 16883 3766 16935
rect 3818 16883 3824 16935
rect 3958 16877 4010 16883
rect 7606 16935 7658 16941
rect 7606 16877 7658 16883
rect 4432 16735 4438 16787
rect 4490 16775 4496 16787
rect 5680 16775 5686 16787
rect 4490 16747 5686 16775
rect 4490 16735 4496 16747
rect 5680 16735 5686 16747
rect 5738 16775 5744 16787
rect 9232 16775 9238 16787
rect 5738 16747 9238 16775
rect 5738 16735 5744 16747
rect 9232 16735 9238 16747
rect 9290 16735 9296 16787
rect 9427 16778 9485 16784
rect 9427 16744 9439 16778
rect 9473 16775 9485 16778
rect 9616 16775 9622 16787
rect 9473 16747 9622 16775
rect 9473 16744 9485 16747
rect 9427 16738 9485 16744
rect 9616 16735 9622 16747
rect 9674 16735 9680 16787
rect 1152 16676 10560 16698
rect 1152 16624 1966 16676
rect 2018 16624 2030 16676
rect 2082 16624 2094 16676
rect 2146 16624 2158 16676
rect 2210 16624 2222 16676
rect 2274 16624 2286 16676
rect 2338 16624 7966 16676
rect 8018 16624 8030 16676
rect 8082 16624 8094 16676
rect 8146 16624 8158 16676
rect 8210 16624 8222 16676
rect 8274 16624 8286 16676
rect 8338 16624 10560 16676
rect 1152 16602 10560 16624
rect 7888 16513 7894 16565
rect 7946 16553 7952 16565
rect 8179 16556 8237 16562
rect 8179 16553 8191 16556
rect 7946 16525 8191 16553
rect 7946 16513 7952 16525
rect 8179 16522 8191 16525
rect 8225 16522 8237 16556
rect 8179 16516 8237 16522
rect 3088 16479 3094 16491
rect 2818 16451 3094 16479
rect 2818 16417 2846 16451
rect 3088 16439 3094 16451
rect 3146 16479 3152 16491
rect 3952 16479 3958 16491
rect 3146 16451 3958 16479
rect 3146 16439 3152 16451
rect 3952 16439 3958 16451
rect 4010 16479 4016 16491
rect 4010 16451 6302 16479
rect 4010 16439 4016 16451
rect 2800 16365 2806 16417
rect 2858 16365 2864 16417
rect 3664 16365 3670 16417
rect 3722 16365 3728 16417
rect 4066 16391 4094 16451
rect 6274 16391 6302 16451
rect 3184 16291 3190 16343
rect 3242 16331 3248 16343
rect 3283 16334 3341 16340
rect 3283 16331 3295 16334
rect 3242 16303 3295 16331
rect 3242 16291 3248 16303
rect 3283 16300 3295 16303
rect 3329 16300 3341 16334
rect 3283 16294 3341 16300
rect 4243 16334 4301 16340
rect 4243 16300 4255 16334
rect 4289 16331 4301 16334
rect 4432 16331 4438 16343
rect 4289 16303 4438 16331
rect 4289 16300 4301 16303
rect 4243 16294 4301 16300
rect 4432 16291 4438 16303
rect 4490 16291 4496 16343
rect 6451 16334 6509 16340
rect 6451 16331 6463 16334
rect 5314 16303 6463 16331
rect 3760 16217 3766 16269
rect 3818 16257 3824 16269
rect 3859 16260 3917 16266
rect 3859 16257 3871 16260
rect 3818 16229 3871 16257
rect 3818 16217 3824 16229
rect 3859 16226 3871 16229
rect 3905 16226 3917 16260
rect 3859 16220 3917 16226
rect 4144 16217 4150 16269
rect 4202 16257 4208 16269
rect 5314 16257 5342 16303
rect 6451 16300 6463 16303
rect 6497 16300 6509 16334
rect 6451 16294 6509 16300
rect 4202 16229 5342 16257
rect 6067 16260 6125 16266
rect 4202 16217 4208 16229
rect 6067 16226 6079 16260
rect 6113 16257 6125 16260
rect 8368 16257 8374 16269
rect 6113 16229 8374 16257
rect 6113 16226 6125 16229
rect 6067 16220 6125 16226
rect 8368 16217 8374 16229
rect 8426 16217 8432 16269
rect 1651 16112 1709 16118
rect 1651 16078 1663 16112
rect 1697 16109 1709 16112
rect 2512 16109 2518 16121
rect 1697 16081 2518 16109
rect 1697 16078 1709 16081
rect 1651 16072 1709 16078
rect 2512 16069 2518 16081
rect 2570 16069 2576 16121
rect 5875 16112 5933 16118
rect 5875 16078 5887 16112
rect 5921 16109 5933 16112
rect 5968 16109 5974 16121
rect 5921 16081 5974 16109
rect 5921 16078 5933 16081
rect 5875 16072 5933 16078
rect 5968 16069 5974 16081
rect 6026 16109 6032 16121
rect 6736 16109 6742 16121
rect 6026 16081 6742 16109
rect 6026 16069 6032 16081
rect 6736 16069 6742 16081
rect 6794 16069 6800 16121
rect 1152 16010 10560 16032
rect 1152 15958 4966 16010
rect 5018 15958 5030 16010
rect 5082 15958 5094 16010
rect 5146 15958 5158 16010
rect 5210 15958 5222 16010
rect 5274 15958 5286 16010
rect 5338 15958 10560 16010
rect 1152 15936 10560 15958
rect 3664 15699 3670 15751
rect 3722 15739 3728 15751
rect 3763 15742 3821 15748
rect 3763 15739 3775 15742
rect 3722 15711 3775 15739
rect 3722 15699 3728 15711
rect 3763 15708 3775 15711
rect 3809 15708 3821 15742
rect 3763 15702 3821 15708
rect 7507 15742 7565 15748
rect 7507 15708 7519 15742
rect 7553 15739 7565 15742
rect 8560 15739 8566 15751
rect 7553 15711 8566 15739
rect 7553 15708 7565 15711
rect 7507 15702 7565 15708
rect 8560 15699 8566 15711
rect 8618 15699 8624 15751
rect 3379 15668 3437 15674
rect 3379 15634 3391 15668
rect 3425 15665 3437 15668
rect 3856 15665 3862 15677
rect 3425 15637 3862 15665
rect 3425 15634 3437 15637
rect 3379 15628 3437 15634
rect 3856 15625 3862 15637
rect 3914 15625 3920 15677
rect 7888 15625 7894 15677
rect 7946 15625 7952 15677
rect 9523 15668 9581 15674
rect 9523 15634 9535 15668
rect 9569 15665 9581 15668
rect 9811 15668 9869 15674
rect 9811 15665 9823 15668
rect 9569 15637 9823 15665
rect 9569 15634 9581 15637
rect 9523 15628 9581 15634
rect 9811 15634 9823 15637
rect 9857 15634 9869 15668
rect 9811 15628 9869 15634
rect 2806 15603 2858 15609
rect 7600 15551 7606 15603
rect 7658 15591 7664 15603
rect 7658 15563 7728 15591
rect 7658 15551 7664 15563
rect 2806 15545 2858 15551
rect 1648 15403 1654 15455
rect 1706 15443 1712 15455
rect 1747 15446 1805 15452
rect 1747 15443 1759 15446
rect 1706 15415 1759 15443
rect 1706 15403 1712 15415
rect 1747 15412 1759 15415
rect 1793 15412 1805 15446
rect 1747 15406 1805 15412
rect 10096 15403 10102 15455
rect 10154 15403 10160 15455
rect 1152 15344 10560 15366
rect 1152 15292 1966 15344
rect 2018 15292 2030 15344
rect 2082 15292 2094 15344
rect 2146 15292 2158 15344
rect 2210 15292 2222 15344
rect 2274 15292 2286 15344
rect 2338 15292 7966 15344
rect 8018 15292 8030 15344
rect 8082 15292 8094 15344
rect 8146 15292 8158 15344
rect 8210 15292 8222 15344
rect 8274 15292 8286 15344
rect 8338 15292 10560 15344
rect 1152 15270 10560 15292
rect 6736 15033 6742 15085
rect 6794 15033 6800 15085
rect 7600 15033 7606 15085
rect 7658 15033 7664 15085
rect 7123 15002 7181 15008
rect 7123 14968 7135 15002
rect 7169 14999 7181 15002
rect 7888 14999 7894 15011
rect 7169 14971 7894 14999
rect 7169 14968 7181 14971
rect 7123 14962 7181 14968
rect 7888 14959 7894 14971
rect 7946 14959 7952 15011
rect 8755 14780 8813 14786
rect 8755 14746 8767 14780
rect 8801 14777 8813 14780
rect 9808 14777 9814 14789
rect 8801 14749 9814 14777
rect 8801 14746 8813 14749
rect 8755 14740 8813 14746
rect 9808 14737 9814 14749
rect 9866 14737 9872 14789
rect 1152 14678 10560 14700
rect 1152 14626 4966 14678
rect 5018 14626 5030 14678
rect 5082 14626 5094 14678
rect 5146 14626 5158 14678
rect 5210 14626 5222 14678
rect 5274 14626 5286 14678
rect 5338 14626 10560 14678
rect 1152 14604 10560 14626
rect 7408 14367 7414 14419
rect 7466 14367 7472 14419
rect 7795 14336 7853 14342
rect 7795 14302 7807 14336
rect 7841 14333 7853 14336
rect 7888 14333 7894 14345
rect 7841 14305 7894 14333
rect 7841 14302 7853 14305
rect 7795 14296 7853 14302
rect 7888 14293 7894 14305
rect 7946 14293 7952 14345
rect 7606 14271 7658 14277
rect 880 14219 886 14271
rect 938 14259 944 14271
rect 1651 14262 1709 14268
rect 1651 14259 1663 14262
rect 938 14231 1663 14259
rect 938 14219 944 14231
rect 1651 14228 1663 14231
rect 1697 14228 1709 14262
rect 1651 14222 1709 14228
rect 1747 14262 1805 14268
rect 1747 14228 1759 14262
rect 1793 14259 1805 14262
rect 3760 14259 3766 14271
rect 1793 14231 3766 14259
rect 1793 14228 1805 14231
rect 1747 14222 1805 14228
rect 3760 14219 3766 14231
rect 3818 14219 3824 14271
rect 5776 14219 5782 14271
rect 5834 14259 5840 14271
rect 5834 14231 7606 14259
rect 5834 14219 5840 14231
rect 7606 14213 7658 14219
rect 9424 14071 9430 14123
rect 9482 14071 9488 14123
rect 1152 14012 10560 14034
rect 1152 13960 1966 14012
rect 2018 13960 2030 14012
rect 2082 13960 2094 14012
rect 2146 13960 2158 14012
rect 2210 13960 2222 14012
rect 2274 13960 2286 14012
rect 2338 13960 7966 14012
rect 8018 13960 8030 14012
rect 8082 13960 8094 14012
rect 8146 13960 8158 14012
rect 8210 13960 8222 14012
rect 8274 13960 8286 14012
rect 8338 13960 10560 14012
rect 1152 13938 10560 13960
rect 9808 13627 9814 13679
rect 9866 13627 9872 13679
rect 10096 13405 10102 13457
rect 10154 13405 10160 13457
rect 1152 13346 10560 13368
rect 1152 13294 4966 13346
rect 5018 13294 5030 13346
rect 5082 13294 5094 13346
rect 5146 13294 5158 13346
rect 5210 13294 5222 13346
rect 5274 13294 5286 13346
rect 5338 13294 10560 13346
rect 1152 13272 10560 13294
rect 4624 13183 4630 13235
rect 4682 13223 4688 13235
rect 4723 13226 4781 13232
rect 4723 13223 4735 13226
rect 4682 13195 4735 13223
rect 4682 13183 4688 13195
rect 4723 13192 4735 13195
rect 4769 13192 4781 13226
rect 4723 13186 4781 13192
rect 2608 13035 2614 13087
rect 2666 13075 2672 13087
rect 2707 13078 2765 13084
rect 2707 13075 2719 13078
rect 2666 13047 2719 13075
rect 2666 13035 2672 13047
rect 2707 13044 2719 13047
rect 2753 13044 2765 13078
rect 2707 13038 2765 13044
rect 3091 13004 3149 13010
rect 3091 12970 3103 13004
rect 3137 13001 3149 13004
rect 4144 13001 4150 13013
rect 3137 12973 4150 13001
rect 3137 12970 3149 12973
rect 3091 12964 3149 12970
rect 4144 12961 4150 12973
rect 4202 12961 4208 13013
rect 2800 12887 2806 12939
rect 2858 12927 2864 12939
rect 2858 12899 2928 12927
rect 2858 12887 2864 12899
rect 1152 12680 10560 12702
rect 1152 12628 1966 12680
rect 2018 12628 2030 12680
rect 2082 12628 2094 12680
rect 2146 12628 2158 12680
rect 2210 12628 2222 12680
rect 2274 12628 2286 12680
rect 2338 12628 7966 12680
rect 8018 12628 8030 12680
rect 8082 12628 8094 12680
rect 8146 12628 8158 12680
rect 8210 12628 8222 12680
rect 8274 12628 8286 12680
rect 8338 12628 10560 12680
rect 1152 12606 10560 12628
rect 5680 12517 5686 12569
rect 5738 12557 5744 12569
rect 7027 12560 7085 12566
rect 7027 12557 7039 12560
rect 5738 12529 7039 12557
rect 5738 12517 5744 12529
rect 7027 12526 7039 12529
rect 7073 12526 7085 12560
rect 7027 12520 7085 12526
rect 2800 12369 2806 12421
rect 2858 12369 2864 12421
rect 4624 12369 4630 12421
rect 4682 12409 4688 12421
rect 5107 12412 5165 12418
rect 5107 12409 5119 12412
rect 4682 12381 5119 12409
rect 4682 12369 4688 12381
rect 5107 12378 5119 12381
rect 5153 12378 5165 12412
rect 7504 12409 7510 12421
rect 6672 12381 7510 12409
rect 5107 12372 5165 12378
rect 7504 12369 7510 12381
rect 7562 12369 7568 12421
rect 1939 12338 1997 12344
rect 1939 12304 1951 12338
rect 1985 12335 1997 12338
rect 2992 12335 2998 12347
rect 1985 12307 2998 12335
rect 1985 12304 1997 12307
rect 1939 12298 1997 12304
rect 2992 12295 2998 12307
rect 3050 12295 3056 12347
rect 4144 12295 4150 12347
rect 4202 12335 4208 12347
rect 5491 12338 5549 12344
rect 5491 12335 5503 12338
rect 4202 12307 5503 12335
rect 4202 12295 4208 12307
rect 5491 12304 5503 12307
rect 5537 12304 5549 12338
rect 5491 12298 5549 12304
rect 1555 12264 1613 12270
rect 1555 12230 1567 12264
rect 1601 12261 1613 12264
rect 3664 12261 3670 12273
rect 1601 12233 3670 12261
rect 1601 12230 1613 12233
rect 1555 12224 1613 12230
rect 3664 12221 3670 12233
rect 3722 12221 3728 12273
rect 3184 12073 3190 12125
rect 3242 12113 3248 12125
rect 3571 12116 3629 12122
rect 3571 12113 3583 12116
rect 3242 12085 3583 12113
rect 3242 12073 3248 12085
rect 3571 12082 3583 12085
rect 3617 12082 3629 12116
rect 3571 12076 3629 12082
rect 1152 12014 10560 12036
rect 1152 11962 4966 12014
rect 5018 11962 5030 12014
rect 5082 11962 5094 12014
rect 5146 11962 5158 12014
rect 5210 11962 5222 12014
rect 5274 11962 5286 12014
rect 5338 11962 10560 12014
rect 1152 11940 10560 11962
rect 2608 11851 2614 11903
rect 2666 11851 2672 11903
rect 8464 11851 8470 11903
rect 8522 11851 8528 11903
rect 2992 11703 2998 11755
rect 3050 11743 3056 11755
rect 4627 11746 4685 11752
rect 4627 11743 4639 11746
rect 3050 11715 4639 11743
rect 3050 11703 3056 11715
rect 4627 11712 4639 11715
rect 4673 11712 4685 11746
rect 4627 11706 4685 11712
rect 5680 11703 5686 11755
rect 5738 11743 5744 11755
rect 6451 11746 6509 11752
rect 6451 11743 6463 11746
rect 5738 11715 6463 11743
rect 5738 11703 5744 11715
rect 6451 11712 6463 11715
rect 6497 11712 6509 11746
rect 6451 11706 6509 11712
rect 4144 11629 4150 11681
rect 4202 11669 4208 11681
rect 4243 11672 4301 11678
rect 4243 11669 4255 11672
rect 4202 11641 4255 11669
rect 4202 11629 4208 11641
rect 4243 11638 4255 11641
rect 4289 11669 4301 11672
rect 6835 11672 6893 11678
rect 6835 11669 6847 11672
rect 4289 11641 6847 11669
rect 4289 11638 4301 11641
rect 4243 11632 4301 11638
rect 6835 11638 6847 11641
rect 6881 11669 6893 11672
rect 7120 11669 7126 11681
rect 6881 11641 7126 11669
rect 6881 11638 6893 11641
rect 6835 11632 6893 11638
rect 7120 11629 7126 11641
rect 7178 11629 7184 11681
rect 2800 11481 2806 11533
rect 2858 11521 2864 11533
rect 4450 11521 4478 11581
rect 7504 11555 7510 11607
rect 7562 11555 7568 11607
rect 6064 11521 6070 11533
rect 2858 11493 6070 11521
rect 2858 11481 2864 11493
rect 6064 11481 6070 11493
rect 6122 11481 6128 11533
rect 1152 11348 10560 11370
rect 1152 11296 1966 11348
rect 2018 11296 2030 11348
rect 2082 11296 2094 11348
rect 2146 11296 2158 11348
rect 2210 11296 2222 11348
rect 2274 11296 2286 11348
rect 2338 11296 7966 11348
rect 8018 11296 8030 11348
rect 8082 11296 8094 11348
rect 8146 11296 8158 11348
rect 8210 11296 8222 11348
rect 8274 11296 8286 11348
rect 8338 11296 10560 11348
rect 1152 11274 10560 11296
rect 6064 11185 6070 11237
rect 6122 11225 6128 11237
rect 7504 11225 7510 11237
rect 6122 11197 7510 11225
rect 6122 11185 6128 11197
rect 7504 11185 7510 11197
rect 7562 11185 7568 11237
rect 8368 11185 8374 11237
rect 8426 11225 8432 11237
rect 8659 11228 8717 11234
rect 8659 11225 8671 11228
rect 8426 11197 8671 11225
rect 8426 11185 8432 11197
rect 8659 11194 8671 11197
rect 8705 11194 8717 11228
rect 8659 11188 8717 11194
rect 2800 11037 2806 11089
rect 2858 11037 2864 11089
rect 3664 11037 3670 11089
rect 3722 11077 3728 11089
rect 4531 11080 4589 11086
rect 4531 11077 4543 11080
rect 3722 11049 4543 11077
rect 3722 11037 3728 11049
rect 4531 11046 4543 11049
rect 4577 11046 4589 11080
rect 6082 11063 6110 11185
rect 6832 11151 6838 11163
rect 6754 11123 6838 11151
rect 6754 11086 6782 11123
rect 6832 11111 6838 11123
rect 6890 11151 6896 11163
rect 8176 11151 8182 11163
rect 6890 11123 8182 11151
rect 6890 11111 6896 11123
rect 8176 11111 8182 11123
rect 8234 11111 8240 11163
rect 6739 11080 6797 11086
rect 4531 11040 4589 11046
rect 6739 11046 6751 11080
rect 6785 11046 6797 11080
rect 6739 11040 6797 11046
rect 7504 11037 7510 11089
rect 7562 11037 7568 11089
rect 1939 11006 1997 11012
rect 1939 10972 1951 11006
rect 1985 11003 1997 11006
rect 2608 11003 2614 11015
rect 1985 10975 2614 11003
rect 1985 10972 1997 10975
rect 1939 10966 1997 10972
rect 2608 10963 2614 10975
rect 2666 10963 2672 11015
rect 4915 11006 4973 11012
rect 4915 10972 4927 11006
rect 4961 11003 4973 11006
rect 5680 11003 5686 11015
rect 4961 10975 5686 11003
rect 4961 10972 4973 10975
rect 4915 10966 4973 10972
rect 5680 10963 5686 10975
rect 5738 10963 5744 11015
rect 7120 10963 7126 11015
rect 7178 10963 7184 11015
rect 9616 10963 9622 11015
rect 9674 11003 9680 11015
rect 9811 11006 9869 11012
rect 9811 11003 9823 11006
rect 9674 10975 9823 11003
rect 9674 10963 9680 10975
rect 9811 10972 9823 10975
rect 9857 10972 9869 11006
rect 9811 10966 9869 10972
rect 1555 10932 1613 10938
rect 1555 10898 1567 10932
rect 1601 10929 1613 10932
rect 3664 10929 3670 10941
rect 1601 10901 3670 10929
rect 1601 10898 1613 10901
rect 1555 10892 1613 10898
rect 3664 10889 3670 10901
rect 3722 10889 3728 10941
rect 3571 10784 3629 10790
rect 3571 10750 3583 10784
rect 3617 10781 3629 10784
rect 4528 10781 4534 10793
rect 3617 10753 4534 10781
rect 3617 10750 3629 10753
rect 3571 10744 3629 10750
rect 4528 10741 4534 10753
rect 4586 10741 4592 10793
rect 6544 10741 6550 10793
rect 6602 10741 6608 10793
rect 10096 10741 10102 10793
rect 10154 10741 10160 10793
rect 1152 10682 10560 10704
rect 1152 10630 4966 10682
rect 5018 10630 5030 10682
rect 5082 10630 5094 10682
rect 5146 10630 5158 10682
rect 5210 10630 5222 10682
rect 5274 10630 5286 10682
rect 5338 10630 10560 10682
rect 1152 10608 10560 10630
rect 1939 10562 1997 10568
rect 1939 10528 1951 10562
rect 1985 10559 1997 10562
rect 4144 10559 4150 10571
rect 1985 10531 4150 10559
rect 1985 10528 1997 10531
rect 1939 10522 1997 10528
rect 4144 10519 4150 10531
rect 4202 10519 4208 10571
rect 7792 10519 7798 10571
rect 7850 10559 7856 10571
rect 8176 10559 8182 10571
rect 7850 10531 8182 10559
rect 7850 10519 7856 10531
rect 8176 10519 8182 10531
rect 8234 10559 8240 10571
rect 8659 10562 8717 10568
rect 8659 10559 8671 10562
rect 8234 10531 8671 10559
rect 8234 10519 8240 10531
rect 8659 10528 8671 10531
rect 8705 10528 8717 10562
rect 8659 10522 8717 10528
rect 880 10371 886 10423
rect 938 10411 944 10423
rect 1651 10414 1709 10420
rect 1651 10411 1663 10414
rect 938 10383 1663 10411
rect 938 10371 944 10383
rect 1651 10380 1663 10383
rect 1697 10380 1709 10414
rect 1651 10374 1709 10380
rect 3379 10414 3437 10420
rect 3379 10380 3391 10414
rect 3425 10411 3437 10414
rect 3664 10411 3670 10423
rect 3425 10383 3670 10411
rect 3425 10380 3437 10383
rect 3379 10374 3437 10380
rect 3664 10371 3670 10383
rect 3722 10411 3728 10423
rect 5872 10411 5878 10423
rect 3722 10383 5878 10411
rect 3722 10371 3728 10383
rect 5872 10371 5878 10383
rect 5930 10371 5936 10423
rect 6640 10371 6646 10423
rect 6698 10371 6704 10423
rect 3763 10340 3821 10346
rect 3763 10306 3775 10340
rect 3809 10337 3821 10340
rect 4624 10337 4630 10349
rect 3809 10309 4630 10337
rect 3809 10306 3821 10309
rect 3763 10300 3821 10306
rect 4624 10297 4630 10309
rect 4682 10297 4688 10349
rect 7027 10340 7085 10346
rect 7027 10306 7039 10340
rect 7073 10337 7085 10340
rect 7120 10337 7126 10349
rect 7073 10309 7126 10337
rect 7073 10306 7085 10309
rect 7027 10300 7085 10306
rect 7120 10297 7126 10309
rect 7178 10297 7184 10349
rect 4930 10189 4958 10249
rect 7522 10201 7550 10249
rect 7504 10189 7510 10201
rect 4930 10161 7510 10189
rect 7504 10149 7510 10161
rect 7562 10149 7568 10201
rect 5395 10118 5453 10124
rect 5395 10084 5407 10118
rect 5441 10115 5453 10118
rect 5584 10115 5590 10127
rect 5441 10087 5590 10115
rect 5441 10084 5453 10087
rect 5395 10078 5453 10084
rect 5584 10075 5590 10087
rect 5642 10075 5648 10127
rect 1152 10016 10560 10038
rect 1152 9964 1966 10016
rect 2018 9964 2030 10016
rect 2082 9964 2094 10016
rect 2146 9964 2158 10016
rect 2210 9964 2222 10016
rect 2274 9964 2286 10016
rect 2338 9964 7966 10016
rect 8018 9964 8030 10016
rect 8082 9964 8094 10016
rect 8146 9964 8158 10016
rect 8210 9964 8222 10016
rect 8274 9964 8286 10016
rect 8338 9964 10560 10016
rect 1152 9942 10560 9964
rect 6640 9853 6646 9905
rect 6698 9893 6704 9905
rect 7120 9893 7126 9905
rect 6698 9865 7126 9893
rect 6698 9853 6704 9865
rect 7120 9853 7126 9865
rect 7178 9893 7184 9905
rect 8467 9896 8525 9902
rect 8467 9893 8479 9896
rect 7178 9865 8479 9893
rect 7178 9853 7184 9865
rect 8467 9862 8479 9865
rect 8513 9862 8525 9896
rect 8467 9856 8525 9862
rect 7510 9757 7562 9763
rect 7510 9699 7562 9705
rect 6931 9674 6989 9680
rect 6931 9640 6943 9674
rect 6977 9671 6989 9674
rect 7024 9671 7030 9683
rect 6977 9643 7030 9671
rect 6977 9640 6989 9643
rect 6931 9634 6989 9640
rect 7024 9631 7030 9643
rect 7082 9631 7088 9683
rect 6352 9557 6358 9609
rect 6410 9597 6416 9609
rect 6547 9600 6605 9606
rect 6547 9597 6559 9600
rect 6410 9569 6559 9597
rect 6410 9557 6416 9569
rect 6547 9566 6559 9569
rect 6593 9597 6605 9600
rect 8464 9597 8470 9609
rect 6593 9569 8470 9597
rect 6593 9566 6605 9569
rect 6547 9560 6605 9566
rect 8464 9557 8470 9569
rect 8522 9557 8528 9609
rect 1152 9350 10560 9372
rect 1152 9298 4966 9350
rect 5018 9298 5030 9350
rect 5082 9298 5094 9350
rect 5146 9298 5158 9350
rect 5210 9298 5222 9350
rect 5274 9298 5286 9350
rect 5338 9298 10560 9350
rect 1152 9276 10560 9298
rect 8179 9008 8237 9014
rect 8179 8974 8191 9008
rect 8225 9005 8237 9008
rect 8368 9005 8374 9017
rect 8225 8977 8374 9005
rect 8225 8974 8237 8977
rect 8179 8968 8237 8974
rect 8368 8965 8374 8977
rect 8426 8965 8432 9017
rect 5872 8891 5878 8943
rect 5930 8931 5936 8943
rect 6736 8931 6742 8943
rect 5930 8903 6742 8931
rect 5930 8891 5936 8903
rect 6736 8891 6742 8903
rect 6794 8931 6800 8943
rect 7795 8934 7853 8940
rect 7795 8931 7807 8934
rect 6794 8903 7807 8931
rect 6794 8891 6800 8903
rect 7795 8900 7807 8903
rect 7841 8900 7853 8934
rect 7795 8894 7853 8900
rect 7504 8817 7510 8869
rect 7562 8857 7568 8869
rect 8002 8857 8030 8917
rect 7562 8829 8030 8857
rect 7562 8817 7568 8829
rect 9520 8743 9526 8795
rect 9578 8783 9584 8795
rect 9715 8786 9773 8792
rect 9715 8783 9727 8786
rect 9578 8755 9727 8783
rect 9578 8743 9584 8755
rect 9715 8752 9727 8755
rect 9761 8752 9773 8786
rect 9715 8746 9773 8752
rect 1152 8684 10560 8706
rect 1152 8632 1966 8684
rect 2018 8632 2030 8684
rect 2082 8632 2094 8684
rect 2146 8632 2158 8684
rect 2210 8632 2222 8684
rect 2274 8632 2286 8684
rect 2338 8632 7966 8684
rect 8018 8632 8030 8684
rect 8082 8632 8094 8684
rect 8146 8632 8158 8684
rect 8210 8632 8222 8684
rect 8274 8632 8286 8684
rect 8338 8632 10560 8684
rect 1152 8610 10560 8632
rect 1840 8299 1846 8351
rect 1898 8339 1904 8351
rect 1954 8339 1982 8399
rect 6736 8373 6742 8425
rect 6794 8373 6800 8425
rect 7504 8373 7510 8425
rect 7562 8373 7568 8425
rect 1898 8311 1982 8339
rect 3667 8342 3725 8348
rect 1898 8299 1904 8311
rect 3667 8308 3679 8342
rect 3713 8339 3725 8342
rect 4240 8339 4246 8351
rect 3713 8311 4246 8339
rect 3713 8308 3725 8311
rect 3667 8302 3725 8308
rect 4240 8299 4246 8311
rect 4298 8299 4304 8351
rect 7120 8299 7126 8351
rect 7178 8299 7184 8351
rect 9424 8299 9430 8351
rect 9482 8339 9488 8351
rect 9811 8342 9869 8348
rect 9811 8339 9823 8342
rect 9482 8311 9823 8339
rect 9482 8299 9488 8311
rect 9811 8308 9823 8311
rect 9857 8308 9869 8342
rect 9811 8302 9869 8308
rect 10096 8299 10102 8351
rect 10154 8299 10160 8351
rect 8755 8120 8813 8126
rect 8755 8086 8767 8120
rect 8801 8117 8813 8120
rect 9232 8117 9238 8129
rect 8801 8089 9238 8117
rect 8801 8086 8813 8089
rect 8755 8080 8813 8086
rect 9232 8077 9238 8089
rect 9290 8077 9296 8129
rect 1152 8018 10560 8040
rect 1152 7966 4966 8018
rect 5018 7966 5030 8018
rect 5082 7966 5094 8018
rect 5146 7966 5158 8018
rect 5210 7966 5222 8018
rect 5274 7966 5286 8018
rect 5338 7966 10560 8018
rect 1152 7944 10560 7966
rect 2896 7855 2902 7907
rect 2954 7895 2960 7907
rect 3667 7898 3725 7904
rect 3667 7895 3679 7898
rect 2954 7867 3679 7895
rect 2954 7855 2960 7867
rect 3667 7864 3679 7867
rect 3713 7864 3725 7898
rect 3667 7858 3725 7864
rect 1456 7781 1462 7833
rect 1514 7821 1520 7833
rect 1514 7793 3902 7821
rect 1514 7781 1520 7793
rect 3187 7750 3245 7756
rect 3187 7747 3199 7750
rect 2626 7719 3199 7747
rect 2626 7682 2654 7719
rect 3187 7716 3199 7719
rect 3233 7747 3245 7750
rect 3874 7747 3902 7793
rect 4435 7750 4493 7756
rect 4435 7747 4447 7750
rect 3233 7719 3806 7747
rect 3874 7719 4447 7747
rect 3233 7716 3245 7719
rect 3187 7710 3245 7716
rect 2611 7676 2669 7682
rect 2611 7642 2623 7676
rect 2657 7642 2669 7676
rect 2611 7636 2669 7642
rect 2704 7633 2710 7685
rect 2762 7673 2768 7685
rect 2803 7676 2861 7682
rect 2803 7673 2815 7676
rect 2762 7645 2815 7673
rect 2762 7633 2768 7645
rect 2803 7642 2815 7645
rect 2849 7642 2861 7676
rect 2803 7636 2861 7642
rect 2899 7676 2957 7682
rect 2899 7642 2911 7676
rect 2945 7642 2957 7676
rect 2899 7636 2957 7642
rect 3571 7676 3629 7682
rect 3571 7642 3583 7676
rect 3617 7642 3629 7676
rect 3571 7636 3629 7642
rect 1936 7559 1942 7611
rect 1994 7599 2000 7611
rect 2914 7599 2942 7636
rect 3472 7599 3478 7611
rect 1994 7571 3478 7599
rect 1994 7559 2000 7571
rect 3472 7559 3478 7571
rect 3530 7559 3536 7611
rect 2416 7411 2422 7463
rect 2474 7411 2480 7463
rect 2992 7411 2998 7463
rect 3050 7411 3056 7463
rect 3586 7451 3614 7636
rect 3778 7608 3806 7719
rect 4435 7716 4447 7719
rect 4481 7747 4493 7750
rect 5776 7747 5782 7759
rect 4481 7719 5782 7747
rect 4481 7716 4493 7719
rect 4435 7710 4493 7716
rect 5776 7707 5782 7719
rect 5834 7707 5840 7759
rect 6736 7707 6742 7759
rect 6794 7747 6800 7759
rect 7411 7750 7469 7756
rect 7411 7747 7423 7750
rect 6794 7719 7423 7747
rect 6794 7707 6800 7719
rect 7411 7716 7423 7719
rect 7457 7716 7469 7750
rect 7411 7710 7469 7716
rect 3856 7633 3862 7685
rect 3914 7673 3920 7685
rect 3955 7676 4013 7682
rect 3955 7673 3967 7676
rect 3914 7645 3967 7673
rect 3914 7633 3920 7645
rect 3955 7642 3967 7645
rect 4001 7642 4013 7676
rect 3955 7636 4013 7642
rect 7792 7633 7798 7685
rect 7850 7633 7856 7685
rect 3763 7602 3821 7608
rect 3763 7568 3775 7602
rect 3809 7568 3821 7602
rect 3763 7562 3821 7568
rect 7504 7559 7510 7611
rect 7562 7599 7568 7611
rect 7562 7571 7632 7599
rect 7562 7559 7568 7571
rect 4051 7454 4109 7460
rect 4051 7451 4063 7454
rect 3586 7423 4063 7451
rect 4051 7420 4063 7423
rect 4097 7451 4109 7454
rect 4624 7451 4630 7463
rect 4097 7423 4630 7451
rect 4097 7420 4109 7423
rect 4051 7414 4109 7420
rect 4624 7411 4630 7423
rect 4682 7411 4688 7463
rect 9427 7454 9485 7460
rect 9427 7420 9439 7454
rect 9473 7451 9485 7454
rect 9616 7451 9622 7463
rect 9473 7423 9622 7451
rect 9473 7420 9485 7423
rect 9427 7414 9485 7420
rect 9616 7411 9622 7423
rect 9674 7411 9680 7463
rect 1152 7352 10560 7374
rect 1152 7300 1966 7352
rect 2018 7300 2030 7352
rect 2082 7300 2094 7352
rect 2146 7300 2158 7352
rect 2210 7300 2222 7352
rect 2274 7300 2286 7352
rect 2338 7300 7966 7352
rect 8018 7300 8030 7352
rect 8082 7300 8094 7352
rect 8146 7300 8158 7352
rect 8210 7300 8222 7352
rect 8274 7300 8286 7352
rect 8338 7300 10560 7352
rect 1152 7278 10560 7300
rect 3472 7189 3478 7241
rect 3530 7189 3536 7241
rect 4624 7189 4630 7241
rect 4682 7229 4688 7241
rect 7504 7229 7510 7241
rect 4682 7201 7510 7229
rect 4682 7189 4688 7201
rect 7504 7189 7510 7201
rect 7562 7189 7568 7241
rect 2992 7155 2998 7167
rect 1666 7127 2998 7155
rect 1666 7016 1694 7127
rect 2992 7115 2998 7127
rect 3050 7115 3056 7167
rect 4144 7115 4150 7167
rect 4202 7155 4208 7167
rect 4202 7127 5438 7155
rect 4202 7115 4208 7127
rect 2323 7084 2381 7090
rect 2323 7050 2335 7084
rect 2369 7081 2381 7084
rect 2416 7081 2422 7093
rect 2369 7053 2422 7081
rect 2369 7050 2381 7053
rect 2323 7044 2381 7050
rect 2416 7041 2422 7053
rect 2474 7041 2480 7093
rect 2704 7081 2710 7093
rect 2530 7053 2710 7081
rect 1651 7010 1709 7016
rect 1651 6976 1663 7010
rect 1697 6976 1709 7010
rect 1651 6970 1709 6976
rect 1840 6967 1846 7019
rect 1898 7007 1904 7019
rect 1939 7010 1997 7016
rect 1939 7007 1951 7010
rect 1898 6979 1951 7007
rect 1898 6967 1904 6979
rect 1939 6976 1951 6979
rect 1985 7007 1997 7010
rect 2224 7007 2230 7019
rect 1985 6979 2230 7007
rect 1985 6976 1997 6979
rect 1939 6970 1997 6976
rect 2224 6967 2230 6979
rect 2282 6967 2288 7019
rect 1552 6893 1558 6945
rect 1610 6933 1616 6945
rect 2530 6933 2558 7053
rect 2704 7041 2710 7053
rect 2762 7081 2768 7093
rect 2762 7053 5246 7081
rect 2762 7041 2768 7053
rect 4051 7010 4109 7016
rect 4051 6976 4063 7010
rect 4097 6976 4109 7010
rect 4051 6970 4109 6976
rect 1610 6905 2558 6933
rect 4066 6933 4094 6970
rect 4144 6967 4150 7019
rect 4202 6967 4208 7019
rect 4720 6967 4726 7019
rect 4778 6967 4784 7019
rect 5218 7016 5246 7053
rect 5410 7016 5438 7127
rect 7522 7067 7550 7189
rect 5011 7010 5069 7016
rect 5011 6976 5023 7010
rect 5057 6976 5069 7010
rect 5011 6970 5069 6976
rect 5203 7010 5261 7016
rect 5203 6976 5215 7010
rect 5249 6976 5261 7010
rect 5203 6970 5261 6976
rect 5395 7010 5453 7016
rect 5395 6976 5407 7010
rect 5441 6976 5453 7010
rect 5395 6970 5453 6976
rect 4432 6933 4438 6945
rect 4066 6905 4438 6933
rect 1610 6893 1616 6905
rect 4432 6893 4438 6905
rect 4490 6893 4496 6945
rect 4531 6936 4589 6942
rect 4531 6902 4543 6936
rect 4577 6933 4589 6936
rect 4816 6933 4822 6945
rect 4577 6905 4822 6933
rect 4577 6902 4589 6905
rect 4531 6896 4589 6902
rect 4816 6893 4822 6905
rect 4874 6893 4880 6945
rect 2800 6819 2806 6871
rect 2858 6859 2864 6871
rect 5026 6859 5054 6970
rect 5218 6933 5246 6970
rect 6352 6967 6358 7019
rect 6410 6967 6416 7019
rect 5680 6933 5686 6945
rect 5218 6905 5686 6933
rect 5680 6893 5686 6905
rect 5738 6893 5744 6945
rect 5971 6936 6029 6942
rect 5971 6902 5983 6936
rect 6017 6933 6029 6936
rect 6736 6933 6742 6945
rect 6017 6905 6742 6933
rect 6017 6902 6029 6905
rect 5971 6896 6029 6902
rect 6736 6893 6742 6905
rect 6794 6893 6800 6945
rect 2858 6831 5054 6859
rect 2858 6819 2864 6831
rect 1843 6788 1901 6794
rect 1843 6754 1855 6788
rect 1889 6785 1901 6788
rect 3280 6785 3286 6797
rect 1889 6757 3286 6785
rect 1889 6754 1901 6757
rect 1843 6748 1901 6754
rect 3280 6745 3286 6757
rect 3338 6745 3344 6797
rect 3856 6745 3862 6797
rect 3914 6745 3920 6797
rect 3952 6745 3958 6797
rect 4010 6785 4016 6797
rect 4819 6788 4877 6794
rect 4819 6785 4831 6788
rect 4010 6757 4831 6785
rect 4010 6745 4016 6757
rect 4819 6754 4831 6757
rect 4865 6754 4877 6788
rect 4819 6748 4877 6754
rect 5299 6788 5357 6794
rect 5299 6754 5311 6788
rect 5345 6785 5357 6788
rect 5392 6785 5398 6797
rect 5345 6757 5398 6785
rect 5345 6754 5357 6757
rect 5299 6748 5357 6754
rect 5392 6745 5398 6757
rect 5450 6745 5456 6797
rect 7888 6745 7894 6797
rect 7946 6785 7952 6797
rect 7987 6788 8045 6794
rect 7987 6785 7999 6788
rect 7946 6757 7999 6785
rect 7946 6745 7952 6757
rect 7987 6754 7999 6757
rect 8033 6754 8045 6788
rect 7987 6748 8045 6754
rect 1152 6686 10560 6708
rect 1152 6634 4966 6686
rect 5018 6634 5030 6686
rect 5082 6634 5094 6686
rect 5146 6634 5158 6686
rect 5210 6634 5222 6686
rect 5274 6634 5286 6686
rect 5338 6634 10560 6686
rect 1152 6612 10560 6634
rect 1456 6523 1462 6575
rect 1514 6563 1520 6575
rect 1939 6566 1997 6572
rect 1939 6563 1951 6566
rect 1514 6535 1951 6563
rect 1514 6523 1520 6535
rect 1939 6532 1951 6535
rect 1985 6532 1997 6566
rect 1939 6526 1997 6532
rect 2323 6566 2381 6572
rect 2323 6532 2335 6566
rect 2369 6563 2381 6566
rect 2515 6566 2573 6572
rect 2515 6563 2527 6566
rect 2369 6535 2527 6563
rect 2369 6532 2381 6535
rect 2323 6526 2381 6532
rect 2515 6532 2527 6535
rect 2561 6563 2573 6566
rect 2896 6563 2902 6575
rect 2561 6535 2902 6563
rect 2561 6532 2573 6535
rect 2515 6526 2573 6532
rect 2896 6523 2902 6535
rect 2954 6523 2960 6575
rect 4624 6523 4630 6575
rect 4682 6523 4688 6575
rect 2416 6489 2422 6501
rect 1858 6461 2422 6489
rect 1552 6375 1558 6427
rect 1610 6375 1616 6427
rect 1744 6301 1750 6353
rect 1802 6301 1808 6353
rect 1858 6350 1886 6461
rect 2416 6449 2422 6461
rect 2474 6449 2480 6501
rect 2800 6449 2806 6501
rect 2858 6449 2864 6501
rect 5299 6492 5357 6498
rect 5299 6489 5311 6492
rect 3202 6461 5311 6489
rect 2131 6418 2189 6424
rect 2131 6384 2143 6418
rect 2177 6384 2189 6418
rect 2131 6378 2189 6384
rect 2611 6418 2669 6424
rect 2611 6384 2623 6418
rect 2657 6415 2669 6418
rect 3202 6415 3230 6461
rect 5299 6458 5311 6461
rect 5345 6458 5357 6492
rect 5299 6452 5357 6458
rect 5680 6449 5686 6501
rect 5738 6449 5744 6501
rect 2657 6387 3230 6415
rect 2657 6384 2669 6387
rect 2611 6378 2669 6384
rect 1843 6344 1901 6350
rect 1843 6310 1855 6344
rect 1889 6310 1901 6344
rect 1843 6304 1901 6310
rect 2146 6267 2174 6378
rect 3280 6375 3286 6427
rect 3338 6375 3344 6427
rect 4816 6375 4822 6427
rect 4874 6375 4880 6427
rect 5587 6418 5645 6424
rect 5587 6415 5599 6418
rect 4930 6387 5599 6415
rect 2224 6301 2230 6353
rect 2282 6341 2288 6353
rect 2899 6344 2957 6350
rect 2899 6341 2911 6344
rect 2282 6313 2911 6341
rect 2282 6301 2288 6313
rect 2899 6310 2911 6313
rect 2945 6310 2957 6344
rect 2899 6304 2957 6310
rect 3856 6301 3862 6353
rect 3914 6341 3920 6353
rect 4930 6341 4958 6387
rect 5587 6384 5599 6387
rect 5633 6384 5645 6418
rect 5587 6378 5645 6384
rect 5776 6375 5782 6427
rect 5834 6375 5840 6427
rect 3914 6313 4958 6341
rect 3914 6301 3920 6313
rect 5104 6301 5110 6353
rect 5162 6301 5168 6353
rect 9712 6301 9718 6353
rect 9770 6341 9776 6353
rect 9811 6344 9869 6350
rect 9811 6341 9823 6344
rect 9770 6313 9823 6341
rect 9770 6301 9776 6313
rect 9811 6310 9823 6313
rect 9857 6310 9869 6344
rect 9811 6304 9869 6310
rect 2146 6239 2894 6267
rect 1843 6196 1901 6202
rect 1843 6162 1855 6196
rect 1889 6193 1901 6196
rect 2866 6193 2894 6239
rect 3856 6193 3862 6205
rect 1889 6165 2462 6193
rect 2866 6165 3862 6193
rect 1889 6162 1901 6165
rect 1843 6156 1901 6162
rect 2434 6119 2462 6165
rect 3856 6153 3862 6165
rect 3914 6153 3920 6205
rect 4240 6119 4246 6131
rect 2434 6091 4246 6119
rect 4240 6079 4246 6091
rect 4298 6079 4304 6131
rect 4432 6079 4438 6131
rect 4490 6119 4496 6131
rect 5488 6119 5494 6131
rect 4490 6091 5494 6119
rect 4490 6079 4496 6091
rect 5488 6079 5494 6091
rect 5546 6079 5552 6131
rect 10096 6079 10102 6131
rect 10154 6079 10160 6131
rect 1152 6020 10560 6042
rect 1152 5968 1966 6020
rect 2018 5968 2030 6020
rect 2082 5968 2094 6020
rect 2146 5968 2158 6020
rect 2210 5968 2222 6020
rect 2274 5968 2286 6020
rect 2338 5968 7966 6020
rect 8018 5968 8030 6020
rect 8082 5968 8094 6020
rect 8146 5968 8158 6020
rect 8210 5968 8222 6020
rect 8274 5968 8286 6020
rect 8338 5968 10560 6020
rect 1152 5946 10560 5968
rect 5104 5857 5110 5909
rect 5162 5897 5168 5909
rect 5779 5900 5837 5906
rect 5779 5897 5791 5900
rect 5162 5869 5791 5897
rect 5162 5857 5168 5869
rect 5779 5866 5791 5869
rect 5825 5866 5837 5900
rect 5779 5860 5837 5866
rect 3952 5823 3958 5835
rect 2530 5795 3958 5823
rect 2530 5758 2558 5795
rect 3952 5783 3958 5795
rect 4010 5783 4016 5835
rect 2515 5752 2573 5758
rect 2515 5718 2527 5752
rect 2561 5718 2573 5752
rect 2515 5712 2573 5718
rect 4528 5709 4534 5761
rect 4586 5709 4592 5761
rect 5872 5709 5878 5761
rect 5930 5749 5936 5761
rect 5930 5721 6686 5749
rect 5930 5709 5936 5721
rect 1744 5635 1750 5687
rect 1802 5635 1808 5687
rect 1840 5635 1846 5687
rect 1898 5675 1904 5687
rect 2131 5678 2189 5684
rect 2131 5675 2143 5678
rect 1898 5647 2143 5675
rect 1898 5635 1904 5647
rect 2131 5644 2143 5647
rect 2177 5644 2189 5678
rect 2131 5638 2189 5644
rect 3856 5635 3862 5687
rect 3914 5635 3920 5687
rect 5680 5635 5686 5687
rect 5738 5675 5744 5687
rect 5971 5678 6029 5684
rect 5971 5675 5983 5678
rect 5738 5647 5983 5675
rect 5738 5635 5744 5647
rect 5971 5644 5983 5647
rect 6017 5675 6029 5678
rect 6547 5678 6605 5684
rect 6017 5647 6398 5675
rect 6017 5644 6029 5647
rect 5971 5638 6029 5644
rect 5872 5561 5878 5613
rect 5930 5601 5936 5613
rect 6370 5610 6398 5647
rect 6547 5644 6559 5678
rect 6593 5644 6605 5678
rect 6547 5638 6605 5644
rect 6067 5604 6125 5610
rect 6067 5601 6079 5604
rect 5930 5573 6079 5601
rect 5930 5561 5936 5573
rect 6067 5570 6079 5573
rect 6113 5570 6125 5604
rect 6067 5564 6125 5570
rect 6355 5604 6413 5610
rect 6355 5570 6367 5604
rect 6401 5570 6413 5604
rect 6355 5564 6413 5570
rect 2416 5487 2422 5539
rect 2474 5527 2480 5539
rect 6451 5530 6509 5536
rect 6451 5527 6463 5530
rect 2474 5499 6463 5527
rect 2474 5487 2480 5499
rect 6451 5496 6463 5499
rect 6497 5496 6509 5530
rect 6451 5490 6509 5496
rect 2035 5456 2093 5462
rect 2035 5422 2047 5456
rect 2081 5453 2093 5456
rect 3568 5453 3574 5465
rect 2081 5425 3574 5453
rect 2081 5422 2093 5425
rect 2035 5416 2093 5422
rect 3568 5413 3574 5425
rect 3626 5413 3632 5465
rect 3667 5456 3725 5462
rect 3667 5422 3679 5456
rect 3713 5453 3725 5456
rect 4816 5453 4822 5465
rect 3713 5425 4822 5453
rect 3713 5422 3725 5425
rect 3667 5416 3725 5422
rect 4816 5413 4822 5425
rect 4874 5413 4880 5465
rect 5488 5413 5494 5465
rect 5546 5453 5552 5465
rect 6067 5456 6125 5462
rect 6067 5453 6079 5456
rect 5546 5425 6079 5453
rect 5546 5413 5552 5425
rect 6067 5422 6079 5425
rect 6113 5453 6125 5456
rect 6562 5453 6590 5638
rect 6658 5610 6686 5721
rect 6643 5604 6701 5610
rect 6643 5570 6655 5604
rect 6689 5570 6701 5604
rect 6643 5564 6701 5570
rect 6113 5425 6590 5453
rect 6113 5422 6125 5425
rect 6067 5416 6125 5422
rect 1152 5354 10560 5376
rect 1152 5302 4966 5354
rect 5018 5302 5030 5354
rect 5082 5302 5094 5354
rect 5146 5302 5158 5354
rect 5210 5302 5222 5354
rect 5274 5302 5286 5354
rect 5338 5302 10560 5354
rect 1152 5280 10560 5302
rect 4720 5191 4726 5243
rect 4778 5231 4784 5243
rect 5395 5234 5453 5240
rect 5395 5231 5407 5234
rect 4778 5203 5407 5231
rect 4778 5191 4784 5203
rect 5395 5200 5407 5203
rect 5441 5231 5453 5234
rect 5680 5231 5686 5243
rect 5441 5203 5686 5231
rect 5441 5200 5453 5203
rect 5395 5194 5453 5200
rect 5680 5191 5686 5203
rect 5738 5191 5744 5243
rect 5776 5191 5782 5243
rect 5834 5231 5840 5243
rect 6739 5234 6797 5240
rect 6739 5231 6751 5234
rect 5834 5203 6751 5231
rect 5834 5191 5840 5203
rect 6739 5200 6751 5203
rect 6785 5200 6797 5234
rect 6739 5194 6797 5200
rect 2227 5160 2285 5166
rect 2227 5126 2239 5160
rect 2273 5157 2285 5160
rect 4144 5157 4150 5169
rect 2273 5129 4150 5157
rect 2273 5126 2285 5129
rect 2227 5120 2285 5126
rect 4144 5117 4150 5129
rect 4202 5157 4208 5169
rect 5872 5157 5878 5169
rect 4202 5129 5878 5157
rect 4202 5117 4208 5129
rect 4240 5043 4246 5095
rect 4298 5043 4304 5095
rect 5488 5043 5494 5095
rect 5546 5043 5552 5095
rect 3763 5012 3821 5018
rect 3763 4978 3775 5012
rect 3809 5009 3821 5012
rect 3856 5009 3862 5021
rect 3809 4981 3862 5009
rect 3809 4978 3821 4981
rect 3763 4972 3821 4978
rect 3856 4969 3862 4981
rect 3914 4969 3920 5021
rect 5794 5018 5822 5129
rect 5872 5117 5878 5129
rect 5930 5117 5936 5169
rect 5971 5160 6029 5166
rect 5971 5126 5983 5160
rect 6017 5157 6029 5160
rect 6017 5129 6686 5157
rect 6017 5126 6029 5129
rect 5971 5120 6029 5126
rect 6658 5092 6686 5129
rect 6643 5086 6701 5092
rect 6643 5052 6655 5086
rect 6689 5052 6701 5086
rect 6643 5046 6701 5052
rect 5779 5012 5837 5018
rect 5779 4978 5791 5012
rect 5825 4978 5837 5012
rect 5779 4972 5837 4978
rect 3379 4938 3437 4944
rect 3379 4904 3391 4938
rect 3425 4935 3437 4938
rect 5392 4935 5398 4947
rect 3425 4907 5398 4935
rect 3425 4904 3437 4907
rect 3379 4898 3437 4904
rect 5392 4895 5398 4907
rect 5450 4895 5456 4947
rect 1744 4821 1750 4873
rect 1802 4861 1808 4873
rect 6451 4864 6509 4870
rect 6451 4861 6463 4864
rect 1802 4833 6463 4861
rect 1802 4821 1808 4833
rect 6451 4830 6463 4833
rect 6497 4830 6509 4864
rect 6451 4824 6509 4830
rect 1152 4688 10560 4710
rect 1152 4636 1966 4688
rect 2018 4636 2030 4688
rect 2082 4636 2094 4688
rect 2146 4636 2158 4688
rect 2210 4636 2222 4688
rect 2274 4636 2286 4688
rect 2338 4636 7966 4688
rect 8018 4636 8030 4688
rect 8082 4636 8094 4688
rect 8146 4636 8158 4688
rect 8210 4636 8222 4688
rect 8274 4636 8286 4688
rect 8338 4636 10560 4688
rect 1152 4614 10560 4636
rect 3856 4377 3862 4429
rect 3914 4417 3920 4429
rect 3914 4389 5040 4417
rect 3914 4377 3920 4389
rect 1648 4303 1654 4355
rect 1706 4343 1712 4355
rect 1747 4346 1805 4352
rect 1747 4343 1759 4346
rect 1706 4315 1759 4343
rect 1706 4303 1712 4315
rect 1747 4312 1759 4315
rect 1793 4312 1805 4346
rect 1747 4306 1805 4312
rect 4528 4303 4534 4355
rect 4586 4303 4592 4355
rect 592 4081 598 4133
rect 650 4121 656 4133
rect 1555 4124 1613 4130
rect 1555 4121 1567 4124
rect 650 4093 1567 4121
rect 650 4081 656 4093
rect 1555 4090 1567 4093
rect 1601 4090 1613 4124
rect 1555 4084 1613 4090
rect 1152 4022 10560 4044
rect 1152 3970 4966 4022
rect 5018 3970 5030 4022
rect 5082 3970 5094 4022
rect 5146 3970 5158 4022
rect 5210 3970 5222 4022
rect 5274 3970 5286 4022
rect 5338 3970 10560 4022
rect 1152 3948 10560 3970
rect 5395 3902 5453 3908
rect 5395 3868 5407 3902
rect 5441 3899 5453 3902
rect 5488 3899 5494 3911
rect 5441 3871 5494 3899
rect 5441 3868 5453 3871
rect 5395 3862 5453 3868
rect 5488 3859 5494 3871
rect 5546 3859 5552 3911
rect 3568 3711 3574 3763
rect 3626 3751 3632 3763
rect 4243 3754 4301 3760
rect 4243 3751 4255 3754
rect 3626 3723 4255 3751
rect 3626 3711 3632 3723
rect 4243 3720 4255 3723
rect 4289 3720 4301 3754
rect 4243 3714 4301 3720
rect 2131 3680 2189 3686
rect 2131 3646 2143 3680
rect 2177 3677 2189 3680
rect 2512 3677 2518 3689
rect 2177 3649 2518 3677
rect 2177 3646 2189 3649
rect 2131 3640 2189 3646
rect 2512 3637 2518 3649
rect 2570 3637 2576 3689
rect 3856 3637 3862 3689
rect 3914 3637 3920 3689
rect 9520 3637 9526 3689
rect 9578 3637 9584 3689
rect 9904 3637 9910 3689
rect 9962 3637 9968 3689
rect 10096 3563 10102 3615
rect 10154 3563 10160 3615
rect 1840 3415 1846 3467
rect 1898 3415 1904 3467
rect 9715 3458 9773 3464
rect 9715 3424 9727 3458
rect 9761 3455 9773 3458
rect 10960 3455 10966 3467
rect 9761 3427 10966 3455
rect 9761 3424 9773 3427
rect 9715 3418 9773 3424
rect 10960 3415 10966 3427
rect 11018 3415 11024 3467
rect 1152 3356 10560 3378
rect 1152 3304 1966 3356
rect 2018 3304 2030 3356
rect 2082 3304 2094 3356
rect 2146 3304 2158 3356
rect 2210 3304 2222 3356
rect 2274 3304 2286 3356
rect 2338 3304 7966 3356
rect 8018 3304 8030 3356
rect 8082 3304 8094 3356
rect 8146 3304 8158 3356
rect 8210 3304 8222 3356
rect 8274 3304 8286 3356
rect 8338 3304 10560 3356
rect 1152 3282 10560 3304
rect 1456 3193 1462 3245
rect 1514 3233 1520 3245
rect 1939 3236 1997 3242
rect 1939 3233 1951 3236
rect 1514 3205 1951 3233
rect 1514 3193 1520 3205
rect 1939 3202 1951 3205
rect 1985 3202 1997 3236
rect 1939 3196 1997 3202
rect 1552 2971 1558 3023
rect 1610 2971 1616 3023
rect 3184 2971 3190 3023
rect 3242 2971 3248 3023
rect 4435 3014 4493 3020
rect 4435 2980 4447 3014
rect 4481 3011 4493 3014
rect 4624 3011 4630 3023
rect 4481 2983 4630 3011
rect 4481 2980 4493 2983
rect 4435 2974 4493 2980
rect 4624 2971 4630 2983
rect 4682 2971 4688 3023
rect 5584 2971 5590 3023
rect 5642 2971 5648 3023
rect 6544 2971 6550 3023
rect 6602 3011 6608 3023
rect 6643 3014 6701 3020
rect 6643 3011 6655 3014
rect 6602 2983 6655 3011
rect 6602 2971 6608 2983
rect 6643 2980 6655 2983
rect 6689 2980 6701 3014
rect 6643 2974 6701 2980
rect 7888 2971 7894 3023
rect 7946 2971 7952 3023
rect 9232 2971 9238 3023
rect 9290 2971 9296 3023
rect 9328 2971 9334 3023
rect 9386 3011 9392 3023
rect 9427 3014 9485 3020
rect 9427 3011 9439 3014
rect 9386 2983 9439 3011
rect 9386 2971 9392 2983
rect 9427 2980 9439 2983
rect 9473 2980 9485 3014
rect 9427 2974 9485 2980
rect 9616 2971 9622 3023
rect 9674 3011 9680 3023
rect 10003 3014 10061 3020
rect 10003 3011 10015 3014
rect 9674 2983 10015 3011
rect 9674 2971 9680 2983
rect 10003 2980 10015 2983
rect 10049 2980 10061 3014
rect 10003 2974 10061 2980
rect 2896 2897 2902 2949
rect 2954 2937 2960 2949
rect 2995 2940 3053 2946
rect 2995 2937 3007 2940
rect 2954 2909 3007 2937
rect 2954 2897 2960 2909
rect 2995 2906 3007 2909
rect 3041 2906 3053 2940
rect 2995 2900 3053 2906
rect 4048 2897 4054 2949
rect 4106 2937 4112 2949
rect 4147 2940 4205 2946
rect 4147 2937 4159 2940
rect 4106 2909 4159 2937
rect 4106 2897 4112 2909
rect 4147 2906 4159 2909
rect 4193 2906 4205 2940
rect 4147 2900 4205 2906
rect 5299 2940 5357 2946
rect 5299 2906 5311 2940
rect 5345 2937 5357 2940
rect 5392 2937 5398 2949
rect 5345 2909 5398 2937
rect 5345 2906 5357 2909
rect 5299 2900 5357 2906
rect 5392 2897 5398 2909
rect 5450 2897 5456 2949
rect 6352 2897 6358 2949
rect 6410 2937 6416 2949
rect 6451 2940 6509 2946
rect 6451 2937 6463 2940
rect 6410 2909 6463 2937
rect 6410 2897 6416 2909
rect 6451 2906 6463 2909
rect 6497 2906 6509 2940
rect 6451 2900 6509 2906
rect 7600 2897 7606 2949
rect 7658 2897 7664 2949
rect 8656 2897 8662 2949
rect 8714 2937 8720 2949
rect 9043 2940 9101 2946
rect 9043 2937 9055 2940
rect 8714 2909 9055 2937
rect 8714 2897 8720 2909
rect 9043 2906 9055 2909
rect 9089 2906 9101 2940
rect 9043 2900 9101 2906
rect 9712 2897 9718 2949
rect 9770 2897 9776 2949
rect 9808 2897 9814 2949
rect 9866 2897 9872 2949
rect 1152 2690 10560 2712
rect 1152 2638 4966 2690
rect 5018 2638 5030 2690
rect 5082 2638 5094 2690
rect 5146 2638 5158 2690
rect 5210 2638 5222 2690
rect 5274 2638 5286 2690
rect 5338 2638 10560 2690
rect 1152 2616 10560 2638
<< via1 >>
rect 1966 25948 2018 26000
rect 2030 25948 2082 26000
rect 2094 25948 2146 26000
rect 2158 25948 2210 26000
rect 2222 25948 2274 26000
rect 2286 25948 2338 26000
rect 7966 25948 8018 26000
rect 8030 25948 8082 26000
rect 8094 25948 8146 26000
rect 8158 25948 8210 26000
rect 8222 25948 8274 26000
rect 8286 25948 8338 26000
rect 1558 25880 1610 25889
rect 1558 25846 1567 25880
rect 1567 25846 1601 25880
rect 1601 25846 1610 25880
rect 1558 25837 1610 25846
rect 1846 25837 1898 25889
rect 2614 25837 2666 25889
rect 3286 25880 3338 25889
rect 3286 25846 3295 25880
rect 3295 25846 3329 25880
rect 3329 25846 3338 25880
rect 3286 25837 3338 25846
rect 3862 25880 3914 25889
rect 3862 25846 3871 25880
rect 3871 25846 3905 25880
rect 3905 25846 3914 25880
rect 3862 25837 3914 25846
rect 4438 25880 4490 25889
rect 4438 25846 4447 25880
rect 4447 25846 4481 25880
rect 4481 25846 4490 25880
rect 4438 25837 4490 25846
rect 5014 25880 5066 25889
rect 5014 25846 5023 25880
rect 5023 25846 5057 25880
rect 5057 25846 5066 25880
rect 5014 25837 5066 25846
rect 5494 25837 5546 25889
rect 6262 25880 6314 25889
rect 6262 25846 6271 25880
rect 6271 25846 6305 25880
rect 6305 25846 6314 25880
rect 6262 25837 6314 25846
rect 6742 25880 6794 25889
rect 6742 25846 6751 25880
rect 6751 25846 6785 25880
rect 6785 25846 6794 25880
rect 6742 25837 6794 25846
rect 7318 25880 7370 25889
rect 7318 25846 7327 25880
rect 7327 25846 7361 25880
rect 7361 25846 7370 25880
rect 7318 25837 7370 25846
rect 7894 25880 7946 25889
rect 7894 25846 7903 25880
rect 7903 25846 7937 25880
rect 7937 25846 7946 25880
rect 7894 25837 7946 25846
rect 8470 25880 8522 25889
rect 8470 25846 8479 25880
rect 8479 25846 8513 25880
rect 8513 25846 8522 25880
rect 8470 25837 8522 25846
rect 9046 25880 9098 25889
rect 9046 25846 9055 25880
rect 9055 25846 9089 25880
rect 9089 25846 9098 25880
rect 9046 25837 9098 25846
rect 9622 25880 9674 25889
rect 9622 25846 9631 25880
rect 9631 25846 9665 25880
rect 9665 25846 9674 25880
rect 9622 25837 9674 25846
rect 1654 25615 1706 25667
rect 2902 25615 2954 25667
rect 2998 25658 3050 25667
rect 2998 25624 3007 25658
rect 3007 25624 3041 25658
rect 3041 25624 3050 25658
rect 2998 25615 3050 25624
rect 5974 25763 6026 25815
rect 3670 25689 3722 25741
rect 5782 25615 5834 25667
rect 5878 25658 5930 25667
rect 5878 25624 5887 25658
rect 5887 25624 5921 25658
rect 5921 25624 5930 25658
rect 5878 25615 5930 25624
rect 6934 25658 6986 25667
rect 6934 25624 6943 25658
rect 6943 25624 6977 25658
rect 6977 25624 6986 25658
rect 6934 25615 6986 25624
rect 7510 25658 7562 25667
rect 7510 25624 7519 25658
rect 7519 25624 7553 25658
rect 7553 25624 7562 25658
rect 7510 25615 7562 25624
rect 8086 25658 8138 25667
rect 8086 25624 8095 25658
rect 8095 25624 8129 25658
rect 8129 25624 8138 25658
rect 8086 25615 8138 25624
rect 7222 25541 7274 25593
rect 6742 25467 6794 25519
rect 5398 25393 5450 25445
rect 9238 25658 9290 25667
rect 9238 25624 9247 25658
rect 9247 25624 9281 25658
rect 9281 25624 9290 25658
rect 9238 25615 9290 25624
rect 9718 25615 9770 25667
rect 4966 25282 5018 25334
rect 5030 25282 5082 25334
rect 5094 25282 5146 25334
rect 5158 25282 5210 25334
rect 5222 25282 5274 25334
rect 5286 25282 5338 25334
rect 1462 25171 1514 25223
rect 3286 25171 3338 25223
rect 6934 25171 6986 25223
rect 9334 25214 9386 25223
rect 9334 25180 9343 25214
rect 9343 25180 9377 25214
rect 9377 25180 9386 25214
rect 9334 25171 9386 25180
rect 10102 25214 10154 25223
rect 10102 25180 10111 25214
rect 10111 25180 10145 25214
rect 10145 25180 10154 25214
rect 10102 25171 10154 25180
rect 310 25097 362 25149
rect 3382 25097 3434 25149
rect 7510 25097 7562 25149
rect 10678 25097 10730 25149
rect 2614 25023 2666 25075
rect 8086 25023 8138 25075
rect 1846 24992 1898 25001
rect 1846 24958 1855 24992
rect 1855 24958 1889 24992
rect 1889 24958 1898 24992
rect 1846 24949 1898 24958
rect 4246 24949 4298 25001
rect 9334 24949 9386 25001
rect 9430 24992 9482 25001
rect 9430 24958 9439 24992
rect 9439 24958 9473 24992
rect 9473 24958 9482 24992
rect 9430 24949 9482 24958
rect 6838 24875 6890 24927
rect 1966 24616 2018 24668
rect 2030 24616 2082 24668
rect 2094 24616 2146 24668
rect 2158 24616 2210 24668
rect 2222 24616 2274 24668
rect 2286 24616 2338 24668
rect 7966 24616 8018 24668
rect 8030 24616 8082 24668
rect 8094 24616 8146 24668
rect 8158 24616 8210 24668
rect 8222 24616 8274 24668
rect 8286 24616 8338 24668
rect 886 24431 938 24483
rect 6742 24474 6794 24483
rect 6742 24440 6751 24474
rect 6751 24440 6785 24474
rect 6785 24440 6794 24474
rect 6742 24431 6794 24440
rect 11254 24431 11306 24483
rect 6070 24357 6122 24409
rect 9718 24357 9770 24409
rect 1750 24326 1802 24335
rect 1750 24292 1759 24326
rect 1759 24292 1793 24326
rect 1793 24292 1802 24326
rect 1750 24283 1802 24292
rect 7798 24283 7850 24335
rect 8470 24283 8522 24335
rect 4150 24209 4202 24261
rect 6742 24061 6794 24113
rect 8566 24061 8618 24113
rect 4966 23950 5018 24002
rect 5030 23950 5082 24002
rect 5094 23950 5146 24002
rect 5158 23950 5210 24002
rect 5222 23950 5274 24002
rect 5286 23950 5338 24002
rect 5878 23839 5930 23891
rect 4150 23586 4202 23595
rect 4150 23552 4159 23586
rect 4159 23552 4193 23586
rect 4193 23552 4202 23586
rect 4150 23543 4202 23552
rect 6070 23543 6122 23595
rect 8374 23617 8426 23669
rect 7894 23543 7946 23595
rect 8470 23469 8522 23521
rect 9814 23395 9866 23447
rect 1966 23284 2018 23336
rect 2030 23284 2082 23336
rect 2094 23284 2146 23336
rect 2158 23284 2210 23336
rect 2222 23284 2274 23336
rect 2286 23284 2338 23336
rect 7966 23284 8018 23336
rect 8030 23284 8082 23336
rect 8094 23284 8146 23336
rect 8158 23284 8210 23336
rect 8222 23284 8274 23336
rect 8286 23284 8338 23336
rect 3478 23025 3530 23077
rect 6070 23025 6122 23077
rect 3382 22951 3434 23003
rect 3766 22877 3818 22929
rect 4150 22877 4202 22929
rect 5782 22951 5834 23003
rect 7126 22994 7178 23003
rect 7126 22960 7135 22994
rect 7135 22960 7169 22994
rect 7169 22960 7178 22994
rect 7126 22951 7178 22960
rect 6838 22877 6890 22929
rect 1654 22772 1706 22781
rect 1654 22738 1663 22772
rect 1663 22738 1697 22772
rect 1697 22738 1706 22772
rect 1654 22729 1706 22738
rect 2710 22729 2762 22781
rect 6070 22729 6122 22781
rect 8278 22920 8330 22929
rect 8278 22886 8287 22920
rect 8287 22886 8321 22920
rect 8321 22886 8330 22920
rect 8278 22877 8330 22886
rect 9334 22994 9386 23003
rect 9334 22960 9343 22994
rect 9343 22960 9377 22994
rect 9377 22960 9386 22994
rect 9334 22951 9386 22960
rect 9814 22994 9866 23003
rect 9814 22960 9823 22994
rect 9823 22960 9857 22994
rect 9857 22960 9866 22994
rect 9814 22951 9866 22960
rect 9430 22729 9482 22781
rect 10102 22772 10154 22781
rect 10102 22738 10111 22772
rect 10111 22738 10145 22772
rect 10145 22738 10154 22772
rect 10102 22729 10154 22738
rect 4966 22618 5018 22670
rect 5030 22618 5082 22670
rect 5094 22618 5146 22670
rect 5158 22618 5210 22670
rect 5222 22618 5274 22670
rect 5286 22618 5338 22670
rect 1270 22507 1322 22559
rect 4246 22550 4298 22559
rect 4246 22516 4255 22550
rect 4255 22516 4289 22550
rect 4289 22516 4298 22550
rect 4246 22507 4298 22516
rect 7798 22507 7850 22559
rect 8470 22507 8522 22559
rect 3766 22359 3818 22411
rect 7126 22359 7178 22411
rect 3670 22285 3722 22337
rect 7318 22285 7370 22337
rect 8278 22285 8330 22337
rect 3478 22211 3530 22263
rect 7894 22211 7946 22263
rect 9814 22063 9866 22115
rect 1966 21952 2018 22004
rect 2030 21952 2082 22004
rect 2094 21952 2146 22004
rect 2158 21952 2210 22004
rect 2222 21952 2274 22004
rect 2286 21952 2338 22004
rect 7966 21952 8018 22004
rect 8030 21952 8082 22004
rect 8094 21952 8146 22004
rect 8158 21952 8210 22004
rect 8222 21952 8274 22004
rect 8286 21952 8338 22004
rect 7222 21841 7274 21893
rect 7510 21841 7562 21893
rect 1750 21736 1802 21745
rect 1750 21702 1759 21736
rect 1759 21702 1793 21736
rect 1793 21702 1802 21736
rect 1750 21693 1802 21702
rect 3478 21693 3530 21745
rect 6070 21693 6122 21745
rect 3286 21662 3338 21671
rect 3286 21628 3295 21662
rect 3295 21628 3329 21662
rect 3329 21628 3338 21662
rect 3286 21619 3338 21628
rect 3766 21619 3818 21671
rect 6742 21619 6794 21671
rect 4966 21286 5018 21338
rect 5030 21286 5082 21338
rect 5094 21286 5146 21338
rect 5158 21286 5210 21338
rect 5222 21286 5274 21338
rect 5286 21286 5338 21338
rect 2902 21175 2954 21227
rect 7414 21175 7466 21227
rect 3766 21027 3818 21079
rect 2614 20996 2666 21005
rect 2614 20962 2623 20996
rect 2623 20962 2657 20996
rect 2657 20962 2666 20996
rect 2614 20953 2666 20962
rect 2710 20953 2762 21005
rect 7318 20996 7370 21005
rect 7318 20962 7327 20996
rect 7327 20962 7361 20996
rect 7361 20962 7370 20996
rect 7318 20953 7370 20962
rect 3478 20879 3530 20931
rect 7894 20879 7946 20931
rect 9718 20731 9770 20783
rect 1966 20620 2018 20672
rect 2030 20620 2082 20672
rect 2094 20620 2146 20672
rect 2158 20620 2210 20672
rect 2222 20620 2274 20672
rect 2286 20620 2338 20672
rect 7966 20620 8018 20672
rect 8030 20620 8082 20672
rect 8094 20620 8146 20672
rect 8158 20620 8210 20672
rect 8222 20620 8274 20672
rect 8286 20620 8338 20672
rect 4246 20361 4298 20413
rect 7894 20361 7946 20413
rect 9814 20330 9866 20339
rect 9814 20296 9823 20330
rect 9823 20296 9857 20330
rect 9857 20296 9866 20330
rect 9814 20287 9866 20296
rect 7318 20213 7370 20265
rect 9334 20139 9386 20191
rect 10102 20182 10154 20191
rect 10102 20148 10111 20182
rect 10111 20148 10145 20182
rect 10145 20148 10154 20182
rect 10102 20139 10154 20148
rect 4966 19954 5018 20006
rect 5030 19954 5082 20006
rect 5094 19954 5146 20006
rect 5158 19954 5210 20006
rect 5222 19954 5274 20006
rect 5286 19954 5338 20006
rect 1750 19695 1802 19747
rect 7318 19664 7370 19673
rect 7318 19630 7327 19664
rect 7327 19630 7361 19664
rect 7361 19630 7370 19664
rect 7318 19621 7370 19630
rect 7894 19547 7946 19599
rect 9910 19399 9962 19451
rect 1966 19288 2018 19340
rect 2030 19288 2082 19340
rect 2094 19288 2146 19340
rect 2158 19288 2210 19340
rect 2222 19288 2274 19340
rect 2286 19288 2338 19340
rect 7966 19288 8018 19340
rect 8030 19288 8082 19340
rect 8094 19288 8146 19340
rect 8158 19288 8210 19340
rect 8222 19288 8274 19340
rect 8286 19288 8338 19340
rect 1654 18924 1706 18933
rect 1654 18890 1663 18924
rect 1663 18890 1697 18924
rect 1697 18890 1706 18924
rect 1654 18881 1706 18890
rect 3670 18733 3722 18785
rect 4966 18622 5018 18674
rect 5030 18622 5082 18674
rect 5094 18622 5146 18674
rect 5158 18622 5210 18674
rect 5222 18622 5274 18674
rect 5286 18622 5338 18674
rect 2902 18511 2954 18563
rect 3382 18511 3434 18563
rect 3286 18363 3338 18415
rect 4246 18363 4298 18415
rect 7510 18406 7562 18415
rect 7510 18372 7519 18406
rect 7519 18372 7553 18406
rect 7553 18372 7562 18406
rect 7510 18363 7562 18372
rect 4150 18289 4202 18341
rect 7318 18289 7370 18341
rect 7894 18332 7946 18341
rect 7894 18298 7903 18332
rect 7903 18298 7937 18332
rect 7937 18298 7946 18332
rect 7894 18289 7946 18298
rect 3478 18215 3530 18267
rect 7798 18215 7850 18267
rect 4054 18141 4106 18193
rect 10102 18110 10154 18119
rect 10102 18076 10111 18110
rect 10111 18076 10145 18110
rect 10145 18076 10154 18110
rect 10102 18067 10154 18076
rect 1966 17956 2018 18008
rect 2030 17956 2082 18008
rect 2094 17956 2146 18008
rect 2158 17956 2210 18008
rect 2222 17956 2274 18008
rect 2286 17956 2338 18008
rect 7966 17956 8018 18008
rect 8030 17956 8082 18008
rect 8094 17956 8146 18008
rect 8158 17956 8210 18008
rect 8222 17956 8274 18008
rect 8286 17956 8338 18008
rect 3574 17888 3626 17897
rect 3574 17854 3583 17888
rect 3583 17854 3617 17888
rect 3617 17854 3626 17888
rect 3574 17845 3626 17854
rect 4246 17845 4298 17897
rect 3094 17697 3146 17749
rect 3862 17740 3914 17749
rect 3862 17706 3871 17740
rect 3871 17706 3905 17740
rect 3905 17706 3914 17740
rect 3862 17697 3914 17706
rect 4054 17697 4106 17749
rect 4150 17623 4202 17675
rect 3094 17549 3146 17601
rect 4966 17290 5018 17342
rect 5030 17290 5082 17342
rect 5094 17290 5146 17342
rect 5158 17290 5210 17342
rect 5222 17290 5274 17342
rect 5286 17290 5338 17342
rect 2998 17179 3050 17231
rect 4630 16957 4682 17009
rect 5398 16957 5450 17009
rect 7894 16957 7946 17009
rect 3766 16926 3818 16935
rect 3766 16892 3775 16926
rect 3775 16892 3809 16926
rect 3809 16892 3818 16926
rect 3766 16883 3818 16892
rect 3958 16883 4010 16935
rect 7606 16883 7658 16935
rect 4438 16735 4490 16787
rect 5686 16735 5738 16787
rect 9238 16735 9290 16787
rect 9622 16735 9674 16787
rect 1966 16624 2018 16676
rect 2030 16624 2082 16676
rect 2094 16624 2146 16676
rect 2158 16624 2210 16676
rect 2222 16624 2274 16676
rect 2286 16624 2338 16676
rect 7966 16624 8018 16676
rect 8030 16624 8082 16676
rect 8094 16624 8146 16676
rect 8158 16624 8210 16676
rect 8222 16624 8274 16676
rect 8286 16624 8338 16676
rect 7894 16513 7946 16565
rect 3094 16439 3146 16491
rect 3958 16439 4010 16491
rect 2806 16365 2858 16417
rect 3670 16408 3722 16417
rect 3670 16374 3679 16408
rect 3679 16374 3713 16408
rect 3713 16374 3722 16408
rect 3670 16365 3722 16374
rect 3190 16291 3242 16343
rect 4438 16291 4490 16343
rect 3766 16217 3818 16269
rect 4150 16217 4202 16269
rect 8374 16217 8426 16269
rect 2518 16069 2570 16121
rect 5974 16069 6026 16121
rect 6742 16069 6794 16121
rect 4966 15958 5018 16010
rect 5030 15958 5082 16010
rect 5094 15958 5146 16010
rect 5158 15958 5210 16010
rect 5222 15958 5274 16010
rect 5286 15958 5338 16010
rect 3670 15699 3722 15751
rect 8566 15699 8618 15751
rect 3862 15625 3914 15677
rect 7894 15668 7946 15677
rect 7894 15634 7903 15668
rect 7903 15634 7937 15668
rect 7937 15634 7946 15668
rect 7894 15625 7946 15634
rect 2806 15551 2858 15603
rect 7606 15551 7658 15603
rect 1654 15403 1706 15455
rect 10102 15446 10154 15455
rect 10102 15412 10111 15446
rect 10111 15412 10145 15446
rect 10145 15412 10154 15446
rect 10102 15403 10154 15412
rect 1966 15292 2018 15344
rect 2030 15292 2082 15344
rect 2094 15292 2146 15344
rect 2158 15292 2210 15344
rect 2222 15292 2274 15344
rect 2286 15292 2338 15344
rect 7966 15292 8018 15344
rect 8030 15292 8082 15344
rect 8094 15292 8146 15344
rect 8158 15292 8210 15344
rect 8222 15292 8274 15344
rect 8286 15292 8338 15344
rect 6742 15076 6794 15085
rect 6742 15042 6751 15076
rect 6751 15042 6785 15076
rect 6785 15042 6794 15076
rect 6742 15033 6794 15042
rect 7606 15033 7658 15085
rect 7894 14959 7946 15011
rect 9814 14737 9866 14789
rect 4966 14626 5018 14678
rect 5030 14626 5082 14678
rect 5094 14626 5146 14678
rect 5158 14626 5210 14678
rect 5222 14626 5274 14678
rect 5286 14626 5338 14678
rect 7414 14410 7466 14419
rect 7414 14376 7423 14410
rect 7423 14376 7457 14410
rect 7457 14376 7466 14410
rect 7414 14367 7466 14376
rect 7894 14293 7946 14345
rect 886 14219 938 14271
rect 3766 14219 3818 14271
rect 5782 14219 5834 14271
rect 7606 14219 7658 14271
rect 9430 14114 9482 14123
rect 9430 14080 9439 14114
rect 9439 14080 9473 14114
rect 9473 14080 9482 14114
rect 9430 14071 9482 14080
rect 1966 13960 2018 14012
rect 2030 13960 2082 14012
rect 2094 13960 2146 14012
rect 2158 13960 2210 14012
rect 2222 13960 2274 14012
rect 2286 13960 2338 14012
rect 7966 13960 8018 14012
rect 8030 13960 8082 14012
rect 8094 13960 8146 14012
rect 8158 13960 8210 14012
rect 8222 13960 8274 14012
rect 8286 13960 8338 14012
rect 9814 13670 9866 13679
rect 9814 13636 9823 13670
rect 9823 13636 9857 13670
rect 9857 13636 9866 13670
rect 9814 13627 9866 13636
rect 10102 13448 10154 13457
rect 10102 13414 10111 13448
rect 10111 13414 10145 13448
rect 10145 13414 10154 13448
rect 10102 13405 10154 13414
rect 4966 13294 5018 13346
rect 5030 13294 5082 13346
rect 5094 13294 5146 13346
rect 5158 13294 5210 13346
rect 5222 13294 5274 13346
rect 5286 13294 5338 13346
rect 4630 13183 4682 13235
rect 2614 13035 2666 13087
rect 4150 12961 4202 13013
rect 2806 12887 2858 12939
rect 1966 12628 2018 12680
rect 2030 12628 2082 12680
rect 2094 12628 2146 12680
rect 2158 12628 2210 12680
rect 2222 12628 2274 12680
rect 2286 12628 2338 12680
rect 7966 12628 8018 12680
rect 8030 12628 8082 12680
rect 8094 12628 8146 12680
rect 8158 12628 8210 12680
rect 8222 12628 8274 12680
rect 8286 12628 8338 12680
rect 5686 12517 5738 12569
rect 2806 12369 2858 12421
rect 4630 12369 4682 12421
rect 7510 12369 7562 12421
rect 2998 12295 3050 12347
rect 4150 12295 4202 12347
rect 3670 12221 3722 12273
rect 3190 12073 3242 12125
rect 4966 11962 5018 12014
rect 5030 11962 5082 12014
rect 5094 11962 5146 12014
rect 5158 11962 5210 12014
rect 5222 11962 5274 12014
rect 5286 11962 5338 12014
rect 2614 11894 2666 11903
rect 2614 11860 2623 11894
rect 2623 11860 2657 11894
rect 2657 11860 2666 11894
rect 2614 11851 2666 11860
rect 8470 11894 8522 11903
rect 8470 11860 8479 11894
rect 8479 11860 8513 11894
rect 8513 11860 8522 11894
rect 8470 11851 8522 11860
rect 2998 11703 3050 11755
rect 5686 11703 5738 11755
rect 4150 11629 4202 11681
rect 7126 11629 7178 11681
rect 2806 11481 2858 11533
rect 7510 11555 7562 11607
rect 6070 11481 6122 11533
rect 1966 11296 2018 11348
rect 2030 11296 2082 11348
rect 2094 11296 2146 11348
rect 2158 11296 2210 11348
rect 2222 11296 2274 11348
rect 2286 11296 2338 11348
rect 7966 11296 8018 11348
rect 8030 11296 8082 11348
rect 8094 11296 8146 11348
rect 8158 11296 8210 11348
rect 8222 11296 8274 11348
rect 8286 11296 8338 11348
rect 6070 11185 6122 11237
rect 7510 11185 7562 11237
rect 8374 11185 8426 11237
rect 2806 11037 2858 11089
rect 3670 11037 3722 11089
rect 6838 11111 6890 11163
rect 8182 11111 8234 11163
rect 7510 11037 7562 11089
rect 2614 10963 2666 11015
rect 5686 10963 5738 11015
rect 7126 11006 7178 11015
rect 7126 10972 7135 11006
rect 7135 10972 7169 11006
rect 7169 10972 7178 11006
rect 7126 10963 7178 10972
rect 9622 10963 9674 11015
rect 3670 10889 3722 10941
rect 4534 10741 4586 10793
rect 6550 10784 6602 10793
rect 6550 10750 6559 10784
rect 6559 10750 6593 10784
rect 6593 10750 6602 10784
rect 6550 10741 6602 10750
rect 10102 10784 10154 10793
rect 10102 10750 10111 10784
rect 10111 10750 10145 10784
rect 10145 10750 10154 10784
rect 10102 10741 10154 10750
rect 4966 10630 5018 10682
rect 5030 10630 5082 10682
rect 5094 10630 5146 10682
rect 5158 10630 5210 10682
rect 5222 10630 5274 10682
rect 5286 10630 5338 10682
rect 4150 10519 4202 10571
rect 7798 10519 7850 10571
rect 8182 10519 8234 10571
rect 886 10371 938 10423
rect 3670 10371 3722 10423
rect 5878 10371 5930 10423
rect 6646 10414 6698 10423
rect 6646 10380 6655 10414
rect 6655 10380 6689 10414
rect 6689 10380 6698 10414
rect 6646 10371 6698 10380
rect 4630 10297 4682 10349
rect 7126 10297 7178 10349
rect 7510 10149 7562 10201
rect 5590 10075 5642 10127
rect 1966 9964 2018 10016
rect 2030 9964 2082 10016
rect 2094 9964 2146 10016
rect 2158 9964 2210 10016
rect 2222 9964 2274 10016
rect 2286 9964 2338 10016
rect 7966 9964 8018 10016
rect 8030 9964 8082 10016
rect 8094 9964 8146 10016
rect 8158 9964 8210 10016
rect 8222 9964 8274 10016
rect 8286 9964 8338 10016
rect 6646 9853 6698 9905
rect 7126 9853 7178 9905
rect 7510 9705 7562 9757
rect 7030 9631 7082 9683
rect 6358 9557 6410 9609
rect 8470 9557 8522 9609
rect 4966 9298 5018 9350
rect 5030 9298 5082 9350
rect 5094 9298 5146 9350
rect 5158 9298 5210 9350
rect 5222 9298 5274 9350
rect 5286 9298 5338 9350
rect 8374 8965 8426 9017
rect 5878 8891 5930 8943
rect 6742 8891 6794 8943
rect 7510 8817 7562 8869
rect 9526 8743 9578 8795
rect 1966 8632 2018 8684
rect 2030 8632 2082 8684
rect 2094 8632 2146 8684
rect 2158 8632 2210 8684
rect 2222 8632 2274 8684
rect 2286 8632 2338 8684
rect 7966 8632 8018 8684
rect 8030 8632 8082 8684
rect 8094 8632 8146 8684
rect 8158 8632 8210 8684
rect 8222 8632 8274 8684
rect 8286 8632 8338 8684
rect 1846 8299 1898 8351
rect 6742 8416 6794 8425
rect 6742 8382 6751 8416
rect 6751 8382 6785 8416
rect 6785 8382 6794 8416
rect 6742 8373 6794 8382
rect 7510 8373 7562 8425
rect 4246 8299 4298 8351
rect 7126 8342 7178 8351
rect 7126 8308 7135 8342
rect 7135 8308 7169 8342
rect 7169 8308 7178 8342
rect 7126 8299 7178 8308
rect 9430 8299 9482 8351
rect 10102 8342 10154 8351
rect 10102 8308 10111 8342
rect 10111 8308 10145 8342
rect 10145 8308 10154 8342
rect 10102 8299 10154 8308
rect 9238 8077 9290 8129
rect 4966 7966 5018 8018
rect 5030 7966 5082 8018
rect 5094 7966 5146 8018
rect 5158 7966 5210 8018
rect 5222 7966 5274 8018
rect 5286 7966 5338 8018
rect 2902 7855 2954 7907
rect 1462 7781 1514 7833
rect 2710 7633 2762 7685
rect 1942 7559 1994 7611
rect 3478 7559 3530 7611
rect 2422 7454 2474 7463
rect 2422 7420 2431 7454
rect 2431 7420 2465 7454
rect 2465 7420 2474 7454
rect 2422 7411 2474 7420
rect 2998 7454 3050 7463
rect 2998 7420 3007 7454
rect 3007 7420 3041 7454
rect 3041 7420 3050 7454
rect 2998 7411 3050 7420
rect 5782 7707 5834 7759
rect 6742 7707 6794 7759
rect 3862 7633 3914 7685
rect 7798 7676 7850 7685
rect 7798 7642 7807 7676
rect 7807 7642 7841 7676
rect 7841 7642 7850 7676
rect 7798 7633 7850 7642
rect 7510 7559 7562 7611
rect 4630 7411 4682 7463
rect 9622 7411 9674 7463
rect 1966 7300 2018 7352
rect 2030 7300 2082 7352
rect 2094 7300 2146 7352
rect 2158 7300 2210 7352
rect 2222 7300 2274 7352
rect 2286 7300 2338 7352
rect 7966 7300 8018 7352
rect 8030 7300 8082 7352
rect 8094 7300 8146 7352
rect 8158 7300 8210 7352
rect 8222 7300 8274 7352
rect 8286 7300 8338 7352
rect 3478 7232 3530 7241
rect 3478 7198 3487 7232
rect 3487 7198 3521 7232
rect 3521 7198 3530 7232
rect 3478 7189 3530 7198
rect 4630 7189 4682 7241
rect 7510 7189 7562 7241
rect 2998 7115 3050 7167
rect 4150 7115 4202 7167
rect 2422 7041 2474 7093
rect 1846 6967 1898 7019
rect 2230 6967 2282 7019
rect 1558 6893 1610 6945
rect 2710 7041 2762 7093
rect 4150 7010 4202 7019
rect 4150 6976 4159 7010
rect 4159 6976 4193 7010
rect 4193 6976 4202 7010
rect 4150 6967 4202 6976
rect 4726 7010 4778 7019
rect 4726 6976 4735 7010
rect 4735 6976 4769 7010
rect 4769 6976 4778 7010
rect 4726 6967 4778 6976
rect 4438 6893 4490 6945
rect 4822 6893 4874 6945
rect 2806 6819 2858 6871
rect 6358 7010 6410 7019
rect 6358 6976 6367 7010
rect 6367 6976 6401 7010
rect 6401 6976 6410 7010
rect 6358 6967 6410 6976
rect 5686 6893 5738 6945
rect 6742 6893 6794 6945
rect 3286 6745 3338 6797
rect 3862 6788 3914 6797
rect 3862 6754 3871 6788
rect 3871 6754 3905 6788
rect 3905 6754 3914 6788
rect 3862 6745 3914 6754
rect 3958 6745 4010 6797
rect 5398 6745 5450 6797
rect 7894 6745 7946 6797
rect 4966 6634 5018 6686
rect 5030 6634 5082 6686
rect 5094 6634 5146 6686
rect 5158 6634 5210 6686
rect 5222 6634 5274 6686
rect 5286 6634 5338 6686
rect 1462 6523 1514 6575
rect 2902 6523 2954 6575
rect 4630 6566 4682 6575
rect 4630 6532 4639 6566
rect 4639 6532 4673 6566
rect 4673 6532 4682 6566
rect 4630 6523 4682 6532
rect 1558 6418 1610 6427
rect 1558 6384 1567 6418
rect 1567 6384 1601 6418
rect 1601 6384 1610 6418
rect 1558 6375 1610 6384
rect 1750 6344 1802 6353
rect 1750 6310 1759 6344
rect 1759 6310 1793 6344
rect 1793 6310 1802 6344
rect 1750 6301 1802 6310
rect 2422 6449 2474 6501
rect 2806 6492 2858 6501
rect 2806 6458 2815 6492
rect 2815 6458 2849 6492
rect 2849 6458 2858 6492
rect 2806 6449 2858 6458
rect 5686 6492 5738 6501
rect 5686 6458 5695 6492
rect 5695 6458 5729 6492
rect 5729 6458 5738 6492
rect 5686 6449 5738 6458
rect 3286 6418 3338 6427
rect 3286 6384 3295 6418
rect 3295 6384 3329 6418
rect 3329 6384 3338 6418
rect 3286 6375 3338 6384
rect 4822 6418 4874 6427
rect 4822 6384 4831 6418
rect 4831 6384 4865 6418
rect 4865 6384 4874 6418
rect 4822 6375 4874 6384
rect 2230 6301 2282 6353
rect 3862 6301 3914 6353
rect 5782 6418 5834 6427
rect 5782 6384 5791 6418
rect 5791 6384 5825 6418
rect 5825 6384 5834 6418
rect 5782 6375 5834 6384
rect 5110 6344 5162 6353
rect 5110 6310 5119 6344
rect 5119 6310 5153 6344
rect 5153 6310 5162 6344
rect 5110 6301 5162 6310
rect 9718 6301 9770 6353
rect 3862 6153 3914 6205
rect 4246 6079 4298 6131
rect 4438 6079 4490 6131
rect 5494 6079 5546 6131
rect 10102 6122 10154 6131
rect 10102 6088 10111 6122
rect 10111 6088 10145 6122
rect 10145 6088 10154 6122
rect 10102 6079 10154 6088
rect 1966 5968 2018 6020
rect 2030 5968 2082 6020
rect 2094 5968 2146 6020
rect 2158 5968 2210 6020
rect 2222 5968 2274 6020
rect 2286 5968 2338 6020
rect 7966 5968 8018 6020
rect 8030 5968 8082 6020
rect 8094 5968 8146 6020
rect 8158 5968 8210 6020
rect 8222 5968 8274 6020
rect 8286 5968 8338 6020
rect 5110 5857 5162 5909
rect 3958 5783 4010 5835
rect 4534 5709 4586 5761
rect 5878 5709 5930 5761
rect 1750 5678 1802 5687
rect 1750 5644 1759 5678
rect 1759 5644 1793 5678
rect 1793 5644 1802 5678
rect 1750 5635 1802 5644
rect 1846 5635 1898 5687
rect 3862 5678 3914 5687
rect 3862 5644 3871 5678
rect 3871 5644 3905 5678
rect 3905 5644 3914 5678
rect 3862 5635 3914 5644
rect 5686 5635 5738 5687
rect 5878 5561 5930 5613
rect 2422 5487 2474 5539
rect 3574 5413 3626 5465
rect 4822 5413 4874 5465
rect 5494 5413 5546 5465
rect 4966 5302 5018 5354
rect 5030 5302 5082 5354
rect 5094 5302 5146 5354
rect 5158 5302 5210 5354
rect 5222 5302 5274 5354
rect 5286 5302 5338 5354
rect 4726 5191 4778 5243
rect 5686 5191 5738 5243
rect 5782 5191 5834 5243
rect 4150 5117 4202 5169
rect 4246 5086 4298 5095
rect 4246 5052 4255 5086
rect 4255 5052 4289 5086
rect 4289 5052 4298 5086
rect 4246 5043 4298 5052
rect 5494 5086 5546 5095
rect 5494 5052 5503 5086
rect 5503 5052 5537 5086
rect 5537 5052 5546 5086
rect 5494 5043 5546 5052
rect 3862 5012 3914 5021
rect 3862 4978 3871 5012
rect 3871 4978 3905 5012
rect 3905 4978 3914 5012
rect 3862 4969 3914 4978
rect 5878 5117 5930 5169
rect 5398 4895 5450 4947
rect 1750 4821 1802 4873
rect 1966 4636 2018 4688
rect 2030 4636 2082 4688
rect 2094 4636 2146 4688
rect 2158 4636 2210 4688
rect 2222 4636 2274 4688
rect 2286 4636 2338 4688
rect 7966 4636 8018 4688
rect 8030 4636 8082 4688
rect 8094 4636 8146 4688
rect 8158 4636 8210 4688
rect 8222 4636 8274 4688
rect 8286 4636 8338 4688
rect 3862 4377 3914 4429
rect 1654 4303 1706 4355
rect 4534 4346 4586 4355
rect 4534 4312 4543 4346
rect 4543 4312 4577 4346
rect 4577 4312 4586 4346
rect 4534 4303 4586 4312
rect 598 4081 650 4133
rect 4966 3970 5018 4022
rect 5030 3970 5082 4022
rect 5094 3970 5146 4022
rect 5158 3970 5210 4022
rect 5222 3970 5274 4022
rect 5286 3970 5338 4022
rect 5494 3859 5546 3911
rect 3574 3711 3626 3763
rect 2518 3637 2570 3689
rect 3862 3680 3914 3689
rect 3862 3646 3871 3680
rect 3871 3646 3905 3680
rect 3905 3646 3914 3680
rect 3862 3637 3914 3646
rect 9526 3680 9578 3689
rect 9526 3646 9535 3680
rect 9535 3646 9569 3680
rect 9569 3646 9578 3680
rect 9526 3637 9578 3646
rect 9910 3680 9962 3689
rect 9910 3646 9919 3680
rect 9919 3646 9953 3680
rect 9953 3646 9962 3680
rect 9910 3637 9962 3646
rect 10102 3606 10154 3615
rect 10102 3572 10111 3606
rect 10111 3572 10145 3606
rect 10145 3572 10154 3606
rect 10102 3563 10154 3572
rect 1846 3458 1898 3467
rect 1846 3424 1855 3458
rect 1855 3424 1889 3458
rect 1889 3424 1898 3458
rect 1846 3415 1898 3424
rect 10966 3415 11018 3467
rect 1966 3304 2018 3356
rect 2030 3304 2082 3356
rect 2094 3304 2146 3356
rect 2158 3304 2210 3356
rect 2222 3304 2274 3356
rect 2286 3304 2338 3356
rect 7966 3304 8018 3356
rect 8030 3304 8082 3356
rect 8094 3304 8146 3356
rect 8158 3304 8210 3356
rect 8222 3304 8274 3356
rect 8286 3304 8338 3356
rect 1462 3193 1514 3245
rect 1558 3014 1610 3023
rect 1558 2980 1567 3014
rect 1567 2980 1601 3014
rect 1601 2980 1610 3014
rect 1558 2971 1610 2980
rect 3190 3014 3242 3023
rect 3190 2980 3199 3014
rect 3199 2980 3233 3014
rect 3233 2980 3242 3014
rect 3190 2971 3242 2980
rect 4630 2971 4682 3023
rect 5590 3014 5642 3023
rect 5590 2980 5599 3014
rect 5599 2980 5633 3014
rect 5633 2980 5642 3014
rect 5590 2971 5642 2980
rect 6550 2971 6602 3023
rect 7894 3014 7946 3023
rect 7894 2980 7903 3014
rect 7903 2980 7937 3014
rect 7937 2980 7946 3014
rect 7894 2971 7946 2980
rect 9238 3014 9290 3023
rect 9238 2980 9247 3014
rect 9247 2980 9281 3014
rect 9281 2980 9290 3014
rect 9238 2971 9290 2980
rect 9334 2971 9386 3023
rect 9622 2971 9674 3023
rect 2902 2897 2954 2949
rect 4054 2897 4106 2949
rect 5398 2897 5450 2949
rect 6358 2897 6410 2949
rect 7606 2940 7658 2949
rect 7606 2906 7615 2940
rect 7615 2906 7649 2940
rect 7649 2906 7658 2940
rect 7606 2897 7658 2906
rect 8662 2897 8714 2949
rect 9718 2940 9770 2949
rect 9718 2906 9727 2940
rect 9727 2906 9761 2940
rect 9761 2906 9770 2940
rect 9718 2897 9770 2906
rect 9814 2940 9866 2949
rect 9814 2906 9823 2940
rect 9823 2906 9857 2940
rect 9857 2906 9866 2940
rect 9814 2897 9866 2906
rect 4966 2638 5018 2690
rect 5030 2638 5082 2690
rect 5094 2638 5146 2690
rect 5158 2638 5210 2690
rect 5222 2638 5274 2690
rect 5286 2638 5338 2690
<< metal2 >>
rect 308 28074 364 28874
rect 884 28074 940 28874
rect 1460 28208 1516 28874
rect 2036 28208 2092 28874
rect 1460 28180 1598 28208
rect 1460 28074 1516 28180
rect 322 25155 350 28074
rect 310 25149 362 25155
rect 310 25091 362 25097
rect 898 24489 926 28074
rect 1460 26742 1516 26751
rect 1460 26677 1516 26686
rect 1474 25229 1502 26677
rect 1570 25895 1598 28180
rect 1858 28180 2092 28208
rect 1858 25895 1886 28180
rect 2036 28074 2092 28180
rect 2612 28074 2668 28874
rect 3188 28208 3244 28874
rect 3764 28208 3820 28874
rect 4340 28208 4396 28874
rect 4916 28208 4972 28874
rect 3188 28180 3326 28208
rect 3188 28074 3244 28180
rect 1964 26002 2340 26011
rect 2020 26000 2044 26002
rect 2100 26000 2124 26002
rect 2180 26000 2204 26002
rect 2260 26000 2284 26002
rect 2020 25948 2030 26000
rect 2274 25948 2284 26000
rect 2020 25946 2044 25948
rect 2100 25946 2124 25948
rect 2180 25946 2204 25948
rect 2260 25946 2284 25948
rect 1964 25937 2340 25946
rect 2626 25895 2654 28074
rect 3298 25895 3326 28180
rect 3764 28180 3902 28208
rect 3764 28074 3820 28180
rect 3874 25895 3902 28180
rect 4340 28180 4478 28208
rect 4340 28074 4396 28180
rect 4450 25895 4478 28180
rect 4916 28180 5054 28208
rect 4916 28074 4972 28180
rect 5026 25895 5054 28180
rect 5492 28074 5548 28874
rect 6068 28208 6124 28874
rect 6644 28208 6700 28874
rect 7220 28208 7276 28874
rect 7796 28208 7852 28874
rect 8372 28208 8428 28874
rect 8948 28208 9004 28874
rect 9524 28208 9580 28874
rect 6068 28180 6302 28208
rect 6068 28074 6124 28180
rect 5506 25895 5534 28074
rect 6274 25895 6302 28180
rect 6644 28180 6782 28208
rect 6644 28074 6700 28180
rect 6754 25895 6782 28180
rect 7220 28180 7358 28208
rect 7220 28074 7276 28180
rect 7330 25895 7358 28180
rect 7796 28180 7934 28208
rect 7796 28074 7852 28180
rect 7906 25895 7934 28180
rect 8372 28180 8510 28208
rect 8372 28074 8428 28180
rect 7964 26002 8340 26011
rect 8020 26000 8044 26002
rect 8100 26000 8124 26002
rect 8180 26000 8204 26002
rect 8260 26000 8284 26002
rect 8020 25948 8030 26000
rect 8274 25948 8284 26000
rect 8020 25946 8044 25948
rect 8100 25946 8124 25948
rect 8180 25946 8204 25948
rect 8260 25946 8284 25948
rect 7964 25937 8340 25946
rect 8482 25895 8510 28180
rect 8948 28180 9086 28208
rect 8948 28074 9004 28180
rect 9058 25895 9086 28180
rect 9524 28180 9662 28208
rect 9524 28074 9580 28180
rect 9332 27334 9388 27343
rect 9332 27269 9388 27278
rect 1558 25889 1610 25895
rect 1558 25831 1610 25837
rect 1846 25889 1898 25895
rect 1846 25831 1898 25837
rect 2614 25889 2666 25895
rect 2614 25831 2666 25837
rect 3286 25889 3338 25895
rect 3286 25831 3338 25837
rect 3862 25889 3914 25895
rect 3862 25831 3914 25837
rect 4438 25889 4490 25895
rect 4438 25831 4490 25837
rect 5014 25889 5066 25895
rect 5014 25831 5066 25837
rect 5494 25889 5546 25895
rect 5494 25831 5546 25837
rect 6262 25889 6314 25895
rect 6262 25831 6314 25837
rect 6742 25889 6794 25895
rect 6742 25831 6794 25837
rect 7318 25889 7370 25895
rect 7318 25831 7370 25837
rect 7894 25889 7946 25895
rect 7894 25831 7946 25837
rect 8470 25889 8522 25895
rect 8470 25831 8522 25837
rect 9046 25889 9098 25895
rect 9046 25831 9098 25837
rect 5974 25815 6026 25821
rect 5974 25757 6026 25763
rect 3670 25741 3722 25747
rect 3670 25683 3722 25689
rect 1654 25667 1706 25673
rect 1654 25609 1706 25615
rect 2902 25667 2954 25673
rect 2902 25609 2954 25615
rect 2998 25667 3050 25673
rect 2998 25609 3050 25615
rect 1462 25223 1514 25229
rect 1462 25165 1514 25171
rect 886 24483 938 24489
rect 886 24425 938 24431
rect 1666 22787 1694 25609
rect 2614 25075 2666 25081
rect 2614 25017 2666 25023
rect 1846 25001 1898 25007
rect 1846 24943 1898 24949
rect 1750 24335 1802 24341
rect 1750 24277 1802 24283
rect 1654 22781 1706 22787
rect 1654 22723 1706 22729
rect 1268 22598 1324 22607
rect 1268 22533 1270 22542
rect 1322 22533 1324 22542
rect 1270 22501 1322 22507
rect 1762 21751 1790 24277
rect 1750 21745 1802 21751
rect 1750 21687 1802 21693
rect 1762 19753 1790 21687
rect 1750 19747 1802 19753
rect 1750 19689 1802 19695
rect 1654 18933 1706 18939
rect 1654 18875 1706 18881
rect 1666 18463 1694 18875
rect 1652 18454 1708 18463
rect 1652 18389 1708 18398
rect 1654 15455 1706 15461
rect 1654 15397 1706 15403
rect 884 14310 940 14319
rect 884 14245 886 14254
rect 938 14245 940 14254
rect 886 14213 938 14219
rect 886 10423 938 10429
rect 886 10365 938 10371
rect 898 10175 926 10365
rect 884 10166 940 10175
rect 884 10101 940 10110
rect 1462 7833 1514 7839
rect 1462 7775 1514 7781
rect 1474 6581 1502 7775
rect 1558 6945 1610 6951
rect 1558 6887 1610 6893
rect 1462 6575 1514 6581
rect 1462 6517 1514 6523
rect 598 4133 650 4139
rect 598 4075 650 4081
rect 610 800 638 4075
rect 1474 3251 1502 6517
rect 1570 6433 1598 6887
rect 1558 6427 1610 6433
rect 1558 6369 1610 6375
rect 1666 4361 1694 15397
rect 1858 8524 1886 24943
rect 1964 24670 2340 24679
rect 2020 24668 2044 24670
rect 2100 24668 2124 24670
rect 2180 24668 2204 24670
rect 2260 24668 2284 24670
rect 2020 24616 2030 24668
rect 2274 24616 2284 24668
rect 2020 24614 2044 24616
rect 2100 24614 2124 24616
rect 2180 24614 2204 24616
rect 2260 24614 2284 24616
rect 1964 24605 2340 24614
rect 1964 23338 2340 23347
rect 2020 23336 2044 23338
rect 2100 23336 2124 23338
rect 2180 23336 2204 23338
rect 2260 23336 2284 23338
rect 2020 23284 2030 23336
rect 2274 23284 2284 23336
rect 2020 23282 2044 23284
rect 2100 23282 2124 23284
rect 2180 23282 2204 23284
rect 2260 23282 2284 23284
rect 1964 23273 2340 23282
rect 1964 22006 2340 22015
rect 2020 22004 2044 22006
rect 2100 22004 2124 22006
rect 2180 22004 2204 22006
rect 2260 22004 2284 22006
rect 2020 21952 2030 22004
rect 2274 21952 2284 22004
rect 2020 21950 2044 21952
rect 2100 21950 2124 21952
rect 2180 21950 2204 21952
rect 2260 21950 2284 21952
rect 1964 21941 2340 21950
rect 2626 21011 2654 25017
rect 2710 22781 2762 22787
rect 2710 22723 2762 22729
rect 2722 21011 2750 22723
rect 2914 21233 2942 25609
rect 2902 21227 2954 21233
rect 2902 21169 2954 21175
rect 2614 21005 2666 21011
rect 2614 20947 2666 20953
rect 2710 21005 2762 21011
rect 2710 20947 2762 20953
rect 1964 20674 2340 20683
rect 2020 20672 2044 20674
rect 2100 20672 2124 20674
rect 2180 20672 2204 20674
rect 2260 20672 2284 20674
rect 2020 20620 2030 20672
rect 2274 20620 2284 20672
rect 2020 20618 2044 20620
rect 2100 20618 2124 20620
rect 2180 20618 2204 20620
rect 2260 20618 2284 20620
rect 1964 20609 2340 20618
rect 1964 19342 2340 19351
rect 2020 19340 2044 19342
rect 2100 19340 2124 19342
rect 2180 19340 2204 19342
rect 2260 19340 2284 19342
rect 2020 19288 2030 19340
rect 2274 19288 2284 19340
rect 2020 19286 2044 19288
rect 2100 19286 2124 19288
rect 2180 19286 2204 19288
rect 2260 19286 2284 19288
rect 1964 19277 2340 19286
rect 1964 18010 2340 18019
rect 2020 18008 2044 18010
rect 2100 18008 2124 18010
rect 2180 18008 2204 18010
rect 2260 18008 2284 18010
rect 2020 17956 2030 18008
rect 2274 17956 2284 18008
rect 2020 17954 2044 17956
rect 2100 17954 2124 17956
rect 2180 17954 2204 17956
rect 2260 17954 2284 17956
rect 1964 17945 2340 17954
rect 1964 16678 2340 16687
rect 2020 16676 2044 16678
rect 2100 16676 2124 16678
rect 2180 16676 2204 16678
rect 2260 16676 2284 16678
rect 2020 16624 2030 16676
rect 2274 16624 2284 16676
rect 2020 16622 2044 16624
rect 2100 16622 2124 16624
rect 2180 16622 2204 16624
rect 2260 16622 2284 16624
rect 1964 16613 2340 16622
rect 2518 16121 2570 16127
rect 2518 16063 2570 16069
rect 1964 15346 2340 15355
rect 2020 15344 2044 15346
rect 2100 15344 2124 15346
rect 2180 15344 2204 15346
rect 2260 15344 2284 15346
rect 2020 15292 2030 15344
rect 2274 15292 2284 15344
rect 2020 15290 2044 15292
rect 2100 15290 2124 15292
rect 2180 15290 2204 15292
rect 2260 15290 2284 15292
rect 1964 15281 2340 15290
rect 1964 14014 2340 14023
rect 2020 14012 2044 14014
rect 2100 14012 2124 14014
rect 2180 14012 2204 14014
rect 2260 14012 2284 14014
rect 2020 13960 2030 14012
rect 2274 13960 2284 14012
rect 2020 13958 2044 13960
rect 2100 13958 2124 13960
rect 2180 13958 2204 13960
rect 2260 13958 2284 13960
rect 1964 13949 2340 13958
rect 1964 12682 2340 12691
rect 2020 12680 2044 12682
rect 2100 12680 2124 12682
rect 2180 12680 2204 12682
rect 2260 12680 2284 12682
rect 2020 12628 2030 12680
rect 2274 12628 2284 12680
rect 2020 12626 2044 12628
rect 2100 12626 2124 12628
rect 2180 12626 2204 12628
rect 2260 12626 2284 12628
rect 1964 12617 2340 12626
rect 1964 11350 2340 11359
rect 2020 11348 2044 11350
rect 2100 11348 2124 11350
rect 2180 11348 2204 11350
rect 2260 11348 2284 11350
rect 2020 11296 2030 11348
rect 2274 11296 2284 11348
rect 2020 11294 2044 11296
rect 2100 11294 2124 11296
rect 2180 11294 2204 11296
rect 2260 11294 2284 11296
rect 1964 11285 2340 11294
rect 1964 10018 2340 10027
rect 2020 10016 2044 10018
rect 2100 10016 2124 10018
rect 2180 10016 2204 10018
rect 2260 10016 2284 10018
rect 2020 9964 2030 10016
rect 2274 9964 2284 10016
rect 2020 9962 2044 9964
rect 2100 9962 2124 9964
rect 2180 9962 2204 9964
rect 2260 9962 2284 9964
rect 1964 9953 2340 9962
rect 1964 8686 2340 8695
rect 2020 8684 2044 8686
rect 2100 8684 2124 8686
rect 2180 8684 2204 8686
rect 2260 8684 2284 8686
rect 2020 8632 2030 8684
rect 2274 8632 2284 8684
rect 2020 8630 2044 8632
rect 2100 8630 2124 8632
rect 2180 8630 2204 8632
rect 2260 8630 2284 8632
rect 1964 8621 2340 8630
rect 1858 8496 1982 8524
rect 1846 8351 1898 8357
rect 1846 8293 1898 8299
rect 1858 7025 1886 8293
rect 1954 7617 1982 8496
rect 1942 7611 1994 7617
rect 1942 7553 1994 7559
rect 2422 7463 2474 7469
rect 2422 7405 2474 7411
rect 1964 7354 2340 7363
rect 2020 7352 2044 7354
rect 2100 7352 2124 7354
rect 2180 7352 2204 7354
rect 2260 7352 2284 7354
rect 2020 7300 2030 7352
rect 2274 7300 2284 7352
rect 2020 7298 2044 7300
rect 2100 7298 2124 7300
rect 2180 7298 2204 7300
rect 2260 7298 2284 7300
rect 1964 7289 2340 7298
rect 2434 7099 2462 7405
rect 2422 7093 2474 7099
rect 2422 7035 2474 7041
rect 1846 7019 1898 7025
rect 1846 6961 1898 6967
rect 2230 7019 2282 7025
rect 2230 6961 2282 6967
rect 1750 6353 1802 6359
rect 1748 6318 1750 6327
rect 1802 6318 1804 6327
rect 1748 6253 1804 6262
rect 1858 5693 1886 6961
rect 2242 6359 2270 6961
rect 2422 6501 2474 6507
rect 2422 6443 2474 6449
rect 2230 6353 2282 6359
rect 2230 6295 2282 6301
rect 1964 6022 2340 6031
rect 2020 6020 2044 6022
rect 2100 6020 2124 6022
rect 2180 6020 2204 6022
rect 2260 6020 2284 6022
rect 2020 5968 2030 6020
rect 2274 5968 2284 6020
rect 2020 5966 2044 5968
rect 2100 5966 2124 5968
rect 2180 5966 2204 5968
rect 2260 5966 2284 5968
rect 1964 5957 2340 5966
rect 1750 5687 1802 5693
rect 1750 5629 1802 5635
rect 1846 5687 1898 5693
rect 1846 5629 1898 5635
rect 1762 4879 1790 5629
rect 2434 5545 2462 6443
rect 2422 5539 2474 5545
rect 2422 5481 2474 5487
rect 1750 4873 1802 4879
rect 1750 4815 1802 4821
rect 1964 4690 2340 4699
rect 2020 4688 2044 4690
rect 2100 4688 2124 4690
rect 2180 4688 2204 4690
rect 2260 4688 2284 4690
rect 2020 4636 2030 4688
rect 2274 4636 2284 4688
rect 2020 4634 2044 4636
rect 2100 4634 2124 4636
rect 2180 4634 2204 4636
rect 2260 4634 2284 4636
rect 1964 4625 2340 4634
rect 1654 4355 1706 4361
rect 1654 4297 1706 4303
rect 2530 3695 2558 16063
rect 2626 13093 2654 20947
rect 2902 18563 2954 18569
rect 2902 18505 2954 18511
rect 2806 16417 2858 16423
rect 2806 16359 2858 16365
rect 2818 15609 2846 16359
rect 2806 15603 2858 15609
rect 2806 15545 2858 15551
rect 2614 13087 2666 13093
rect 2614 13029 2666 13035
rect 2626 11909 2654 13029
rect 2818 12945 2846 15545
rect 2914 13112 2942 18505
rect 3010 17237 3038 25609
rect 3286 25223 3338 25229
rect 3286 25165 3338 25171
rect 3298 21677 3326 25165
rect 3382 25149 3434 25155
rect 3382 25091 3434 25097
rect 3394 23009 3422 25091
rect 3478 23077 3530 23083
rect 3478 23019 3530 23025
rect 3382 23003 3434 23009
rect 3382 22945 3434 22951
rect 3286 21671 3338 21677
rect 3286 21613 3338 21619
rect 3298 18421 3326 21613
rect 3394 18569 3422 22945
rect 3490 22269 3518 23019
rect 3682 22343 3710 25683
rect 5782 25667 5834 25673
rect 5782 25609 5834 25615
rect 5878 25667 5930 25673
rect 5878 25609 5930 25615
rect 5398 25445 5450 25451
rect 5398 25387 5450 25393
rect 4964 25336 5340 25345
rect 5020 25334 5044 25336
rect 5100 25334 5124 25336
rect 5180 25334 5204 25336
rect 5260 25334 5284 25336
rect 5020 25282 5030 25334
rect 5274 25282 5284 25334
rect 5020 25280 5044 25282
rect 5100 25280 5124 25282
rect 5180 25280 5204 25282
rect 5260 25280 5284 25282
rect 4964 25271 5340 25280
rect 4246 25001 4298 25007
rect 4246 24943 4298 24949
rect 4150 24261 4202 24267
rect 4150 24203 4202 24209
rect 4162 23601 4190 24203
rect 4150 23595 4202 23601
rect 4150 23537 4202 23543
rect 4162 22935 4190 23537
rect 3766 22929 3818 22935
rect 3766 22871 3818 22877
rect 4150 22929 4202 22935
rect 4150 22871 4202 22877
rect 3778 22417 3806 22871
rect 4258 22565 4286 24943
rect 4964 24004 5340 24013
rect 5020 24002 5044 24004
rect 5100 24002 5124 24004
rect 5180 24002 5204 24004
rect 5260 24002 5284 24004
rect 5020 23950 5030 24002
rect 5274 23950 5284 24002
rect 5020 23948 5044 23950
rect 5100 23948 5124 23950
rect 5180 23948 5204 23950
rect 5260 23948 5284 23950
rect 4964 23939 5340 23948
rect 4964 22672 5340 22681
rect 5020 22670 5044 22672
rect 5100 22670 5124 22672
rect 5180 22670 5204 22672
rect 5260 22670 5284 22672
rect 5020 22618 5030 22670
rect 5274 22618 5284 22670
rect 5020 22616 5044 22618
rect 5100 22616 5124 22618
rect 5180 22616 5204 22618
rect 5260 22616 5284 22618
rect 4964 22607 5340 22616
rect 4246 22559 4298 22565
rect 4246 22501 4298 22507
rect 3766 22411 3818 22417
rect 3766 22353 3818 22359
rect 3670 22337 3722 22343
rect 3586 22297 3670 22325
rect 3478 22263 3530 22269
rect 3478 22205 3530 22211
rect 3490 21751 3518 22205
rect 3478 21745 3530 21751
rect 3478 21687 3530 21693
rect 3490 20937 3518 21687
rect 3478 20931 3530 20937
rect 3478 20873 3530 20879
rect 3382 18563 3434 18569
rect 3382 18505 3434 18511
rect 3286 18415 3338 18421
rect 3202 18375 3286 18403
rect 3094 17749 3146 17755
rect 3094 17691 3146 17697
rect 3106 17607 3134 17691
rect 3094 17601 3146 17607
rect 3094 17543 3146 17549
rect 2998 17231 3050 17237
rect 2998 17173 3050 17179
rect 3106 16497 3134 17543
rect 3094 16491 3146 16497
rect 3094 16433 3146 16439
rect 3202 16349 3230 18375
rect 3286 18357 3338 18363
rect 3490 18273 3518 20873
rect 3478 18267 3530 18273
rect 3478 18209 3530 18215
rect 3586 17903 3614 22297
rect 3670 22279 3722 22285
rect 3778 21677 3806 22353
rect 3766 21671 3818 21677
rect 3766 21613 3818 21619
rect 3778 21085 3806 21613
rect 3766 21079 3818 21085
rect 3766 21021 3818 21027
rect 3670 18785 3722 18791
rect 3670 18727 3722 18733
rect 3574 17897 3626 17903
rect 3574 17839 3626 17845
rect 3682 16423 3710 18727
rect 3778 16941 3806 21021
rect 4258 20419 4286 22501
rect 4964 21340 5340 21349
rect 5020 21338 5044 21340
rect 5100 21338 5124 21340
rect 5180 21338 5204 21340
rect 5260 21338 5284 21340
rect 5020 21286 5030 21338
rect 5274 21286 5284 21338
rect 5020 21284 5044 21286
rect 5100 21284 5124 21286
rect 5180 21284 5204 21286
rect 5260 21284 5284 21286
rect 4964 21275 5340 21284
rect 4246 20413 4298 20419
rect 4246 20355 4298 20361
rect 4964 20008 5340 20017
rect 5020 20006 5044 20008
rect 5100 20006 5124 20008
rect 5180 20006 5204 20008
rect 5260 20006 5284 20008
rect 5020 19954 5030 20006
rect 5274 19954 5284 20006
rect 5020 19952 5044 19954
rect 5100 19952 5124 19954
rect 5180 19952 5204 19954
rect 5260 19952 5284 19954
rect 4964 19943 5340 19952
rect 4964 18676 5340 18685
rect 5020 18674 5044 18676
rect 5100 18674 5124 18676
rect 5180 18674 5204 18676
rect 5260 18674 5284 18676
rect 5020 18622 5030 18674
rect 5274 18622 5284 18674
rect 5020 18620 5044 18622
rect 5100 18620 5124 18622
rect 5180 18620 5204 18622
rect 5260 18620 5284 18622
rect 4964 18611 5340 18620
rect 4246 18415 4298 18421
rect 4246 18357 4298 18363
rect 4150 18341 4202 18347
rect 4150 18283 4202 18289
rect 4054 18193 4106 18199
rect 4054 18135 4106 18141
rect 4066 17755 4094 18135
rect 3862 17749 3914 17755
rect 3862 17691 3914 17697
rect 4054 17749 4106 17755
rect 4054 17691 4106 17697
rect 3766 16935 3818 16941
rect 3766 16877 3818 16883
rect 3670 16417 3722 16423
rect 3670 16359 3722 16365
rect 3190 16343 3242 16349
rect 3190 16285 3242 16291
rect 3682 15757 3710 16359
rect 3778 16275 3806 16877
rect 3766 16269 3818 16275
rect 3766 16211 3818 16217
rect 3670 15751 3722 15757
rect 3670 15693 3722 15699
rect 2914 13084 3038 13112
rect 2806 12939 2858 12945
rect 2806 12881 2858 12887
rect 2818 12427 2846 12881
rect 2806 12421 2858 12427
rect 2806 12363 2858 12369
rect 2614 11903 2666 11909
rect 2614 11845 2666 11851
rect 2626 11021 2654 11845
rect 2818 11539 2846 12363
rect 3010 12353 3038 13084
rect 2998 12347 3050 12353
rect 2998 12289 3050 12295
rect 3010 11761 3038 12289
rect 3682 12279 3710 15693
rect 3778 14277 3806 16211
rect 3874 15683 3902 17691
rect 3958 16935 4010 16941
rect 4066 16923 4094 17691
rect 4162 17681 4190 18283
rect 4258 17903 4286 18357
rect 4246 17897 4298 17903
rect 4246 17839 4298 17845
rect 4150 17675 4202 17681
rect 4150 17617 4202 17623
rect 4010 16895 4094 16923
rect 3958 16877 4010 16883
rect 3970 16497 3998 16877
rect 3958 16491 4010 16497
rect 3958 16433 4010 16439
rect 4162 16275 4190 17617
rect 4964 17344 5340 17353
rect 5020 17342 5044 17344
rect 5100 17342 5124 17344
rect 5180 17342 5204 17344
rect 5260 17342 5284 17344
rect 5020 17290 5030 17342
rect 5274 17290 5284 17342
rect 5020 17288 5044 17290
rect 5100 17288 5124 17290
rect 5180 17288 5204 17290
rect 5260 17288 5284 17290
rect 4964 17279 5340 17288
rect 5410 17015 5438 25387
rect 5794 23009 5822 25609
rect 5890 23897 5918 25609
rect 5878 23891 5930 23897
rect 5878 23833 5930 23839
rect 5782 23003 5834 23009
rect 5782 22945 5834 22951
rect 4630 17009 4682 17015
rect 4630 16951 4682 16957
rect 5398 17009 5450 17015
rect 5398 16951 5450 16957
rect 4438 16787 4490 16793
rect 4438 16729 4490 16735
rect 4450 16349 4478 16729
rect 4438 16343 4490 16349
rect 4438 16285 4490 16291
rect 4150 16269 4202 16275
rect 4150 16211 4202 16217
rect 3862 15677 3914 15683
rect 3862 15619 3914 15625
rect 3766 14271 3818 14277
rect 3766 14213 3818 14219
rect 4162 13019 4190 16211
rect 4642 13241 4670 16951
rect 5686 16787 5738 16793
rect 5686 16729 5738 16735
rect 4964 16012 5340 16021
rect 5020 16010 5044 16012
rect 5100 16010 5124 16012
rect 5180 16010 5204 16012
rect 5260 16010 5284 16012
rect 5020 15958 5030 16010
rect 5274 15958 5284 16010
rect 5020 15956 5044 15958
rect 5100 15956 5124 15958
rect 5180 15956 5204 15958
rect 5260 15956 5284 15958
rect 4964 15947 5340 15956
rect 4964 14680 5340 14689
rect 5020 14678 5044 14680
rect 5100 14678 5124 14680
rect 5180 14678 5204 14680
rect 5260 14678 5284 14680
rect 5020 14626 5030 14678
rect 5274 14626 5284 14678
rect 5020 14624 5044 14626
rect 5100 14624 5124 14626
rect 5180 14624 5204 14626
rect 5260 14624 5284 14626
rect 4964 14615 5340 14624
rect 4964 13348 5340 13357
rect 5020 13346 5044 13348
rect 5100 13346 5124 13348
rect 5180 13346 5204 13348
rect 5260 13346 5284 13348
rect 5020 13294 5030 13346
rect 5274 13294 5284 13346
rect 5020 13292 5044 13294
rect 5100 13292 5124 13294
rect 5180 13292 5204 13294
rect 5260 13292 5284 13294
rect 4964 13283 5340 13292
rect 4630 13235 4682 13241
rect 4630 13177 4682 13183
rect 4150 13013 4202 13019
rect 4150 12955 4202 12961
rect 4162 12353 4190 12955
rect 4642 12427 4670 13177
rect 5698 12575 5726 16729
rect 5986 16127 6014 25757
rect 6934 25667 6986 25673
rect 6934 25609 6986 25615
rect 7510 25667 7562 25673
rect 7510 25609 7562 25615
rect 8086 25667 8138 25673
rect 8086 25609 8138 25615
rect 9238 25667 9290 25673
rect 9238 25609 9290 25615
rect 6742 25519 6794 25525
rect 6742 25461 6794 25467
rect 6754 24489 6782 25461
rect 6946 25229 6974 25609
rect 7222 25593 7274 25599
rect 7222 25535 7274 25541
rect 6934 25223 6986 25229
rect 6934 25165 6986 25171
rect 6838 24927 6890 24933
rect 6838 24869 6890 24875
rect 6742 24483 6794 24489
rect 6742 24425 6794 24431
rect 6070 24409 6122 24415
rect 6070 24351 6122 24357
rect 6082 23601 6110 24351
rect 6754 24119 6782 24425
rect 6742 24113 6794 24119
rect 6742 24055 6794 24061
rect 6850 23916 6878 24869
rect 6754 23888 6878 23916
rect 6070 23595 6122 23601
rect 6070 23537 6122 23543
rect 6082 23083 6110 23537
rect 6070 23077 6122 23083
rect 6070 23019 6122 23025
rect 6082 22787 6110 23019
rect 6070 22781 6122 22787
rect 6070 22723 6122 22729
rect 6082 21751 6110 22723
rect 6070 21745 6122 21751
rect 6070 21687 6122 21693
rect 6754 21677 6782 23888
rect 7126 23003 7178 23009
rect 7126 22945 7178 22951
rect 6838 22929 6890 22935
rect 6838 22871 6890 22877
rect 6742 21671 6794 21677
rect 6742 21613 6794 21619
rect 6754 17294 6782 21613
rect 6658 17266 6782 17294
rect 5974 16121 6026 16127
rect 5974 16063 6026 16069
rect 5782 14271 5834 14277
rect 5782 14213 5834 14219
rect 5686 12569 5738 12575
rect 5686 12511 5738 12517
rect 4630 12421 4682 12427
rect 4630 12363 4682 12369
rect 4150 12347 4202 12353
rect 4150 12289 4202 12295
rect 3670 12273 3722 12279
rect 3670 12215 3722 12221
rect 3190 12125 3242 12131
rect 3190 12067 3242 12073
rect 2998 11755 3050 11761
rect 2998 11697 3050 11703
rect 2806 11533 2858 11539
rect 2806 11475 2858 11481
rect 2818 11095 2846 11475
rect 2806 11089 2858 11095
rect 2806 11031 2858 11037
rect 2614 11015 2666 11021
rect 2614 10957 2666 10963
rect 2902 7907 2954 7913
rect 2902 7849 2954 7855
rect 2710 7685 2762 7691
rect 2710 7627 2762 7633
rect 2722 7099 2750 7627
rect 2710 7093 2762 7099
rect 2710 7035 2762 7041
rect 2806 6871 2858 6877
rect 2806 6813 2858 6819
rect 2818 6507 2846 6813
rect 2914 6581 2942 7849
rect 2998 7463 3050 7469
rect 2998 7405 3050 7411
rect 3010 7173 3038 7405
rect 2998 7167 3050 7173
rect 2998 7109 3050 7115
rect 2902 6575 2954 6581
rect 2902 6517 2954 6523
rect 2806 6501 2858 6507
rect 2806 6443 2858 6449
rect 2518 3689 2570 3695
rect 2518 3631 2570 3637
rect 1846 3467 1898 3473
rect 1846 3409 1898 3415
rect 1462 3245 1514 3251
rect 1462 3187 1514 3193
rect 1558 3023 1610 3029
rect 1558 2965 1610 2971
rect 1570 1887 1598 2965
rect 1556 1878 1612 1887
rect 1556 1813 1612 1822
rect 596 0 652 800
rect 1748 680 1804 800
rect 1858 680 1886 3409
rect 1964 3358 2340 3367
rect 2020 3356 2044 3358
rect 2100 3356 2124 3358
rect 2180 3356 2204 3358
rect 2260 3356 2284 3358
rect 2020 3304 2030 3356
rect 2274 3304 2284 3356
rect 2020 3302 2044 3304
rect 2100 3302 2124 3304
rect 2180 3302 2204 3304
rect 2260 3302 2284 3304
rect 1964 3293 2340 3302
rect 3202 3029 3230 12067
rect 3682 11095 3710 12215
rect 4162 11687 4190 12289
rect 4150 11681 4202 11687
rect 4150 11623 4202 11629
rect 3670 11089 3722 11095
rect 3670 11031 3722 11037
rect 3682 10947 3710 11031
rect 3670 10941 3722 10947
rect 3670 10883 3722 10889
rect 3682 10429 3710 10883
rect 4162 10577 4190 11623
rect 4534 10793 4586 10799
rect 4534 10735 4586 10741
rect 4150 10571 4202 10577
rect 4150 10513 4202 10519
rect 3670 10423 3722 10429
rect 3670 10365 3722 10371
rect 4246 8351 4298 8357
rect 4246 8293 4298 8299
rect 3862 7685 3914 7691
rect 3862 7627 3914 7633
rect 3478 7611 3530 7617
rect 3478 7553 3530 7559
rect 3490 7247 3518 7553
rect 3478 7241 3530 7247
rect 3478 7183 3530 7189
rect 3874 6803 3902 7627
rect 4258 7214 4286 8293
rect 4258 7186 4382 7214
rect 4150 7167 4202 7173
rect 4150 7109 4202 7115
rect 4162 7025 4190 7109
rect 4150 7019 4202 7025
rect 4150 6961 4202 6967
rect 3286 6797 3338 6803
rect 3286 6739 3338 6745
rect 3862 6797 3914 6803
rect 3862 6739 3914 6745
rect 3958 6797 4010 6803
rect 3958 6739 4010 6745
rect 3298 6433 3326 6739
rect 3286 6427 3338 6433
rect 3286 6369 3338 6375
rect 3874 6359 3902 6739
rect 3862 6353 3914 6359
rect 3862 6295 3914 6301
rect 3874 6211 3902 6295
rect 3862 6205 3914 6211
rect 3862 6147 3914 6153
rect 3860 5874 3916 5883
rect 3970 5841 3998 6739
rect 3860 5809 3916 5818
rect 3958 5835 4010 5841
rect 3874 5693 3902 5809
rect 3958 5777 4010 5783
rect 3862 5687 3914 5693
rect 3862 5629 3914 5635
rect 3574 5465 3626 5471
rect 3574 5407 3626 5413
rect 3586 3769 3614 5407
rect 4162 5175 4190 6961
rect 4246 6131 4298 6137
rect 4246 6073 4298 6079
rect 4150 5169 4202 5175
rect 4150 5111 4202 5117
rect 4258 5101 4286 6073
rect 4354 5712 4382 7186
rect 4438 6945 4490 6951
rect 4438 6887 4490 6893
rect 4450 6137 4478 6887
rect 4438 6131 4490 6137
rect 4438 6073 4490 6079
rect 4546 5860 4574 10735
rect 4642 10355 4670 12363
rect 4964 12016 5340 12025
rect 5020 12014 5044 12016
rect 5100 12014 5124 12016
rect 5180 12014 5204 12016
rect 5260 12014 5284 12016
rect 5020 11962 5030 12014
rect 5274 11962 5284 12014
rect 5020 11960 5044 11962
rect 5100 11960 5124 11962
rect 5180 11960 5204 11962
rect 5260 11960 5284 11962
rect 4964 11951 5340 11960
rect 5698 11761 5726 12511
rect 5686 11755 5738 11761
rect 5686 11697 5738 11703
rect 5698 11021 5726 11697
rect 5686 11015 5738 11021
rect 5686 10957 5738 10963
rect 4964 10684 5340 10693
rect 5020 10682 5044 10684
rect 5100 10682 5124 10684
rect 5180 10682 5204 10684
rect 5260 10682 5284 10684
rect 5020 10630 5030 10682
rect 5274 10630 5284 10682
rect 5020 10628 5044 10630
rect 5100 10628 5124 10630
rect 5180 10628 5204 10630
rect 5260 10628 5284 10630
rect 4964 10619 5340 10628
rect 4630 10349 4682 10355
rect 4630 10291 4682 10297
rect 5590 10127 5642 10133
rect 5590 10069 5642 10075
rect 4964 9352 5340 9361
rect 5020 9350 5044 9352
rect 5100 9350 5124 9352
rect 5180 9350 5204 9352
rect 5260 9350 5284 9352
rect 5020 9298 5030 9350
rect 5274 9298 5284 9350
rect 5020 9296 5044 9298
rect 5100 9296 5124 9298
rect 5180 9296 5204 9298
rect 5260 9296 5284 9298
rect 4964 9287 5340 9296
rect 4964 8020 5340 8029
rect 5020 8018 5044 8020
rect 5100 8018 5124 8020
rect 5180 8018 5204 8020
rect 5260 8018 5284 8020
rect 5020 7966 5030 8018
rect 5274 7966 5284 8018
rect 5020 7964 5044 7966
rect 5100 7964 5124 7966
rect 5180 7964 5204 7966
rect 5260 7964 5284 7966
rect 4964 7955 5340 7964
rect 4630 7463 4682 7469
rect 4630 7405 4682 7411
rect 4642 7247 4670 7405
rect 4630 7241 4682 7247
rect 4630 7183 4682 7189
rect 4642 6581 4670 7183
rect 4726 7019 4778 7025
rect 4726 6961 4778 6967
rect 4630 6575 4682 6581
rect 4630 6517 4682 6523
rect 4546 5832 4670 5860
rect 4534 5761 4586 5767
rect 4354 5709 4534 5712
rect 4354 5703 4586 5709
rect 4354 5684 4574 5703
rect 4246 5095 4298 5101
rect 4246 5037 4298 5043
rect 3862 5021 3914 5027
rect 3862 4963 3914 4969
rect 3874 4435 3902 4963
rect 3862 4429 3914 4435
rect 3862 4371 3914 4377
rect 3574 3763 3626 3769
rect 3574 3705 3626 3711
rect 3874 3695 3902 4371
rect 4546 4361 4574 5684
rect 4534 4355 4586 4361
rect 4534 4297 4586 4303
rect 3862 3689 3914 3695
rect 3862 3631 3914 3637
rect 4642 3029 4670 5832
rect 4738 5249 4766 6961
rect 4822 6945 4874 6951
rect 4822 6887 4874 6893
rect 4834 6433 4862 6887
rect 5398 6797 5450 6803
rect 5398 6739 5450 6745
rect 4964 6688 5340 6697
rect 5020 6686 5044 6688
rect 5100 6686 5124 6688
rect 5180 6686 5204 6688
rect 5260 6686 5284 6688
rect 5020 6634 5030 6686
rect 5274 6634 5284 6686
rect 5020 6632 5044 6634
rect 5100 6632 5124 6634
rect 5180 6632 5204 6634
rect 5260 6632 5284 6634
rect 4964 6623 5340 6632
rect 4822 6427 4874 6433
rect 4822 6369 4874 6375
rect 4834 5471 4862 6369
rect 5110 6353 5162 6359
rect 5108 6318 5110 6327
rect 5162 6318 5164 6327
rect 5108 6253 5164 6262
rect 5122 5915 5150 6253
rect 5110 5909 5162 5915
rect 5110 5851 5162 5857
rect 4822 5465 4874 5471
rect 4822 5407 4874 5413
rect 4964 5356 5340 5365
rect 5020 5354 5044 5356
rect 5100 5354 5124 5356
rect 5180 5354 5204 5356
rect 5260 5354 5284 5356
rect 5020 5302 5030 5354
rect 5274 5302 5284 5354
rect 5020 5300 5044 5302
rect 5100 5300 5124 5302
rect 5180 5300 5204 5302
rect 5260 5300 5284 5302
rect 4964 5291 5340 5300
rect 4726 5243 4778 5249
rect 4726 5185 4778 5191
rect 5410 4953 5438 6739
rect 5494 6131 5546 6137
rect 5494 6073 5546 6079
rect 5506 5471 5534 6073
rect 5494 5465 5546 5471
rect 5494 5407 5546 5413
rect 5506 5101 5534 5407
rect 5494 5095 5546 5101
rect 5494 5037 5546 5043
rect 5398 4947 5450 4953
rect 5398 4889 5450 4895
rect 4964 4024 5340 4033
rect 5020 4022 5044 4024
rect 5100 4022 5124 4024
rect 5180 4022 5204 4024
rect 5260 4022 5284 4024
rect 5020 3970 5030 4022
rect 5274 3970 5284 4022
rect 5020 3968 5044 3970
rect 5100 3968 5124 3970
rect 5180 3968 5204 3970
rect 5260 3968 5284 3970
rect 4964 3959 5340 3968
rect 5506 3917 5534 5037
rect 5494 3911 5546 3917
rect 5494 3853 5546 3859
rect 5602 3029 5630 10069
rect 5794 7765 5822 14213
rect 6070 11533 6122 11539
rect 6070 11475 6122 11481
rect 6082 11243 6110 11475
rect 6070 11237 6122 11243
rect 6070 11179 6122 11185
rect 6550 10793 6602 10799
rect 6550 10735 6602 10741
rect 5878 10423 5930 10429
rect 5878 10365 5930 10371
rect 5890 8949 5918 10365
rect 6358 9609 6410 9615
rect 6358 9551 6410 9557
rect 5878 8943 5930 8949
rect 5878 8885 5930 8891
rect 5782 7759 5834 7765
rect 5782 7701 5834 7707
rect 5686 6945 5738 6951
rect 5686 6887 5738 6893
rect 5698 6507 5726 6887
rect 5686 6501 5738 6507
rect 5686 6443 5738 6449
rect 5794 6433 5822 7701
rect 6370 7025 6398 9551
rect 6358 7019 6410 7025
rect 6358 6961 6410 6967
rect 5782 6427 5834 6433
rect 5782 6369 5834 6375
rect 5686 5687 5738 5693
rect 5686 5629 5738 5635
rect 5698 5249 5726 5629
rect 5794 5249 5822 6369
rect 5878 5761 5930 5767
rect 5878 5703 5930 5709
rect 5890 5619 5918 5703
rect 5878 5613 5930 5619
rect 5878 5555 5930 5561
rect 5686 5243 5738 5249
rect 5686 5185 5738 5191
rect 5782 5243 5834 5249
rect 5782 5185 5834 5191
rect 5890 5175 5918 5555
rect 5878 5169 5930 5175
rect 5878 5111 5930 5117
rect 6562 3029 6590 10735
rect 6658 10429 6686 17266
rect 6742 16121 6794 16127
rect 6742 16063 6794 16069
rect 6754 15091 6782 16063
rect 6742 15085 6794 15091
rect 6742 15027 6794 15033
rect 6850 11169 6878 22871
rect 7138 22417 7166 22945
rect 7126 22411 7178 22417
rect 7126 22353 7178 22359
rect 7234 21899 7262 25535
rect 7522 25155 7550 25609
rect 7510 25149 7562 25155
rect 7510 25091 7562 25097
rect 8098 25081 8126 25609
rect 8086 25075 8138 25081
rect 8086 25017 8138 25023
rect 7964 24670 8340 24679
rect 8020 24668 8044 24670
rect 8100 24668 8124 24670
rect 8180 24668 8204 24670
rect 8260 24668 8284 24670
rect 8020 24616 8030 24668
rect 8274 24616 8284 24668
rect 8020 24614 8044 24616
rect 8100 24614 8124 24616
rect 8180 24614 8204 24616
rect 8260 24614 8284 24616
rect 7964 24605 8340 24614
rect 7798 24335 7850 24341
rect 7798 24277 7850 24283
rect 8470 24335 8522 24341
rect 8470 24277 8522 24283
rect 7810 22565 7838 24277
rect 8374 23669 8426 23675
rect 8374 23611 8426 23617
rect 7894 23595 7946 23601
rect 7894 23537 7946 23543
rect 7798 22559 7850 22565
rect 7798 22501 7850 22507
rect 7318 22337 7370 22343
rect 7318 22279 7370 22285
rect 7222 21893 7274 21899
rect 7222 21835 7274 21841
rect 7330 21011 7358 22279
rect 7906 22269 7934 23537
rect 7964 23338 8340 23347
rect 8020 23336 8044 23338
rect 8100 23336 8124 23338
rect 8180 23336 8204 23338
rect 8260 23336 8284 23338
rect 8020 23284 8030 23336
rect 8274 23284 8284 23336
rect 8020 23282 8044 23284
rect 8100 23282 8124 23284
rect 8180 23282 8204 23284
rect 8260 23282 8284 23284
rect 7964 23273 8340 23282
rect 8278 22929 8330 22935
rect 8386 22917 8414 23611
rect 8482 23527 8510 24277
rect 8566 24113 8618 24119
rect 8566 24055 8618 24061
rect 8470 23521 8522 23527
rect 8470 23463 8522 23469
rect 8330 22889 8414 22917
rect 8278 22871 8330 22877
rect 8290 22343 8318 22871
rect 8482 22732 8510 23463
rect 8386 22704 8510 22732
rect 8278 22337 8330 22343
rect 8278 22279 8330 22285
rect 7894 22263 7946 22269
rect 7894 22205 7946 22211
rect 7510 21893 7562 21899
rect 7510 21835 7562 21841
rect 7414 21227 7466 21233
rect 7414 21169 7466 21175
rect 7318 21005 7370 21011
rect 7318 20947 7370 20953
rect 7330 20271 7358 20947
rect 7318 20265 7370 20271
rect 7318 20207 7370 20213
rect 7330 19679 7358 20207
rect 7318 19673 7370 19679
rect 7318 19615 7370 19621
rect 7330 18347 7358 19615
rect 7318 18341 7370 18347
rect 7318 18283 7370 18289
rect 7426 14425 7454 21169
rect 7522 18421 7550 21835
rect 7906 20937 7934 22205
rect 7964 22006 8340 22015
rect 8020 22004 8044 22006
rect 8100 22004 8124 22006
rect 8180 22004 8204 22006
rect 8260 22004 8284 22006
rect 8020 21952 8030 22004
rect 8274 21952 8284 22004
rect 8020 21950 8044 21952
rect 8100 21950 8124 21952
rect 8180 21950 8204 21952
rect 8260 21950 8284 21952
rect 7964 21941 8340 21950
rect 7894 20931 7946 20937
rect 7894 20873 7946 20879
rect 7906 20419 7934 20873
rect 7964 20674 8340 20683
rect 8020 20672 8044 20674
rect 8100 20672 8124 20674
rect 8180 20672 8204 20674
rect 8260 20672 8284 20674
rect 8020 20620 8030 20672
rect 8274 20620 8284 20672
rect 8020 20618 8044 20620
rect 8100 20618 8124 20620
rect 8180 20618 8204 20620
rect 8260 20618 8284 20620
rect 7964 20609 8340 20618
rect 7894 20413 7946 20419
rect 7894 20355 7946 20361
rect 7906 19605 7934 20355
rect 7894 19599 7946 19605
rect 7894 19541 7946 19547
rect 7906 19476 7934 19541
rect 7810 19448 7934 19476
rect 7510 18415 7562 18421
rect 7510 18357 7562 18363
rect 7810 18273 7838 19448
rect 7964 19342 8340 19351
rect 8020 19340 8044 19342
rect 8100 19340 8124 19342
rect 8180 19340 8204 19342
rect 8260 19340 8284 19342
rect 8020 19288 8030 19340
rect 8274 19288 8284 19340
rect 8020 19286 8044 19288
rect 8100 19286 8124 19288
rect 8180 19286 8204 19288
rect 8260 19286 8284 19288
rect 7964 19277 8340 19286
rect 7894 18341 7946 18347
rect 7894 18283 7946 18289
rect 7798 18267 7850 18273
rect 7798 18209 7850 18215
rect 7810 18144 7838 18209
rect 7618 18116 7838 18144
rect 7618 16941 7646 18116
rect 7906 17015 7934 18283
rect 7964 18010 8340 18019
rect 8020 18008 8044 18010
rect 8100 18008 8124 18010
rect 8180 18008 8204 18010
rect 8260 18008 8284 18010
rect 8020 17956 8030 18008
rect 8274 17956 8284 18008
rect 8020 17954 8044 17956
rect 8100 17954 8124 17956
rect 8180 17954 8204 17956
rect 8260 17954 8284 17956
rect 7964 17945 8340 17954
rect 7894 17009 7946 17015
rect 7894 16951 7946 16957
rect 7606 16935 7658 16941
rect 7606 16877 7658 16883
rect 7618 15609 7646 16877
rect 7906 16571 7934 16951
rect 7964 16678 8340 16687
rect 8020 16676 8044 16678
rect 8100 16676 8124 16678
rect 8180 16676 8204 16678
rect 8260 16676 8284 16678
rect 8020 16624 8030 16676
rect 8274 16624 8284 16676
rect 8020 16622 8044 16624
rect 8100 16622 8124 16624
rect 8180 16622 8204 16624
rect 8260 16622 8284 16624
rect 7964 16613 8340 16622
rect 7894 16565 7946 16571
rect 7894 16507 7946 16513
rect 7906 15683 7934 16507
rect 8386 16275 8414 22704
rect 8470 22559 8522 22565
rect 8470 22501 8522 22507
rect 8374 16269 8426 16275
rect 8374 16211 8426 16217
rect 7894 15677 7946 15683
rect 7894 15619 7946 15625
rect 7606 15603 7658 15609
rect 7606 15545 7658 15551
rect 7618 15091 7646 15545
rect 7606 15085 7658 15091
rect 7606 15027 7658 15033
rect 7414 14419 7466 14425
rect 7414 14361 7466 14367
rect 7618 14277 7646 15027
rect 7906 15017 7934 15619
rect 7964 15346 8340 15355
rect 8020 15344 8044 15346
rect 8100 15344 8124 15346
rect 8180 15344 8204 15346
rect 8260 15344 8284 15346
rect 8020 15292 8030 15344
rect 8274 15292 8284 15344
rect 8020 15290 8044 15292
rect 8100 15290 8124 15292
rect 8180 15290 8204 15292
rect 8260 15290 8284 15292
rect 7964 15281 8340 15290
rect 7894 15011 7946 15017
rect 7894 14953 7946 14959
rect 7906 14351 7934 14953
rect 7894 14345 7946 14351
rect 7894 14287 7946 14293
rect 7606 14271 7658 14277
rect 7606 14213 7658 14219
rect 7964 14014 8340 14023
rect 8020 14012 8044 14014
rect 8100 14012 8124 14014
rect 8180 14012 8204 14014
rect 8260 14012 8284 14014
rect 8020 13960 8030 14012
rect 8274 13960 8284 14012
rect 8020 13958 8044 13960
rect 8100 13958 8124 13960
rect 8180 13958 8204 13960
rect 8260 13958 8284 13960
rect 7964 13949 8340 13958
rect 7964 12682 8340 12691
rect 8020 12680 8044 12682
rect 8100 12680 8124 12682
rect 8180 12680 8204 12682
rect 8260 12680 8284 12682
rect 8020 12628 8030 12680
rect 8274 12628 8284 12680
rect 8020 12626 8044 12628
rect 8100 12626 8124 12628
rect 8180 12626 8204 12628
rect 8260 12626 8284 12628
rect 7964 12617 8340 12626
rect 7510 12421 7562 12427
rect 7510 12363 7562 12369
rect 7126 11681 7178 11687
rect 7126 11623 7178 11629
rect 6838 11163 6890 11169
rect 6838 11105 6890 11111
rect 7138 11021 7166 11623
rect 7522 11613 7550 12363
rect 7510 11607 7562 11613
rect 7510 11549 7562 11555
rect 7522 11243 7550 11549
rect 7964 11350 8340 11359
rect 8020 11348 8044 11350
rect 8100 11348 8124 11350
rect 8180 11348 8204 11350
rect 8260 11348 8284 11350
rect 8020 11296 8030 11348
rect 8274 11296 8284 11348
rect 8020 11294 8044 11296
rect 8100 11294 8124 11296
rect 8180 11294 8204 11296
rect 8260 11294 8284 11296
rect 7964 11285 8340 11294
rect 8386 11243 8414 16211
rect 8482 11909 8510 22501
rect 8578 15757 8606 24055
rect 9250 16793 9278 25609
rect 9346 25229 9374 27269
rect 9634 25895 9662 28180
rect 10100 28074 10156 28874
rect 10676 28074 10732 28874
rect 11252 28074 11308 28874
rect 9622 25889 9674 25895
rect 9622 25831 9674 25837
rect 9718 25667 9770 25673
rect 9718 25609 9770 25615
rect 9334 25223 9386 25229
rect 9334 25165 9386 25171
rect 9334 25001 9386 25007
rect 9334 24943 9386 24949
rect 9430 25001 9482 25007
rect 9430 24943 9482 24949
rect 9346 23009 9374 24943
rect 9334 23003 9386 23009
rect 9334 22945 9386 22951
rect 9442 22787 9470 24943
rect 9730 24415 9758 25609
rect 10114 25229 10142 28074
rect 10102 25223 10154 25229
rect 10102 25165 10154 25171
rect 10690 25155 10718 28074
rect 10678 25149 10730 25155
rect 10678 25091 10730 25097
rect 11266 24489 11294 28074
rect 11254 24483 11306 24489
rect 11254 24425 11306 24431
rect 9718 24409 9770 24415
rect 9718 24351 9770 24357
rect 9814 23447 9866 23453
rect 9814 23389 9866 23395
rect 9826 23009 9854 23389
rect 9814 23003 9866 23009
rect 9814 22945 9866 22951
rect 9430 22781 9482 22787
rect 9430 22723 9482 22729
rect 10102 22781 10154 22787
rect 10102 22723 10154 22729
rect 10114 22607 10142 22723
rect 10100 22598 10156 22607
rect 10100 22533 10156 22542
rect 9814 22115 9866 22121
rect 9814 22057 9866 22063
rect 9718 20783 9770 20789
rect 9718 20725 9770 20731
rect 9334 20191 9386 20197
rect 9334 20133 9386 20139
rect 9238 16787 9290 16793
rect 9238 16729 9290 16735
rect 8566 15751 8618 15757
rect 8566 15693 8618 15699
rect 8470 11903 8522 11909
rect 8470 11845 8522 11851
rect 7510 11237 7562 11243
rect 7510 11179 7562 11185
rect 8374 11237 8426 11243
rect 8374 11179 8426 11185
rect 7522 11095 7550 11179
rect 8182 11163 8234 11169
rect 8182 11105 8234 11111
rect 7510 11089 7562 11095
rect 7510 11031 7562 11037
rect 7126 11015 7178 11021
rect 7126 10957 7178 10963
rect 6646 10423 6698 10429
rect 6646 10365 6698 10371
rect 6658 9911 6686 10365
rect 7138 10355 7166 10957
rect 7126 10349 7178 10355
rect 7126 10291 7178 10297
rect 7138 10004 7166 10291
rect 7522 10207 7550 11031
rect 8194 10577 8222 11105
rect 7798 10571 7850 10577
rect 7798 10513 7850 10519
rect 8182 10571 8234 10577
rect 8182 10513 8234 10519
rect 7510 10201 7562 10207
rect 7510 10143 7562 10149
rect 7042 9976 7166 10004
rect 6646 9905 6698 9911
rect 6646 9847 6698 9853
rect 7042 9689 7070 9976
rect 7126 9905 7178 9911
rect 7126 9847 7178 9853
rect 7030 9683 7082 9689
rect 7030 9625 7082 9631
rect 6742 8943 6794 8949
rect 6742 8885 6794 8891
rect 6754 8431 6782 8885
rect 6742 8425 6794 8431
rect 6742 8367 6794 8373
rect 6754 7765 6782 8367
rect 7138 8357 7166 9847
rect 7522 9763 7550 10143
rect 7510 9757 7562 9763
rect 7510 9699 7562 9705
rect 7522 8875 7550 9699
rect 7510 8869 7562 8875
rect 7510 8811 7562 8817
rect 7522 8431 7550 8811
rect 7510 8425 7562 8431
rect 7510 8367 7562 8373
rect 7126 8351 7178 8357
rect 7126 8293 7178 8299
rect 6742 7759 6794 7765
rect 6742 7701 6794 7707
rect 6754 6951 6782 7701
rect 7522 7617 7550 8367
rect 7810 7691 7838 10513
rect 7964 10018 8340 10027
rect 8020 10016 8044 10018
rect 8100 10016 8124 10018
rect 8180 10016 8204 10018
rect 8260 10016 8284 10018
rect 8020 9964 8030 10016
rect 8274 9964 8284 10016
rect 8020 9962 8044 9964
rect 8100 9962 8124 9964
rect 8180 9962 8204 9964
rect 8260 9962 8284 9964
rect 7964 9953 8340 9962
rect 8386 9023 8414 11179
rect 8482 9615 8510 11845
rect 8470 9609 8522 9615
rect 8470 9551 8522 9557
rect 8374 9017 8426 9023
rect 8374 8959 8426 8965
rect 7964 8686 8340 8695
rect 8020 8684 8044 8686
rect 8100 8684 8124 8686
rect 8180 8684 8204 8686
rect 8260 8684 8284 8686
rect 8020 8632 8030 8684
rect 8274 8632 8284 8684
rect 8020 8630 8044 8632
rect 8100 8630 8124 8632
rect 8180 8630 8204 8632
rect 8260 8630 8284 8632
rect 7964 8621 8340 8630
rect 9238 8129 9290 8135
rect 9238 8071 9290 8077
rect 7798 7685 7850 7691
rect 7798 7627 7850 7633
rect 7510 7611 7562 7617
rect 7510 7553 7562 7559
rect 7522 7247 7550 7553
rect 7964 7354 8340 7363
rect 8020 7352 8044 7354
rect 8100 7352 8124 7354
rect 8180 7352 8204 7354
rect 8260 7352 8284 7354
rect 8020 7300 8030 7352
rect 8274 7300 8284 7352
rect 8020 7298 8044 7300
rect 8100 7298 8124 7300
rect 8180 7298 8204 7300
rect 8260 7298 8284 7300
rect 7964 7289 8340 7298
rect 7510 7241 7562 7247
rect 7510 7183 7562 7189
rect 6742 6945 6794 6951
rect 6742 6887 6794 6893
rect 7894 6797 7946 6803
rect 7894 6739 7946 6745
rect 7906 3029 7934 6739
rect 7964 6022 8340 6031
rect 8020 6020 8044 6022
rect 8100 6020 8124 6022
rect 8180 6020 8204 6022
rect 8260 6020 8284 6022
rect 8020 5968 8030 6020
rect 8274 5968 8284 6020
rect 8020 5966 8044 5968
rect 8100 5966 8124 5968
rect 8180 5966 8204 5968
rect 8260 5966 8284 5968
rect 7964 5957 8340 5966
rect 7964 4690 8340 4699
rect 8020 4688 8044 4690
rect 8100 4688 8124 4690
rect 8180 4688 8204 4690
rect 8260 4688 8284 4690
rect 8020 4636 8030 4688
rect 8274 4636 8284 4688
rect 8020 4634 8044 4636
rect 8100 4634 8124 4636
rect 8180 4634 8204 4636
rect 8260 4634 8284 4636
rect 7964 4625 8340 4634
rect 7964 3358 8340 3367
rect 8020 3356 8044 3358
rect 8100 3356 8124 3358
rect 8180 3356 8204 3358
rect 8260 3356 8284 3358
rect 8020 3304 8030 3356
rect 8274 3304 8284 3356
rect 8020 3302 8044 3304
rect 8100 3302 8124 3304
rect 8180 3302 8204 3304
rect 8260 3302 8284 3304
rect 7964 3293 8340 3302
rect 9250 3029 9278 8071
rect 9346 3029 9374 20133
rect 9622 16787 9674 16793
rect 9622 16729 9674 16735
rect 9430 14123 9482 14129
rect 9430 14065 9482 14071
rect 9442 8357 9470 14065
rect 9634 11021 9662 16729
rect 9622 11015 9674 11021
rect 9622 10957 9674 10963
rect 9526 8795 9578 8801
rect 9526 8737 9578 8743
rect 9430 8351 9482 8357
rect 9430 8293 9482 8299
rect 9538 3695 9566 8737
rect 9622 7463 9674 7469
rect 9622 7405 9674 7411
rect 9526 3689 9578 3695
rect 9526 3631 9578 3637
rect 9634 3029 9662 7405
rect 9730 6359 9758 20725
rect 9826 20345 9854 22057
rect 9814 20339 9866 20345
rect 9814 20281 9866 20287
rect 10100 20230 10156 20239
rect 10100 20165 10102 20174
rect 10154 20165 10156 20174
rect 10102 20133 10154 20139
rect 9910 19451 9962 19457
rect 9910 19393 9962 19399
rect 9814 14789 9866 14795
rect 9814 14731 9866 14737
rect 9826 13685 9854 14731
rect 9814 13679 9866 13685
rect 9814 13621 9866 13627
rect 9718 6353 9770 6359
rect 9718 6295 9770 6301
rect 9922 3695 9950 19393
rect 10102 18119 10154 18125
rect 10102 18061 10154 18067
rect 10114 17871 10142 18061
rect 10100 17862 10156 17871
rect 10100 17797 10156 17806
rect 10100 15494 10156 15503
rect 10100 15429 10102 15438
rect 10154 15429 10156 15438
rect 10102 15397 10154 15403
rect 10102 13457 10154 13463
rect 10102 13399 10154 13405
rect 10114 13135 10142 13399
rect 10100 13126 10156 13135
rect 10100 13061 10156 13070
rect 10102 10793 10154 10799
rect 10100 10758 10102 10767
rect 10154 10758 10156 10767
rect 10100 10693 10156 10702
rect 10100 8390 10156 8399
rect 10100 8325 10102 8334
rect 10154 8325 10156 8334
rect 10102 8293 10154 8299
rect 10102 6131 10154 6137
rect 10102 6073 10154 6079
rect 10114 6031 10142 6073
rect 10100 6022 10156 6031
rect 10100 5957 10156 5966
rect 9910 3689 9962 3695
rect 9910 3631 9962 3637
rect 10100 3654 10156 3663
rect 10100 3589 10102 3598
rect 10154 3589 10156 3598
rect 10102 3557 10154 3563
rect 10966 3467 11018 3473
rect 10966 3409 11018 3415
rect 3190 3023 3242 3029
rect 3190 2965 3242 2971
rect 4630 3023 4682 3029
rect 4630 2965 4682 2971
rect 5590 3023 5642 3029
rect 5590 2965 5642 2971
rect 6550 3023 6602 3029
rect 6550 2965 6602 2971
rect 7894 3023 7946 3029
rect 7894 2965 7946 2971
rect 9238 3023 9290 3029
rect 9238 2965 9290 2971
rect 9334 3023 9386 3029
rect 9334 2965 9386 2971
rect 9622 3023 9674 3029
rect 9622 2965 9674 2971
rect 2902 2949 2954 2955
rect 2902 2891 2954 2897
rect 4054 2949 4106 2955
rect 4054 2891 4106 2897
rect 5398 2949 5450 2955
rect 5398 2891 5450 2897
rect 6358 2949 6410 2955
rect 6358 2891 6410 2897
rect 7606 2949 7658 2955
rect 7606 2891 7658 2897
rect 8662 2949 8714 2955
rect 8662 2891 8714 2897
rect 9718 2949 9770 2955
rect 9718 2891 9770 2897
rect 9814 2949 9866 2955
rect 9814 2891 9866 2897
rect 2914 800 2942 2891
rect 4066 800 4094 2891
rect 4964 2692 5340 2701
rect 5020 2690 5044 2692
rect 5100 2690 5124 2692
rect 5180 2690 5204 2692
rect 5260 2690 5284 2692
rect 5020 2638 5030 2690
rect 5274 2638 5284 2690
rect 5020 2636 5044 2638
rect 5100 2636 5124 2638
rect 5180 2636 5204 2638
rect 5260 2636 5284 2638
rect 4964 2627 5340 2636
rect 5410 1420 5438 2891
rect 5218 1392 5438 1420
rect 5218 800 5246 1392
rect 6370 800 6398 2891
rect 1748 652 1886 680
rect 1748 0 1804 652
rect 2900 0 2956 800
rect 4052 0 4108 800
rect 5204 0 5260 800
rect 6356 0 6412 800
rect 7508 680 7564 800
rect 7618 680 7646 2891
rect 8674 800 8702 2891
rect 9730 1295 9758 2891
rect 9716 1286 9772 1295
rect 9716 1221 9772 1230
rect 9826 800 9854 2891
rect 10978 800 11006 3409
rect 7508 652 7646 680
rect 7508 0 7564 652
rect 8660 0 8716 800
rect 9812 0 9868 800
rect 10964 0 11020 800
<< via2 >>
rect 1460 26686 1516 26742
rect 1964 26000 2020 26002
rect 2044 26000 2100 26002
rect 2124 26000 2180 26002
rect 2204 26000 2260 26002
rect 2284 26000 2340 26002
rect 1964 25948 1966 26000
rect 1966 25948 2018 26000
rect 2018 25948 2020 26000
rect 2044 25948 2082 26000
rect 2082 25948 2094 26000
rect 2094 25948 2100 26000
rect 2124 25948 2146 26000
rect 2146 25948 2158 26000
rect 2158 25948 2180 26000
rect 2204 25948 2210 26000
rect 2210 25948 2222 26000
rect 2222 25948 2260 26000
rect 2284 25948 2286 26000
rect 2286 25948 2338 26000
rect 2338 25948 2340 26000
rect 1964 25946 2020 25948
rect 2044 25946 2100 25948
rect 2124 25946 2180 25948
rect 2204 25946 2260 25948
rect 2284 25946 2340 25948
rect 7964 26000 8020 26002
rect 8044 26000 8100 26002
rect 8124 26000 8180 26002
rect 8204 26000 8260 26002
rect 8284 26000 8340 26002
rect 7964 25948 7966 26000
rect 7966 25948 8018 26000
rect 8018 25948 8020 26000
rect 8044 25948 8082 26000
rect 8082 25948 8094 26000
rect 8094 25948 8100 26000
rect 8124 25948 8146 26000
rect 8146 25948 8158 26000
rect 8158 25948 8180 26000
rect 8204 25948 8210 26000
rect 8210 25948 8222 26000
rect 8222 25948 8260 26000
rect 8284 25948 8286 26000
rect 8286 25948 8338 26000
rect 8338 25948 8340 26000
rect 7964 25946 8020 25948
rect 8044 25946 8100 25948
rect 8124 25946 8180 25948
rect 8204 25946 8260 25948
rect 8284 25946 8340 25948
rect 9332 27278 9388 27334
rect 1268 22559 1324 22598
rect 1268 22542 1270 22559
rect 1270 22542 1322 22559
rect 1322 22542 1324 22559
rect 1652 18398 1708 18454
rect 884 14271 940 14310
rect 884 14254 886 14271
rect 886 14254 938 14271
rect 938 14254 940 14271
rect 884 10110 940 10166
rect 1964 24668 2020 24670
rect 2044 24668 2100 24670
rect 2124 24668 2180 24670
rect 2204 24668 2260 24670
rect 2284 24668 2340 24670
rect 1964 24616 1966 24668
rect 1966 24616 2018 24668
rect 2018 24616 2020 24668
rect 2044 24616 2082 24668
rect 2082 24616 2094 24668
rect 2094 24616 2100 24668
rect 2124 24616 2146 24668
rect 2146 24616 2158 24668
rect 2158 24616 2180 24668
rect 2204 24616 2210 24668
rect 2210 24616 2222 24668
rect 2222 24616 2260 24668
rect 2284 24616 2286 24668
rect 2286 24616 2338 24668
rect 2338 24616 2340 24668
rect 1964 24614 2020 24616
rect 2044 24614 2100 24616
rect 2124 24614 2180 24616
rect 2204 24614 2260 24616
rect 2284 24614 2340 24616
rect 1964 23336 2020 23338
rect 2044 23336 2100 23338
rect 2124 23336 2180 23338
rect 2204 23336 2260 23338
rect 2284 23336 2340 23338
rect 1964 23284 1966 23336
rect 1966 23284 2018 23336
rect 2018 23284 2020 23336
rect 2044 23284 2082 23336
rect 2082 23284 2094 23336
rect 2094 23284 2100 23336
rect 2124 23284 2146 23336
rect 2146 23284 2158 23336
rect 2158 23284 2180 23336
rect 2204 23284 2210 23336
rect 2210 23284 2222 23336
rect 2222 23284 2260 23336
rect 2284 23284 2286 23336
rect 2286 23284 2338 23336
rect 2338 23284 2340 23336
rect 1964 23282 2020 23284
rect 2044 23282 2100 23284
rect 2124 23282 2180 23284
rect 2204 23282 2260 23284
rect 2284 23282 2340 23284
rect 1964 22004 2020 22006
rect 2044 22004 2100 22006
rect 2124 22004 2180 22006
rect 2204 22004 2260 22006
rect 2284 22004 2340 22006
rect 1964 21952 1966 22004
rect 1966 21952 2018 22004
rect 2018 21952 2020 22004
rect 2044 21952 2082 22004
rect 2082 21952 2094 22004
rect 2094 21952 2100 22004
rect 2124 21952 2146 22004
rect 2146 21952 2158 22004
rect 2158 21952 2180 22004
rect 2204 21952 2210 22004
rect 2210 21952 2222 22004
rect 2222 21952 2260 22004
rect 2284 21952 2286 22004
rect 2286 21952 2338 22004
rect 2338 21952 2340 22004
rect 1964 21950 2020 21952
rect 2044 21950 2100 21952
rect 2124 21950 2180 21952
rect 2204 21950 2260 21952
rect 2284 21950 2340 21952
rect 1964 20672 2020 20674
rect 2044 20672 2100 20674
rect 2124 20672 2180 20674
rect 2204 20672 2260 20674
rect 2284 20672 2340 20674
rect 1964 20620 1966 20672
rect 1966 20620 2018 20672
rect 2018 20620 2020 20672
rect 2044 20620 2082 20672
rect 2082 20620 2094 20672
rect 2094 20620 2100 20672
rect 2124 20620 2146 20672
rect 2146 20620 2158 20672
rect 2158 20620 2180 20672
rect 2204 20620 2210 20672
rect 2210 20620 2222 20672
rect 2222 20620 2260 20672
rect 2284 20620 2286 20672
rect 2286 20620 2338 20672
rect 2338 20620 2340 20672
rect 1964 20618 2020 20620
rect 2044 20618 2100 20620
rect 2124 20618 2180 20620
rect 2204 20618 2260 20620
rect 2284 20618 2340 20620
rect 1964 19340 2020 19342
rect 2044 19340 2100 19342
rect 2124 19340 2180 19342
rect 2204 19340 2260 19342
rect 2284 19340 2340 19342
rect 1964 19288 1966 19340
rect 1966 19288 2018 19340
rect 2018 19288 2020 19340
rect 2044 19288 2082 19340
rect 2082 19288 2094 19340
rect 2094 19288 2100 19340
rect 2124 19288 2146 19340
rect 2146 19288 2158 19340
rect 2158 19288 2180 19340
rect 2204 19288 2210 19340
rect 2210 19288 2222 19340
rect 2222 19288 2260 19340
rect 2284 19288 2286 19340
rect 2286 19288 2338 19340
rect 2338 19288 2340 19340
rect 1964 19286 2020 19288
rect 2044 19286 2100 19288
rect 2124 19286 2180 19288
rect 2204 19286 2260 19288
rect 2284 19286 2340 19288
rect 1964 18008 2020 18010
rect 2044 18008 2100 18010
rect 2124 18008 2180 18010
rect 2204 18008 2260 18010
rect 2284 18008 2340 18010
rect 1964 17956 1966 18008
rect 1966 17956 2018 18008
rect 2018 17956 2020 18008
rect 2044 17956 2082 18008
rect 2082 17956 2094 18008
rect 2094 17956 2100 18008
rect 2124 17956 2146 18008
rect 2146 17956 2158 18008
rect 2158 17956 2180 18008
rect 2204 17956 2210 18008
rect 2210 17956 2222 18008
rect 2222 17956 2260 18008
rect 2284 17956 2286 18008
rect 2286 17956 2338 18008
rect 2338 17956 2340 18008
rect 1964 17954 2020 17956
rect 2044 17954 2100 17956
rect 2124 17954 2180 17956
rect 2204 17954 2260 17956
rect 2284 17954 2340 17956
rect 1964 16676 2020 16678
rect 2044 16676 2100 16678
rect 2124 16676 2180 16678
rect 2204 16676 2260 16678
rect 2284 16676 2340 16678
rect 1964 16624 1966 16676
rect 1966 16624 2018 16676
rect 2018 16624 2020 16676
rect 2044 16624 2082 16676
rect 2082 16624 2094 16676
rect 2094 16624 2100 16676
rect 2124 16624 2146 16676
rect 2146 16624 2158 16676
rect 2158 16624 2180 16676
rect 2204 16624 2210 16676
rect 2210 16624 2222 16676
rect 2222 16624 2260 16676
rect 2284 16624 2286 16676
rect 2286 16624 2338 16676
rect 2338 16624 2340 16676
rect 1964 16622 2020 16624
rect 2044 16622 2100 16624
rect 2124 16622 2180 16624
rect 2204 16622 2260 16624
rect 2284 16622 2340 16624
rect 1964 15344 2020 15346
rect 2044 15344 2100 15346
rect 2124 15344 2180 15346
rect 2204 15344 2260 15346
rect 2284 15344 2340 15346
rect 1964 15292 1966 15344
rect 1966 15292 2018 15344
rect 2018 15292 2020 15344
rect 2044 15292 2082 15344
rect 2082 15292 2094 15344
rect 2094 15292 2100 15344
rect 2124 15292 2146 15344
rect 2146 15292 2158 15344
rect 2158 15292 2180 15344
rect 2204 15292 2210 15344
rect 2210 15292 2222 15344
rect 2222 15292 2260 15344
rect 2284 15292 2286 15344
rect 2286 15292 2338 15344
rect 2338 15292 2340 15344
rect 1964 15290 2020 15292
rect 2044 15290 2100 15292
rect 2124 15290 2180 15292
rect 2204 15290 2260 15292
rect 2284 15290 2340 15292
rect 1964 14012 2020 14014
rect 2044 14012 2100 14014
rect 2124 14012 2180 14014
rect 2204 14012 2260 14014
rect 2284 14012 2340 14014
rect 1964 13960 1966 14012
rect 1966 13960 2018 14012
rect 2018 13960 2020 14012
rect 2044 13960 2082 14012
rect 2082 13960 2094 14012
rect 2094 13960 2100 14012
rect 2124 13960 2146 14012
rect 2146 13960 2158 14012
rect 2158 13960 2180 14012
rect 2204 13960 2210 14012
rect 2210 13960 2222 14012
rect 2222 13960 2260 14012
rect 2284 13960 2286 14012
rect 2286 13960 2338 14012
rect 2338 13960 2340 14012
rect 1964 13958 2020 13960
rect 2044 13958 2100 13960
rect 2124 13958 2180 13960
rect 2204 13958 2260 13960
rect 2284 13958 2340 13960
rect 1964 12680 2020 12682
rect 2044 12680 2100 12682
rect 2124 12680 2180 12682
rect 2204 12680 2260 12682
rect 2284 12680 2340 12682
rect 1964 12628 1966 12680
rect 1966 12628 2018 12680
rect 2018 12628 2020 12680
rect 2044 12628 2082 12680
rect 2082 12628 2094 12680
rect 2094 12628 2100 12680
rect 2124 12628 2146 12680
rect 2146 12628 2158 12680
rect 2158 12628 2180 12680
rect 2204 12628 2210 12680
rect 2210 12628 2222 12680
rect 2222 12628 2260 12680
rect 2284 12628 2286 12680
rect 2286 12628 2338 12680
rect 2338 12628 2340 12680
rect 1964 12626 2020 12628
rect 2044 12626 2100 12628
rect 2124 12626 2180 12628
rect 2204 12626 2260 12628
rect 2284 12626 2340 12628
rect 1964 11348 2020 11350
rect 2044 11348 2100 11350
rect 2124 11348 2180 11350
rect 2204 11348 2260 11350
rect 2284 11348 2340 11350
rect 1964 11296 1966 11348
rect 1966 11296 2018 11348
rect 2018 11296 2020 11348
rect 2044 11296 2082 11348
rect 2082 11296 2094 11348
rect 2094 11296 2100 11348
rect 2124 11296 2146 11348
rect 2146 11296 2158 11348
rect 2158 11296 2180 11348
rect 2204 11296 2210 11348
rect 2210 11296 2222 11348
rect 2222 11296 2260 11348
rect 2284 11296 2286 11348
rect 2286 11296 2338 11348
rect 2338 11296 2340 11348
rect 1964 11294 2020 11296
rect 2044 11294 2100 11296
rect 2124 11294 2180 11296
rect 2204 11294 2260 11296
rect 2284 11294 2340 11296
rect 1964 10016 2020 10018
rect 2044 10016 2100 10018
rect 2124 10016 2180 10018
rect 2204 10016 2260 10018
rect 2284 10016 2340 10018
rect 1964 9964 1966 10016
rect 1966 9964 2018 10016
rect 2018 9964 2020 10016
rect 2044 9964 2082 10016
rect 2082 9964 2094 10016
rect 2094 9964 2100 10016
rect 2124 9964 2146 10016
rect 2146 9964 2158 10016
rect 2158 9964 2180 10016
rect 2204 9964 2210 10016
rect 2210 9964 2222 10016
rect 2222 9964 2260 10016
rect 2284 9964 2286 10016
rect 2286 9964 2338 10016
rect 2338 9964 2340 10016
rect 1964 9962 2020 9964
rect 2044 9962 2100 9964
rect 2124 9962 2180 9964
rect 2204 9962 2260 9964
rect 2284 9962 2340 9964
rect 1964 8684 2020 8686
rect 2044 8684 2100 8686
rect 2124 8684 2180 8686
rect 2204 8684 2260 8686
rect 2284 8684 2340 8686
rect 1964 8632 1966 8684
rect 1966 8632 2018 8684
rect 2018 8632 2020 8684
rect 2044 8632 2082 8684
rect 2082 8632 2094 8684
rect 2094 8632 2100 8684
rect 2124 8632 2146 8684
rect 2146 8632 2158 8684
rect 2158 8632 2180 8684
rect 2204 8632 2210 8684
rect 2210 8632 2222 8684
rect 2222 8632 2260 8684
rect 2284 8632 2286 8684
rect 2286 8632 2338 8684
rect 2338 8632 2340 8684
rect 1964 8630 2020 8632
rect 2044 8630 2100 8632
rect 2124 8630 2180 8632
rect 2204 8630 2260 8632
rect 2284 8630 2340 8632
rect 1964 7352 2020 7354
rect 2044 7352 2100 7354
rect 2124 7352 2180 7354
rect 2204 7352 2260 7354
rect 2284 7352 2340 7354
rect 1964 7300 1966 7352
rect 1966 7300 2018 7352
rect 2018 7300 2020 7352
rect 2044 7300 2082 7352
rect 2082 7300 2094 7352
rect 2094 7300 2100 7352
rect 2124 7300 2146 7352
rect 2146 7300 2158 7352
rect 2158 7300 2180 7352
rect 2204 7300 2210 7352
rect 2210 7300 2222 7352
rect 2222 7300 2260 7352
rect 2284 7300 2286 7352
rect 2286 7300 2338 7352
rect 2338 7300 2340 7352
rect 1964 7298 2020 7300
rect 2044 7298 2100 7300
rect 2124 7298 2180 7300
rect 2204 7298 2260 7300
rect 2284 7298 2340 7300
rect 1748 6301 1750 6318
rect 1750 6301 1802 6318
rect 1802 6301 1804 6318
rect 1748 6262 1804 6301
rect 1964 6020 2020 6022
rect 2044 6020 2100 6022
rect 2124 6020 2180 6022
rect 2204 6020 2260 6022
rect 2284 6020 2340 6022
rect 1964 5968 1966 6020
rect 1966 5968 2018 6020
rect 2018 5968 2020 6020
rect 2044 5968 2082 6020
rect 2082 5968 2094 6020
rect 2094 5968 2100 6020
rect 2124 5968 2146 6020
rect 2146 5968 2158 6020
rect 2158 5968 2180 6020
rect 2204 5968 2210 6020
rect 2210 5968 2222 6020
rect 2222 5968 2260 6020
rect 2284 5968 2286 6020
rect 2286 5968 2338 6020
rect 2338 5968 2340 6020
rect 1964 5966 2020 5968
rect 2044 5966 2100 5968
rect 2124 5966 2180 5968
rect 2204 5966 2260 5968
rect 2284 5966 2340 5968
rect 1964 4688 2020 4690
rect 2044 4688 2100 4690
rect 2124 4688 2180 4690
rect 2204 4688 2260 4690
rect 2284 4688 2340 4690
rect 1964 4636 1966 4688
rect 1966 4636 2018 4688
rect 2018 4636 2020 4688
rect 2044 4636 2082 4688
rect 2082 4636 2094 4688
rect 2094 4636 2100 4688
rect 2124 4636 2146 4688
rect 2146 4636 2158 4688
rect 2158 4636 2180 4688
rect 2204 4636 2210 4688
rect 2210 4636 2222 4688
rect 2222 4636 2260 4688
rect 2284 4636 2286 4688
rect 2286 4636 2338 4688
rect 2338 4636 2340 4688
rect 1964 4634 2020 4636
rect 2044 4634 2100 4636
rect 2124 4634 2180 4636
rect 2204 4634 2260 4636
rect 2284 4634 2340 4636
rect 4964 25334 5020 25336
rect 5044 25334 5100 25336
rect 5124 25334 5180 25336
rect 5204 25334 5260 25336
rect 5284 25334 5340 25336
rect 4964 25282 4966 25334
rect 4966 25282 5018 25334
rect 5018 25282 5020 25334
rect 5044 25282 5082 25334
rect 5082 25282 5094 25334
rect 5094 25282 5100 25334
rect 5124 25282 5146 25334
rect 5146 25282 5158 25334
rect 5158 25282 5180 25334
rect 5204 25282 5210 25334
rect 5210 25282 5222 25334
rect 5222 25282 5260 25334
rect 5284 25282 5286 25334
rect 5286 25282 5338 25334
rect 5338 25282 5340 25334
rect 4964 25280 5020 25282
rect 5044 25280 5100 25282
rect 5124 25280 5180 25282
rect 5204 25280 5260 25282
rect 5284 25280 5340 25282
rect 4964 24002 5020 24004
rect 5044 24002 5100 24004
rect 5124 24002 5180 24004
rect 5204 24002 5260 24004
rect 5284 24002 5340 24004
rect 4964 23950 4966 24002
rect 4966 23950 5018 24002
rect 5018 23950 5020 24002
rect 5044 23950 5082 24002
rect 5082 23950 5094 24002
rect 5094 23950 5100 24002
rect 5124 23950 5146 24002
rect 5146 23950 5158 24002
rect 5158 23950 5180 24002
rect 5204 23950 5210 24002
rect 5210 23950 5222 24002
rect 5222 23950 5260 24002
rect 5284 23950 5286 24002
rect 5286 23950 5338 24002
rect 5338 23950 5340 24002
rect 4964 23948 5020 23950
rect 5044 23948 5100 23950
rect 5124 23948 5180 23950
rect 5204 23948 5260 23950
rect 5284 23948 5340 23950
rect 4964 22670 5020 22672
rect 5044 22670 5100 22672
rect 5124 22670 5180 22672
rect 5204 22670 5260 22672
rect 5284 22670 5340 22672
rect 4964 22618 4966 22670
rect 4966 22618 5018 22670
rect 5018 22618 5020 22670
rect 5044 22618 5082 22670
rect 5082 22618 5094 22670
rect 5094 22618 5100 22670
rect 5124 22618 5146 22670
rect 5146 22618 5158 22670
rect 5158 22618 5180 22670
rect 5204 22618 5210 22670
rect 5210 22618 5222 22670
rect 5222 22618 5260 22670
rect 5284 22618 5286 22670
rect 5286 22618 5338 22670
rect 5338 22618 5340 22670
rect 4964 22616 5020 22618
rect 5044 22616 5100 22618
rect 5124 22616 5180 22618
rect 5204 22616 5260 22618
rect 5284 22616 5340 22618
rect 4964 21338 5020 21340
rect 5044 21338 5100 21340
rect 5124 21338 5180 21340
rect 5204 21338 5260 21340
rect 5284 21338 5340 21340
rect 4964 21286 4966 21338
rect 4966 21286 5018 21338
rect 5018 21286 5020 21338
rect 5044 21286 5082 21338
rect 5082 21286 5094 21338
rect 5094 21286 5100 21338
rect 5124 21286 5146 21338
rect 5146 21286 5158 21338
rect 5158 21286 5180 21338
rect 5204 21286 5210 21338
rect 5210 21286 5222 21338
rect 5222 21286 5260 21338
rect 5284 21286 5286 21338
rect 5286 21286 5338 21338
rect 5338 21286 5340 21338
rect 4964 21284 5020 21286
rect 5044 21284 5100 21286
rect 5124 21284 5180 21286
rect 5204 21284 5260 21286
rect 5284 21284 5340 21286
rect 4964 20006 5020 20008
rect 5044 20006 5100 20008
rect 5124 20006 5180 20008
rect 5204 20006 5260 20008
rect 5284 20006 5340 20008
rect 4964 19954 4966 20006
rect 4966 19954 5018 20006
rect 5018 19954 5020 20006
rect 5044 19954 5082 20006
rect 5082 19954 5094 20006
rect 5094 19954 5100 20006
rect 5124 19954 5146 20006
rect 5146 19954 5158 20006
rect 5158 19954 5180 20006
rect 5204 19954 5210 20006
rect 5210 19954 5222 20006
rect 5222 19954 5260 20006
rect 5284 19954 5286 20006
rect 5286 19954 5338 20006
rect 5338 19954 5340 20006
rect 4964 19952 5020 19954
rect 5044 19952 5100 19954
rect 5124 19952 5180 19954
rect 5204 19952 5260 19954
rect 5284 19952 5340 19954
rect 4964 18674 5020 18676
rect 5044 18674 5100 18676
rect 5124 18674 5180 18676
rect 5204 18674 5260 18676
rect 5284 18674 5340 18676
rect 4964 18622 4966 18674
rect 4966 18622 5018 18674
rect 5018 18622 5020 18674
rect 5044 18622 5082 18674
rect 5082 18622 5094 18674
rect 5094 18622 5100 18674
rect 5124 18622 5146 18674
rect 5146 18622 5158 18674
rect 5158 18622 5180 18674
rect 5204 18622 5210 18674
rect 5210 18622 5222 18674
rect 5222 18622 5260 18674
rect 5284 18622 5286 18674
rect 5286 18622 5338 18674
rect 5338 18622 5340 18674
rect 4964 18620 5020 18622
rect 5044 18620 5100 18622
rect 5124 18620 5180 18622
rect 5204 18620 5260 18622
rect 5284 18620 5340 18622
rect 4964 17342 5020 17344
rect 5044 17342 5100 17344
rect 5124 17342 5180 17344
rect 5204 17342 5260 17344
rect 5284 17342 5340 17344
rect 4964 17290 4966 17342
rect 4966 17290 5018 17342
rect 5018 17290 5020 17342
rect 5044 17290 5082 17342
rect 5082 17290 5094 17342
rect 5094 17290 5100 17342
rect 5124 17290 5146 17342
rect 5146 17290 5158 17342
rect 5158 17290 5180 17342
rect 5204 17290 5210 17342
rect 5210 17290 5222 17342
rect 5222 17290 5260 17342
rect 5284 17290 5286 17342
rect 5286 17290 5338 17342
rect 5338 17290 5340 17342
rect 4964 17288 5020 17290
rect 5044 17288 5100 17290
rect 5124 17288 5180 17290
rect 5204 17288 5260 17290
rect 5284 17288 5340 17290
rect 4964 16010 5020 16012
rect 5044 16010 5100 16012
rect 5124 16010 5180 16012
rect 5204 16010 5260 16012
rect 5284 16010 5340 16012
rect 4964 15958 4966 16010
rect 4966 15958 5018 16010
rect 5018 15958 5020 16010
rect 5044 15958 5082 16010
rect 5082 15958 5094 16010
rect 5094 15958 5100 16010
rect 5124 15958 5146 16010
rect 5146 15958 5158 16010
rect 5158 15958 5180 16010
rect 5204 15958 5210 16010
rect 5210 15958 5222 16010
rect 5222 15958 5260 16010
rect 5284 15958 5286 16010
rect 5286 15958 5338 16010
rect 5338 15958 5340 16010
rect 4964 15956 5020 15958
rect 5044 15956 5100 15958
rect 5124 15956 5180 15958
rect 5204 15956 5260 15958
rect 5284 15956 5340 15958
rect 4964 14678 5020 14680
rect 5044 14678 5100 14680
rect 5124 14678 5180 14680
rect 5204 14678 5260 14680
rect 5284 14678 5340 14680
rect 4964 14626 4966 14678
rect 4966 14626 5018 14678
rect 5018 14626 5020 14678
rect 5044 14626 5082 14678
rect 5082 14626 5094 14678
rect 5094 14626 5100 14678
rect 5124 14626 5146 14678
rect 5146 14626 5158 14678
rect 5158 14626 5180 14678
rect 5204 14626 5210 14678
rect 5210 14626 5222 14678
rect 5222 14626 5260 14678
rect 5284 14626 5286 14678
rect 5286 14626 5338 14678
rect 5338 14626 5340 14678
rect 4964 14624 5020 14626
rect 5044 14624 5100 14626
rect 5124 14624 5180 14626
rect 5204 14624 5260 14626
rect 5284 14624 5340 14626
rect 4964 13346 5020 13348
rect 5044 13346 5100 13348
rect 5124 13346 5180 13348
rect 5204 13346 5260 13348
rect 5284 13346 5340 13348
rect 4964 13294 4966 13346
rect 4966 13294 5018 13346
rect 5018 13294 5020 13346
rect 5044 13294 5082 13346
rect 5082 13294 5094 13346
rect 5094 13294 5100 13346
rect 5124 13294 5146 13346
rect 5146 13294 5158 13346
rect 5158 13294 5180 13346
rect 5204 13294 5210 13346
rect 5210 13294 5222 13346
rect 5222 13294 5260 13346
rect 5284 13294 5286 13346
rect 5286 13294 5338 13346
rect 5338 13294 5340 13346
rect 4964 13292 5020 13294
rect 5044 13292 5100 13294
rect 5124 13292 5180 13294
rect 5204 13292 5260 13294
rect 5284 13292 5340 13294
rect 1556 1822 1612 1878
rect 1964 3356 2020 3358
rect 2044 3356 2100 3358
rect 2124 3356 2180 3358
rect 2204 3356 2260 3358
rect 2284 3356 2340 3358
rect 1964 3304 1966 3356
rect 1966 3304 2018 3356
rect 2018 3304 2020 3356
rect 2044 3304 2082 3356
rect 2082 3304 2094 3356
rect 2094 3304 2100 3356
rect 2124 3304 2146 3356
rect 2146 3304 2158 3356
rect 2158 3304 2180 3356
rect 2204 3304 2210 3356
rect 2210 3304 2222 3356
rect 2222 3304 2260 3356
rect 2284 3304 2286 3356
rect 2286 3304 2338 3356
rect 2338 3304 2340 3356
rect 1964 3302 2020 3304
rect 2044 3302 2100 3304
rect 2124 3302 2180 3304
rect 2204 3302 2260 3304
rect 2284 3302 2340 3304
rect 3860 5818 3916 5874
rect 4964 12014 5020 12016
rect 5044 12014 5100 12016
rect 5124 12014 5180 12016
rect 5204 12014 5260 12016
rect 5284 12014 5340 12016
rect 4964 11962 4966 12014
rect 4966 11962 5018 12014
rect 5018 11962 5020 12014
rect 5044 11962 5082 12014
rect 5082 11962 5094 12014
rect 5094 11962 5100 12014
rect 5124 11962 5146 12014
rect 5146 11962 5158 12014
rect 5158 11962 5180 12014
rect 5204 11962 5210 12014
rect 5210 11962 5222 12014
rect 5222 11962 5260 12014
rect 5284 11962 5286 12014
rect 5286 11962 5338 12014
rect 5338 11962 5340 12014
rect 4964 11960 5020 11962
rect 5044 11960 5100 11962
rect 5124 11960 5180 11962
rect 5204 11960 5260 11962
rect 5284 11960 5340 11962
rect 4964 10682 5020 10684
rect 5044 10682 5100 10684
rect 5124 10682 5180 10684
rect 5204 10682 5260 10684
rect 5284 10682 5340 10684
rect 4964 10630 4966 10682
rect 4966 10630 5018 10682
rect 5018 10630 5020 10682
rect 5044 10630 5082 10682
rect 5082 10630 5094 10682
rect 5094 10630 5100 10682
rect 5124 10630 5146 10682
rect 5146 10630 5158 10682
rect 5158 10630 5180 10682
rect 5204 10630 5210 10682
rect 5210 10630 5222 10682
rect 5222 10630 5260 10682
rect 5284 10630 5286 10682
rect 5286 10630 5338 10682
rect 5338 10630 5340 10682
rect 4964 10628 5020 10630
rect 5044 10628 5100 10630
rect 5124 10628 5180 10630
rect 5204 10628 5260 10630
rect 5284 10628 5340 10630
rect 4964 9350 5020 9352
rect 5044 9350 5100 9352
rect 5124 9350 5180 9352
rect 5204 9350 5260 9352
rect 5284 9350 5340 9352
rect 4964 9298 4966 9350
rect 4966 9298 5018 9350
rect 5018 9298 5020 9350
rect 5044 9298 5082 9350
rect 5082 9298 5094 9350
rect 5094 9298 5100 9350
rect 5124 9298 5146 9350
rect 5146 9298 5158 9350
rect 5158 9298 5180 9350
rect 5204 9298 5210 9350
rect 5210 9298 5222 9350
rect 5222 9298 5260 9350
rect 5284 9298 5286 9350
rect 5286 9298 5338 9350
rect 5338 9298 5340 9350
rect 4964 9296 5020 9298
rect 5044 9296 5100 9298
rect 5124 9296 5180 9298
rect 5204 9296 5260 9298
rect 5284 9296 5340 9298
rect 4964 8018 5020 8020
rect 5044 8018 5100 8020
rect 5124 8018 5180 8020
rect 5204 8018 5260 8020
rect 5284 8018 5340 8020
rect 4964 7966 4966 8018
rect 4966 7966 5018 8018
rect 5018 7966 5020 8018
rect 5044 7966 5082 8018
rect 5082 7966 5094 8018
rect 5094 7966 5100 8018
rect 5124 7966 5146 8018
rect 5146 7966 5158 8018
rect 5158 7966 5180 8018
rect 5204 7966 5210 8018
rect 5210 7966 5222 8018
rect 5222 7966 5260 8018
rect 5284 7966 5286 8018
rect 5286 7966 5338 8018
rect 5338 7966 5340 8018
rect 4964 7964 5020 7966
rect 5044 7964 5100 7966
rect 5124 7964 5180 7966
rect 5204 7964 5260 7966
rect 5284 7964 5340 7966
rect 4964 6686 5020 6688
rect 5044 6686 5100 6688
rect 5124 6686 5180 6688
rect 5204 6686 5260 6688
rect 5284 6686 5340 6688
rect 4964 6634 4966 6686
rect 4966 6634 5018 6686
rect 5018 6634 5020 6686
rect 5044 6634 5082 6686
rect 5082 6634 5094 6686
rect 5094 6634 5100 6686
rect 5124 6634 5146 6686
rect 5146 6634 5158 6686
rect 5158 6634 5180 6686
rect 5204 6634 5210 6686
rect 5210 6634 5222 6686
rect 5222 6634 5260 6686
rect 5284 6634 5286 6686
rect 5286 6634 5338 6686
rect 5338 6634 5340 6686
rect 4964 6632 5020 6634
rect 5044 6632 5100 6634
rect 5124 6632 5180 6634
rect 5204 6632 5260 6634
rect 5284 6632 5340 6634
rect 5108 6301 5110 6318
rect 5110 6301 5162 6318
rect 5162 6301 5164 6318
rect 5108 6262 5164 6301
rect 4964 5354 5020 5356
rect 5044 5354 5100 5356
rect 5124 5354 5180 5356
rect 5204 5354 5260 5356
rect 5284 5354 5340 5356
rect 4964 5302 4966 5354
rect 4966 5302 5018 5354
rect 5018 5302 5020 5354
rect 5044 5302 5082 5354
rect 5082 5302 5094 5354
rect 5094 5302 5100 5354
rect 5124 5302 5146 5354
rect 5146 5302 5158 5354
rect 5158 5302 5180 5354
rect 5204 5302 5210 5354
rect 5210 5302 5222 5354
rect 5222 5302 5260 5354
rect 5284 5302 5286 5354
rect 5286 5302 5338 5354
rect 5338 5302 5340 5354
rect 4964 5300 5020 5302
rect 5044 5300 5100 5302
rect 5124 5300 5180 5302
rect 5204 5300 5260 5302
rect 5284 5300 5340 5302
rect 4964 4022 5020 4024
rect 5044 4022 5100 4024
rect 5124 4022 5180 4024
rect 5204 4022 5260 4024
rect 5284 4022 5340 4024
rect 4964 3970 4966 4022
rect 4966 3970 5018 4022
rect 5018 3970 5020 4022
rect 5044 3970 5082 4022
rect 5082 3970 5094 4022
rect 5094 3970 5100 4022
rect 5124 3970 5146 4022
rect 5146 3970 5158 4022
rect 5158 3970 5180 4022
rect 5204 3970 5210 4022
rect 5210 3970 5222 4022
rect 5222 3970 5260 4022
rect 5284 3970 5286 4022
rect 5286 3970 5338 4022
rect 5338 3970 5340 4022
rect 4964 3968 5020 3970
rect 5044 3968 5100 3970
rect 5124 3968 5180 3970
rect 5204 3968 5260 3970
rect 5284 3968 5340 3970
rect 7964 24668 8020 24670
rect 8044 24668 8100 24670
rect 8124 24668 8180 24670
rect 8204 24668 8260 24670
rect 8284 24668 8340 24670
rect 7964 24616 7966 24668
rect 7966 24616 8018 24668
rect 8018 24616 8020 24668
rect 8044 24616 8082 24668
rect 8082 24616 8094 24668
rect 8094 24616 8100 24668
rect 8124 24616 8146 24668
rect 8146 24616 8158 24668
rect 8158 24616 8180 24668
rect 8204 24616 8210 24668
rect 8210 24616 8222 24668
rect 8222 24616 8260 24668
rect 8284 24616 8286 24668
rect 8286 24616 8338 24668
rect 8338 24616 8340 24668
rect 7964 24614 8020 24616
rect 8044 24614 8100 24616
rect 8124 24614 8180 24616
rect 8204 24614 8260 24616
rect 8284 24614 8340 24616
rect 7964 23336 8020 23338
rect 8044 23336 8100 23338
rect 8124 23336 8180 23338
rect 8204 23336 8260 23338
rect 8284 23336 8340 23338
rect 7964 23284 7966 23336
rect 7966 23284 8018 23336
rect 8018 23284 8020 23336
rect 8044 23284 8082 23336
rect 8082 23284 8094 23336
rect 8094 23284 8100 23336
rect 8124 23284 8146 23336
rect 8146 23284 8158 23336
rect 8158 23284 8180 23336
rect 8204 23284 8210 23336
rect 8210 23284 8222 23336
rect 8222 23284 8260 23336
rect 8284 23284 8286 23336
rect 8286 23284 8338 23336
rect 8338 23284 8340 23336
rect 7964 23282 8020 23284
rect 8044 23282 8100 23284
rect 8124 23282 8180 23284
rect 8204 23282 8260 23284
rect 8284 23282 8340 23284
rect 7964 22004 8020 22006
rect 8044 22004 8100 22006
rect 8124 22004 8180 22006
rect 8204 22004 8260 22006
rect 8284 22004 8340 22006
rect 7964 21952 7966 22004
rect 7966 21952 8018 22004
rect 8018 21952 8020 22004
rect 8044 21952 8082 22004
rect 8082 21952 8094 22004
rect 8094 21952 8100 22004
rect 8124 21952 8146 22004
rect 8146 21952 8158 22004
rect 8158 21952 8180 22004
rect 8204 21952 8210 22004
rect 8210 21952 8222 22004
rect 8222 21952 8260 22004
rect 8284 21952 8286 22004
rect 8286 21952 8338 22004
rect 8338 21952 8340 22004
rect 7964 21950 8020 21952
rect 8044 21950 8100 21952
rect 8124 21950 8180 21952
rect 8204 21950 8260 21952
rect 8284 21950 8340 21952
rect 7964 20672 8020 20674
rect 8044 20672 8100 20674
rect 8124 20672 8180 20674
rect 8204 20672 8260 20674
rect 8284 20672 8340 20674
rect 7964 20620 7966 20672
rect 7966 20620 8018 20672
rect 8018 20620 8020 20672
rect 8044 20620 8082 20672
rect 8082 20620 8094 20672
rect 8094 20620 8100 20672
rect 8124 20620 8146 20672
rect 8146 20620 8158 20672
rect 8158 20620 8180 20672
rect 8204 20620 8210 20672
rect 8210 20620 8222 20672
rect 8222 20620 8260 20672
rect 8284 20620 8286 20672
rect 8286 20620 8338 20672
rect 8338 20620 8340 20672
rect 7964 20618 8020 20620
rect 8044 20618 8100 20620
rect 8124 20618 8180 20620
rect 8204 20618 8260 20620
rect 8284 20618 8340 20620
rect 7964 19340 8020 19342
rect 8044 19340 8100 19342
rect 8124 19340 8180 19342
rect 8204 19340 8260 19342
rect 8284 19340 8340 19342
rect 7964 19288 7966 19340
rect 7966 19288 8018 19340
rect 8018 19288 8020 19340
rect 8044 19288 8082 19340
rect 8082 19288 8094 19340
rect 8094 19288 8100 19340
rect 8124 19288 8146 19340
rect 8146 19288 8158 19340
rect 8158 19288 8180 19340
rect 8204 19288 8210 19340
rect 8210 19288 8222 19340
rect 8222 19288 8260 19340
rect 8284 19288 8286 19340
rect 8286 19288 8338 19340
rect 8338 19288 8340 19340
rect 7964 19286 8020 19288
rect 8044 19286 8100 19288
rect 8124 19286 8180 19288
rect 8204 19286 8260 19288
rect 8284 19286 8340 19288
rect 7964 18008 8020 18010
rect 8044 18008 8100 18010
rect 8124 18008 8180 18010
rect 8204 18008 8260 18010
rect 8284 18008 8340 18010
rect 7964 17956 7966 18008
rect 7966 17956 8018 18008
rect 8018 17956 8020 18008
rect 8044 17956 8082 18008
rect 8082 17956 8094 18008
rect 8094 17956 8100 18008
rect 8124 17956 8146 18008
rect 8146 17956 8158 18008
rect 8158 17956 8180 18008
rect 8204 17956 8210 18008
rect 8210 17956 8222 18008
rect 8222 17956 8260 18008
rect 8284 17956 8286 18008
rect 8286 17956 8338 18008
rect 8338 17956 8340 18008
rect 7964 17954 8020 17956
rect 8044 17954 8100 17956
rect 8124 17954 8180 17956
rect 8204 17954 8260 17956
rect 8284 17954 8340 17956
rect 7964 16676 8020 16678
rect 8044 16676 8100 16678
rect 8124 16676 8180 16678
rect 8204 16676 8260 16678
rect 8284 16676 8340 16678
rect 7964 16624 7966 16676
rect 7966 16624 8018 16676
rect 8018 16624 8020 16676
rect 8044 16624 8082 16676
rect 8082 16624 8094 16676
rect 8094 16624 8100 16676
rect 8124 16624 8146 16676
rect 8146 16624 8158 16676
rect 8158 16624 8180 16676
rect 8204 16624 8210 16676
rect 8210 16624 8222 16676
rect 8222 16624 8260 16676
rect 8284 16624 8286 16676
rect 8286 16624 8338 16676
rect 8338 16624 8340 16676
rect 7964 16622 8020 16624
rect 8044 16622 8100 16624
rect 8124 16622 8180 16624
rect 8204 16622 8260 16624
rect 8284 16622 8340 16624
rect 7964 15344 8020 15346
rect 8044 15344 8100 15346
rect 8124 15344 8180 15346
rect 8204 15344 8260 15346
rect 8284 15344 8340 15346
rect 7964 15292 7966 15344
rect 7966 15292 8018 15344
rect 8018 15292 8020 15344
rect 8044 15292 8082 15344
rect 8082 15292 8094 15344
rect 8094 15292 8100 15344
rect 8124 15292 8146 15344
rect 8146 15292 8158 15344
rect 8158 15292 8180 15344
rect 8204 15292 8210 15344
rect 8210 15292 8222 15344
rect 8222 15292 8260 15344
rect 8284 15292 8286 15344
rect 8286 15292 8338 15344
rect 8338 15292 8340 15344
rect 7964 15290 8020 15292
rect 8044 15290 8100 15292
rect 8124 15290 8180 15292
rect 8204 15290 8260 15292
rect 8284 15290 8340 15292
rect 7964 14012 8020 14014
rect 8044 14012 8100 14014
rect 8124 14012 8180 14014
rect 8204 14012 8260 14014
rect 8284 14012 8340 14014
rect 7964 13960 7966 14012
rect 7966 13960 8018 14012
rect 8018 13960 8020 14012
rect 8044 13960 8082 14012
rect 8082 13960 8094 14012
rect 8094 13960 8100 14012
rect 8124 13960 8146 14012
rect 8146 13960 8158 14012
rect 8158 13960 8180 14012
rect 8204 13960 8210 14012
rect 8210 13960 8222 14012
rect 8222 13960 8260 14012
rect 8284 13960 8286 14012
rect 8286 13960 8338 14012
rect 8338 13960 8340 14012
rect 7964 13958 8020 13960
rect 8044 13958 8100 13960
rect 8124 13958 8180 13960
rect 8204 13958 8260 13960
rect 8284 13958 8340 13960
rect 7964 12680 8020 12682
rect 8044 12680 8100 12682
rect 8124 12680 8180 12682
rect 8204 12680 8260 12682
rect 8284 12680 8340 12682
rect 7964 12628 7966 12680
rect 7966 12628 8018 12680
rect 8018 12628 8020 12680
rect 8044 12628 8082 12680
rect 8082 12628 8094 12680
rect 8094 12628 8100 12680
rect 8124 12628 8146 12680
rect 8146 12628 8158 12680
rect 8158 12628 8180 12680
rect 8204 12628 8210 12680
rect 8210 12628 8222 12680
rect 8222 12628 8260 12680
rect 8284 12628 8286 12680
rect 8286 12628 8338 12680
rect 8338 12628 8340 12680
rect 7964 12626 8020 12628
rect 8044 12626 8100 12628
rect 8124 12626 8180 12628
rect 8204 12626 8260 12628
rect 8284 12626 8340 12628
rect 7964 11348 8020 11350
rect 8044 11348 8100 11350
rect 8124 11348 8180 11350
rect 8204 11348 8260 11350
rect 8284 11348 8340 11350
rect 7964 11296 7966 11348
rect 7966 11296 8018 11348
rect 8018 11296 8020 11348
rect 8044 11296 8082 11348
rect 8082 11296 8094 11348
rect 8094 11296 8100 11348
rect 8124 11296 8146 11348
rect 8146 11296 8158 11348
rect 8158 11296 8180 11348
rect 8204 11296 8210 11348
rect 8210 11296 8222 11348
rect 8222 11296 8260 11348
rect 8284 11296 8286 11348
rect 8286 11296 8338 11348
rect 8338 11296 8340 11348
rect 7964 11294 8020 11296
rect 8044 11294 8100 11296
rect 8124 11294 8180 11296
rect 8204 11294 8260 11296
rect 8284 11294 8340 11296
rect 10100 22542 10156 22598
rect 7964 10016 8020 10018
rect 8044 10016 8100 10018
rect 8124 10016 8180 10018
rect 8204 10016 8260 10018
rect 8284 10016 8340 10018
rect 7964 9964 7966 10016
rect 7966 9964 8018 10016
rect 8018 9964 8020 10016
rect 8044 9964 8082 10016
rect 8082 9964 8094 10016
rect 8094 9964 8100 10016
rect 8124 9964 8146 10016
rect 8146 9964 8158 10016
rect 8158 9964 8180 10016
rect 8204 9964 8210 10016
rect 8210 9964 8222 10016
rect 8222 9964 8260 10016
rect 8284 9964 8286 10016
rect 8286 9964 8338 10016
rect 8338 9964 8340 10016
rect 7964 9962 8020 9964
rect 8044 9962 8100 9964
rect 8124 9962 8180 9964
rect 8204 9962 8260 9964
rect 8284 9962 8340 9964
rect 7964 8684 8020 8686
rect 8044 8684 8100 8686
rect 8124 8684 8180 8686
rect 8204 8684 8260 8686
rect 8284 8684 8340 8686
rect 7964 8632 7966 8684
rect 7966 8632 8018 8684
rect 8018 8632 8020 8684
rect 8044 8632 8082 8684
rect 8082 8632 8094 8684
rect 8094 8632 8100 8684
rect 8124 8632 8146 8684
rect 8146 8632 8158 8684
rect 8158 8632 8180 8684
rect 8204 8632 8210 8684
rect 8210 8632 8222 8684
rect 8222 8632 8260 8684
rect 8284 8632 8286 8684
rect 8286 8632 8338 8684
rect 8338 8632 8340 8684
rect 7964 8630 8020 8632
rect 8044 8630 8100 8632
rect 8124 8630 8180 8632
rect 8204 8630 8260 8632
rect 8284 8630 8340 8632
rect 7964 7352 8020 7354
rect 8044 7352 8100 7354
rect 8124 7352 8180 7354
rect 8204 7352 8260 7354
rect 8284 7352 8340 7354
rect 7964 7300 7966 7352
rect 7966 7300 8018 7352
rect 8018 7300 8020 7352
rect 8044 7300 8082 7352
rect 8082 7300 8094 7352
rect 8094 7300 8100 7352
rect 8124 7300 8146 7352
rect 8146 7300 8158 7352
rect 8158 7300 8180 7352
rect 8204 7300 8210 7352
rect 8210 7300 8222 7352
rect 8222 7300 8260 7352
rect 8284 7300 8286 7352
rect 8286 7300 8338 7352
rect 8338 7300 8340 7352
rect 7964 7298 8020 7300
rect 8044 7298 8100 7300
rect 8124 7298 8180 7300
rect 8204 7298 8260 7300
rect 8284 7298 8340 7300
rect 7964 6020 8020 6022
rect 8044 6020 8100 6022
rect 8124 6020 8180 6022
rect 8204 6020 8260 6022
rect 8284 6020 8340 6022
rect 7964 5968 7966 6020
rect 7966 5968 8018 6020
rect 8018 5968 8020 6020
rect 8044 5968 8082 6020
rect 8082 5968 8094 6020
rect 8094 5968 8100 6020
rect 8124 5968 8146 6020
rect 8146 5968 8158 6020
rect 8158 5968 8180 6020
rect 8204 5968 8210 6020
rect 8210 5968 8222 6020
rect 8222 5968 8260 6020
rect 8284 5968 8286 6020
rect 8286 5968 8338 6020
rect 8338 5968 8340 6020
rect 7964 5966 8020 5968
rect 8044 5966 8100 5968
rect 8124 5966 8180 5968
rect 8204 5966 8260 5968
rect 8284 5966 8340 5968
rect 7964 4688 8020 4690
rect 8044 4688 8100 4690
rect 8124 4688 8180 4690
rect 8204 4688 8260 4690
rect 8284 4688 8340 4690
rect 7964 4636 7966 4688
rect 7966 4636 8018 4688
rect 8018 4636 8020 4688
rect 8044 4636 8082 4688
rect 8082 4636 8094 4688
rect 8094 4636 8100 4688
rect 8124 4636 8146 4688
rect 8146 4636 8158 4688
rect 8158 4636 8180 4688
rect 8204 4636 8210 4688
rect 8210 4636 8222 4688
rect 8222 4636 8260 4688
rect 8284 4636 8286 4688
rect 8286 4636 8338 4688
rect 8338 4636 8340 4688
rect 7964 4634 8020 4636
rect 8044 4634 8100 4636
rect 8124 4634 8180 4636
rect 8204 4634 8260 4636
rect 8284 4634 8340 4636
rect 7964 3356 8020 3358
rect 8044 3356 8100 3358
rect 8124 3356 8180 3358
rect 8204 3356 8260 3358
rect 8284 3356 8340 3358
rect 7964 3304 7966 3356
rect 7966 3304 8018 3356
rect 8018 3304 8020 3356
rect 8044 3304 8082 3356
rect 8082 3304 8094 3356
rect 8094 3304 8100 3356
rect 8124 3304 8146 3356
rect 8146 3304 8158 3356
rect 8158 3304 8180 3356
rect 8204 3304 8210 3356
rect 8210 3304 8222 3356
rect 8222 3304 8260 3356
rect 8284 3304 8286 3356
rect 8286 3304 8338 3356
rect 8338 3304 8340 3356
rect 7964 3302 8020 3304
rect 8044 3302 8100 3304
rect 8124 3302 8180 3304
rect 8204 3302 8260 3304
rect 8284 3302 8340 3304
rect 10100 20191 10156 20230
rect 10100 20174 10102 20191
rect 10102 20174 10154 20191
rect 10154 20174 10156 20191
rect 10100 17806 10156 17862
rect 10100 15455 10156 15494
rect 10100 15438 10102 15455
rect 10102 15438 10154 15455
rect 10154 15438 10156 15455
rect 10100 13070 10156 13126
rect 10100 10741 10102 10758
rect 10102 10741 10154 10758
rect 10154 10741 10156 10758
rect 10100 10702 10156 10741
rect 10100 8351 10156 8390
rect 10100 8334 10102 8351
rect 10102 8334 10154 8351
rect 10154 8334 10156 8351
rect 10100 5966 10156 6022
rect 10100 3615 10156 3654
rect 10100 3598 10102 3615
rect 10102 3598 10154 3615
rect 10154 3598 10156 3615
rect 4964 2690 5020 2692
rect 5044 2690 5100 2692
rect 5124 2690 5180 2692
rect 5204 2690 5260 2692
rect 5284 2690 5340 2692
rect 4964 2638 4966 2690
rect 4966 2638 5018 2690
rect 5018 2638 5020 2690
rect 5044 2638 5082 2690
rect 5082 2638 5094 2690
rect 5094 2638 5100 2690
rect 5124 2638 5146 2690
rect 5146 2638 5158 2690
rect 5158 2638 5180 2690
rect 5204 2638 5210 2690
rect 5210 2638 5222 2690
rect 5222 2638 5260 2690
rect 5284 2638 5286 2690
rect 5286 2638 5338 2690
rect 5338 2638 5340 2690
rect 4964 2636 5020 2638
rect 5044 2636 5100 2638
rect 5124 2636 5180 2638
rect 5204 2636 5260 2638
rect 5284 2636 5340 2638
rect 9716 1230 9772 1286
<< metal3 >>
rect 9327 27336 9393 27339
rect 10922 27336 11722 27366
rect 9327 27334 11722 27336
rect 9327 27278 9332 27334
rect 9388 27278 11722 27334
rect 9327 27276 11722 27278
rect 9327 27273 9393 27276
rect 10922 27246 11722 27276
rect 0 26744 800 26774
rect 1455 26744 1521 26747
rect 0 26742 1521 26744
rect 0 26686 1460 26742
rect 1516 26686 1521 26742
rect 0 26684 1521 26686
rect 0 26654 800 26684
rect 1455 26681 1521 26684
rect 1954 26006 2350 26007
rect 1954 25942 1960 26006
rect 2024 25942 2040 26006
rect 2104 25942 2120 26006
rect 2184 25942 2200 26006
rect 2264 25942 2280 26006
rect 2344 25942 2350 26006
rect 1954 25941 2350 25942
rect 7954 26006 8350 26007
rect 7954 25942 7960 26006
rect 8024 25942 8040 26006
rect 8104 25942 8120 26006
rect 8184 25942 8200 26006
rect 8264 25942 8280 26006
rect 8344 25942 8350 26006
rect 7954 25941 8350 25942
rect 4954 25340 5350 25341
rect 4954 25276 4960 25340
rect 5024 25276 5040 25340
rect 5104 25276 5120 25340
rect 5184 25276 5200 25340
rect 5264 25276 5280 25340
rect 5344 25276 5350 25340
rect 4954 25275 5350 25276
rect 1954 24674 2350 24675
rect 1954 24610 1960 24674
rect 2024 24610 2040 24674
rect 2104 24610 2120 24674
rect 2184 24610 2200 24674
rect 2264 24610 2280 24674
rect 2344 24610 2350 24674
rect 1954 24609 2350 24610
rect 7954 24674 8350 24675
rect 7954 24610 7960 24674
rect 8024 24610 8040 24674
rect 8104 24610 8120 24674
rect 8184 24610 8200 24674
rect 8264 24610 8280 24674
rect 8344 24610 8350 24674
rect 7954 24609 8350 24610
rect 4954 24008 5350 24009
rect 4954 23944 4960 24008
rect 5024 23944 5040 24008
rect 5104 23944 5120 24008
rect 5184 23944 5200 24008
rect 5264 23944 5280 24008
rect 5344 23944 5350 24008
rect 4954 23943 5350 23944
rect 1954 23342 2350 23343
rect 1954 23278 1960 23342
rect 2024 23278 2040 23342
rect 2104 23278 2120 23342
rect 2184 23278 2200 23342
rect 2264 23278 2280 23342
rect 2344 23278 2350 23342
rect 1954 23277 2350 23278
rect 7954 23342 8350 23343
rect 7954 23278 7960 23342
rect 8024 23278 8040 23342
rect 8104 23278 8120 23342
rect 8184 23278 8200 23342
rect 8264 23278 8280 23342
rect 8344 23278 8350 23342
rect 7954 23277 8350 23278
rect 4954 22676 5350 22677
rect 0 22600 800 22630
rect 4954 22612 4960 22676
rect 5024 22612 5040 22676
rect 5104 22612 5120 22676
rect 5184 22612 5200 22676
rect 5264 22612 5280 22676
rect 5344 22612 5350 22676
rect 4954 22611 5350 22612
rect 1263 22600 1329 22603
rect 0 22598 1329 22600
rect 0 22542 1268 22598
rect 1324 22542 1329 22598
rect 0 22540 1329 22542
rect 0 22510 800 22540
rect 1263 22537 1329 22540
rect 10095 22600 10161 22603
rect 10922 22600 11722 22630
rect 10095 22598 11722 22600
rect 10095 22542 10100 22598
rect 10156 22542 11722 22598
rect 10095 22540 11722 22542
rect 10095 22537 10161 22540
rect 10922 22510 11722 22540
rect 1954 22010 2350 22011
rect 1954 21946 1960 22010
rect 2024 21946 2040 22010
rect 2104 21946 2120 22010
rect 2184 21946 2200 22010
rect 2264 21946 2280 22010
rect 2344 21946 2350 22010
rect 1954 21945 2350 21946
rect 7954 22010 8350 22011
rect 7954 21946 7960 22010
rect 8024 21946 8040 22010
rect 8104 21946 8120 22010
rect 8184 21946 8200 22010
rect 8264 21946 8280 22010
rect 8344 21946 8350 22010
rect 7954 21945 8350 21946
rect 4954 21344 5350 21345
rect 4954 21280 4960 21344
rect 5024 21280 5040 21344
rect 5104 21280 5120 21344
rect 5184 21280 5200 21344
rect 5264 21280 5280 21344
rect 5344 21280 5350 21344
rect 4954 21279 5350 21280
rect 1954 20678 2350 20679
rect 1954 20614 1960 20678
rect 2024 20614 2040 20678
rect 2104 20614 2120 20678
rect 2184 20614 2200 20678
rect 2264 20614 2280 20678
rect 2344 20614 2350 20678
rect 1954 20613 2350 20614
rect 7954 20678 8350 20679
rect 7954 20614 7960 20678
rect 8024 20614 8040 20678
rect 8104 20614 8120 20678
rect 8184 20614 8200 20678
rect 8264 20614 8280 20678
rect 8344 20614 8350 20678
rect 7954 20613 8350 20614
rect 10095 20232 10161 20235
rect 10922 20232 11722 20262
rect 10095 20230 11722 20232
rect 10095 20174 10100 20230
rect 10156 20174 11722 20230
rect 10095 20172 11722 20174
rect 10095 20169 10161 20172
rect 10922 20142 11722 20172
rect 4954 20012 5350 20013
rect 4954 19948 4960 20012
rect 5024 19948 5040 20012
rect 5104 19948 5120 20012
rect 5184 19948 5200 20012
rect 5264 19948 5280 20012
rect 5344 19948 5350 20012
rect 4954 19947 5350 19948
rect 1954 19346 2350 19347
rect 1954 19282 1960 19346
rect 2024 19282 2040 19346
rect 2104 19282 2120 19346
rect 2184 19282 2200 19346
rect 2264 19282 2280 19346
rect 2344 19282 2350 19346
rect 1954 19281 2350 19282
rect 7954 19346 8350 19347
rect 7954 19282 7960 19346
rect 8024 19282 8040 19346
rect 8104 19282 8120 19346
rect 8184 19282 8200 19346
rect 8264 19282 8280 19346
rect 8344 19282 8350 19346
rect 7954 19281 8350 19282
rect 4954 18680 5350 18681
rect 4954 18616 4960 18680
rect 5024 18616 5040 18680
rect 5104 18616 5120 18680
rect 5184 18616 5200 18680
rect 5264 18616 5280 18680
rect 5344 18616 5350 18680
rect 4954 18615 5350 18616
rect 0 18456 800 18486
rect 1647 18456 1713 18459
rect 0 18454 1713 18456
rect 0 18398 1652 18454
rect 1708 18398 1713 18454
rect 0 18396 1713 18398
rect 0 18366 800 18396
rect 1647 18393 1713 18396
rect 1954 18014 2350 18015
rect 1954 17950 1960 18014
rect 2024 17950 2040 18014
rect 2104 17950 2120 18014
rect 2184 17950 2200 18014
rect 2264 17950 2280 18014
rect 2344 17950 2350 18014
rect 1954 17949 2350 17950
rect 7954 18014 8350 18015
rect 7954 17950 7960 18014
rect 8024 17950 8040 18014
rect 8104 17950 8120 18014
rect 8184 17950 8200 18014
rect 8264 17950 8280 18014
rect 8344 17950 8350 18014
rect 7954 17949 8350 17950
rect 10095 17864 10161 17867
rect 10922 17864 11722 17894
rect 10095 17862 11722 17864
rect 10095 17806 10100 17862
rect 10156 17806 11722 17862
rect 10095 17804 11722 17806
rect 10095 17801 10161 17804
rect 10922 17774 11722 17804
rect 4954 17348 5350 17349
rect 4954 17284 4960 17348
rect 5024 17284 5040 17348
rect 5104 17284 5120 17348
rect 5184 17284 5200 17348
rect 5264 17284 5280 17348
rect 5344 17284 5350 17348
rect 4954 17283 5350 17284
rect 1954 16682 2350 16683
rect 1954 16618 1960 16682
rect 2024 16618 2040 16682
rect 2104 16618 2120 16682
rect 2184 16618 2200 16682
rect 2264 16618 2280 16682
rect 2344 16618 2350 16682
rect 1954 16617 2350 16618
rect 7954 16682 8350 16683
rect 7954 16618 7960 16682
rect 8024 16618 8040 16682
rect 8104 16618 8120 16682
rect 8184 16618 8200 16682
rect 8264 16618 8280 16682
rect 8344 16618 8350 16682
rect 7954 16617 8350 16618
rect 4954 16016 5350 16017
rect 4954 15952 4960 16016
rect 5024 15952 5040 16016
rect 5104 15952 5120 16016
rect 5184 15952 5200 16016
rect 5264 15952 5280 16016
rect 5344 15952 5350 16016
rect 4954 15951 5350 15952
rect 10095 15496 10161 15499
rect 10922 15496 11722 15526
rect 10095 15494 11722 15496
rect 10095 15438 10100 15494
rect 10156 15438 11722 15494
rect 10095 15436 11722 15438
rect 10095 15433 10161 15436
rect 10922 15406 11722 15436
rect 1954 15350 2350 15351
rect 1954 15286 1960 15350
rect 2024 15286 2040 15350
rect 2104 15286 2120 15350
rect 2184 15286 2200 15350
rect 2264 15286 2280 15350
rect 2344 15286 2350 15350
rect 1954 15285 2350 15286
rect 7954 15350 8350 15351
rect 7954 15286 7960 15350
rect 8024 15286 8040 15350
rect 8104 15286 8120 15350
rect 8184 15286 8200 15350
rect 8264 15286 8280 15350
rect 8344 15286 8350 15350
rect 7954 15285 8350 15286
rect 4954 14684 5350 14685
rect 4954 14620 4960 14684
rect 5024 14620 5040 14684
rect 5104 14620 5120 14684
rect 5184 14620 5200 14684
rect 5264 14620 5280 14684
rect 5344 14620 5350 14684
rect 4954 14619 5350 14620
rect 0 14312 800 14342
rect 879 14312 945 14315
rect 0 14310 945 14312
rect 0 14254 884 14310
rect 940 14254 945 14310
rect 0 14252 945 14254
rect 0 14222 800 14252
rect 879 14249 945 14252
rect 1954 14018 2350 14019
rect 1954 13954 1960 14018
rect 2024 13954 2040 14018
rect 2104 13954 2120 14018
rect 2184 13954 2200 14018
rect 2264 13954 2280 14018
rect 2344 13954 2350 14018
rect 1954 13953 2350 13954
rect 7954 14018 8350 14019
rect 7954 13954 7960 14018
rect 8024 13954 8040 14018
rect 8104 13954 8120 14018
rect 8184 13954 8200 14018
rect 8264 13954 8280 14018
rect 8344 13954 8350 14018
rect 7954 13953 8350 13954
rect 4954 13352 5350 13353
rect 4954 13288 4960 13352
rect 5024 13288 5040 13352
rect 5104 13288 5120 13352
rect 5184 13288 5200 13352
rect 5264 13288 5280 13352
rect 5344 13288 5350 13352
rect 4954 13287 5350 13288
rect 10095 13128 10161 13131
rect 10922 13128 11722 13158
rect 10095 13126 11722 13128
rect 10095 13070 10100 13126
rect 10156 13070 11722 13126
rect 10095 13068 11722 13070
rect 10095 13065 10161 13068
rect 10922 13038 11722 13068
rect 1954 12686 2350 12687
rect 1954 12622 1960 12686
rect 2024 12622 2040 12686
rect 2104 12622 2120 12686
rect 2184 12622 2200 12686
rect 2264 12622 2280 12686
rect 2344 12622 2350 12686
rect 1954 12621 2350 12622
rect 7954 12686 8350 12687
rect 7954 12622 7960 12686
rect 8024 12622 8040 12686
rect 8104 12622 8120 12686
rect 8184 12622 8200 12686
rect 8264 12622 8280 12686
rect 8344 12622 8350 12686
rect 7954 12621 8350 12622
rect 4954 12020 5350 12021
rect 4954 11956 4960 12020
rect 5024 11956 5040 12020
rect 5104 11956 5120 12020
rect 5184 11956 5200 12020
rect 5264 11956 5280 12020
rect 5344 11956 5350 12020
rect 4954 11955 5350 11956
rect 1954 11354 2350 11355
rect 1954 11290 1960 11354
rect 2024 11290 2040 11354
rect 2104 11290 2120 11354
rect 2184 11290 2200 11354
rect 2264 11290 2280 11354
rect 2344 11290 2350 11354
rect 1954 11289 2350 11290
rect 7954 11354 8350 11355
rect 7954 11290 7960 11354
rect 8024 11290 8040 11354
rect 8104 11290 8120 11354
rect 8184 11290 8200 11354
rect 8264 11290 8280 11354
rect 8344 11290 8350 11354
rect 7954 11289 8350 11290
rect 10095 10760 10161 10763
rect 10922 10760 11722 10790
rect 10095 10758 11722 10760
rect 10095 10702 10100 10758
rect 10156 10702 11722 10758
rect 10095 10700 11722 10702
rect 10095 10697 10161 10700
rect 4954 10688 5350 10689
rect 4954 10624 4960 10688
rect 5024 10624 5040 10688
rect 5104 10624 5120 10688
rect 5184 10624 5200 10688
rect 5264 10624 5280 10688
rect 5344 10624 5350 10688
rect 10922 10670 11722 10700
rect 4954 10623 5350 10624
rect 0 10168 800 10198
rect 879 10168 945 10171
rect 0 10166 945 10168
rect 0 10110 884 10166
rect 940 10110 945 10166
rect 0 10108 945 10110
rect 0 10078 800 10108
rect 879 10105 945 10108
rect 1954 10022 2350 10023
rect 1954 9958 1960 10022
rect 2024 9958 2040 10022
rect 2104 9958 2120 10022
rect 2184 9958 2200 10022
rect 2264 9958 2280 10022
rect 2344 9958 2350 10022
rect 1954 9957 2350 9958
rect 7954 10022 8350 10023
rect 7954 9958 7960 10022
rect 8024 9958 8040 10022
rect 8104 9958 8120 10022
rect 8184 9958 8200 10022
rect 8264 9958 8280 10022
rect 8344 9958 8350 10022
rect 7954 9957 8350 9958
rect 4954 9356 5350 9357
rect 4954 9292 4960 9356
rect 5024 9292 5040 9356
rect 5104 9292 5120 9356
rect 5184 9292 5200 9356
rect 5264 9292 5280 9356
rect 5344 9292 5350 9356
rect 4954 9291 5350 9292
rect 1954 8690 2350 8691
rect 1954 8626 1960 8690
rect 2024 8626 2040 8690
rect 2104 8626 2120 8690
rect 2184 8626 2200 8690
rect 2264 8626 2280 8690
rect 2344 8626 2350 8690
rect 1954 8625 2350 8626
rect 7954 8690 8350 8691
rect 7954 8626 7960 8690
rect 8024 8626 8040 8690
rect 8104 8626 8120 8690
rect 8184 8626 8200 8690
rect 8264 8626 8280 8690
rect 8344 8626 8350 8690
rect 7954 8625 8350 8626
rect 10095 8392 10161 8395
rect 10922 8392 11722 8422
rect 10095 8390 11722 8392
rect 10095 8334 10100 8390
rect 10156 8334 11722 8390
rect 10095 8332 11722 8334
rect 10095 8329 10161 8332
rect 10922 8302 11722 8332
rect 4954 8024 5350 8025
rect 4954 7960 4960 8024
rect 5024 7960 5040 8024
rect 5104 7960 5120 8024
rect 5184 7960 5200 8024
rect 5264 7960 5280 8024
rect 5344 7960 5350 8024
rect 4954 7959 5350 7960
rect 1954 7358 2350 7359
rect 1954 7294 1960 7358
rect 2024 7294 2040 7358
rect 2104 7294 2120 7358
rect 2184 7294 2200 7358
rect 2264 7294 2280 7358
rect 2344 7294 2350 7358
rect 1954 7293 2350 7294
rect 7954 7358 8350 7359
rect 7954 7294 7960 7358
rect 8024 7294 8040 7358
rect 8104 7294 8120 7358
rect 8184 7294 8200 7358
rect 8264 7294 8280 7358
rect 8344 7294 8350 7358
rect 7954 7293 8350 7294
rect 4954 6692 5350 6693
rect 4954 6628 4960 6692
rect 5024 6628 5040 6692
rect 5104 6628 5120 6692
rect 5184 6628 5200 6692
rect 5264 6628 5280 6692
rect 5344 6628 5350 6692
rect 4954 6627 5350 6628
rect 1743 6320 1809 6323
rect 5103 6320 5169 6323
rect 1743 6318 5169 6320
rect 1743 6262 1748 6318
rect 1804 6262 5108 6318
rect 5164 6262 5169 6318
rect 1743 6260 5169 6262
rect 1743 6257 1809 6260
rect 5103 6257 5169 6260
rect 0 6024 800 6054
rect 1954 6026 2350 6027
rect 0 5964 1470 6024
rect 0 5934 800 5964
rect 1410 5876 1470 5964
rect 1954 5962 1960 6026
rect 2024 5962 2040 6026
rect 2104 5962 2120 6026
rect 2184 5962 2200 6026
rect 2264 5962 2280 6026
rect 2344 5962 2350 6026
rect 1954 5961 2350 5962
rect 7954 6026 8350 6027
rect 7954 5962 7960 6026
rect 8024 5962 8040 6026
rect 8104 5962 8120 6026
rect 8184 5962 8200 6026
rect 8264 5962 8280 6026
rect 8344 5962 8350 6026
rect 7954 5961 8350 5962
rect 10095 6024 10161 6027
rect 10922 6024 11722 6054
rect 10095 6022 11722 6024
rect 10095 5966 10100 6022
rect 10156 5966 11722 6022
rect 10095 5964 11722 5966
rect 10095 5961 10161 5964
rect 10922 5934 11722 5964
rect 3855 5876 3921 5879
rect 1410 5874 3921 5876
rect 1410 5818 3860 5874
rect 3916 5818 3921 5874
rect 1410 5816 3921 5818
rect 3855 5813 3921 5816
rect 4954 5360 5350 5361
rect 4954 5296 4960 5360
rect 5024 5296 5040 5360
rect 5104 5296 5120 5360
rect 5184 5296 5200 5360
rect 5264 5296 5280 5360
rect 5344 5296 5350 5360
rect 4954 5295 5350 5296
rect 1954 4694 2350 4695
rect 1954 4630 1960 4694
rect 2024 4630 2040 4694
rect 2104 4630 2120 4694
rect 2184 4630 2200 4694
rect 2264 4630 2280 4694
rect 2344 4630 2350 4694
rect 1954 4629 2350 4630
rect 7954 4694 8350 4695
rect 7954 4630 7960 4694
rect 8024 4630 8040 4694
rect 8104 4630 8120 4694
rect 8184 4630 8200 4694
rect 8264 4630 8280 4694
rect 8344 4630 8350 4694
rect 7954 4629 8350 4630
rect 4954 4028 5350 4029
rect 4954 3964 4960 4028
rect 5024 3964 5040 4028
rect 5104 3964 5120 4028
rect 5184 3964 5200 4028
rect 5264 3964 5280 4028
rect 5344 3964 5350 4028
rect 4954 3963 5350 3964
rect 10095 3656 10161 3659
rect 10922 3656 11722 3686
rect 10095 3654 11722 3656
rect 10095 3598 10100 3654
rect 10156 3598 11722 3654
rect 10095 3596 11722 3598
rect 10095 3593 10161 3596
rect 10922 3566 11722 3596
rect 1954 3362 2350 3363
rect 1954 3298 1960 3362
rect 2024 3298 2040 3362
rect 2104 3298 2120 3362
rect 2184 3298 2200 3362
rect 2264 3298 2280 3362
rect 2344 3298 2350 3362
rect 1954 3297 2350 3298
rect 7954 3362 8350 3363
rect 7954 3298 7960 3362
rect 8024 3298 8040 3362
rect 8104 3298 8120 3362
rect 8184 3298 8200 3362
rect 8264 3298 8280 3362
rect 8344 3298 8350 3362
rect 7954 3297 8350 3298
rect 4954 2696 5350 2697
rect 4954 2632 4960 2696
rect 5024 2632 5040 2696
rect 5104 2632 5120 2696
rect 5184 2632 5200 2696
rect 5264 2632 5280 2696
rect 5344 2632 5350 2696
rect 4954 2631 5350 2632
rect 0 1880 800 1910
rect 1551 1880 1617 1883
rect 0 1878 1617 1880
rect 0 1822 1556 1878
rect 1612 1822 1617 1878
rect 0 1820 1617 1822
rect 0 1790 800 1820
rect 1551 1817 1617 1820
rect 9711 1288 9777 1291
rect 10922 1288 11722 1318
rect 9711 1286 11722 1288
rect 9711 1230 9716 1286
rect 9772 1230 11722 1286
rect 9711 1228 11722 1230
rect 9711 1225 9777 1228
rect 10922 1198 11722 1228
<< via3 >>
rect 1960 26002 2024 26006
rect 1960 25946 1964 26002
rect 1964 25946 2020 26002
rect 2020 25946 2024 26002
rect 1960 25942 2024 25946
rect 2040 26002 2104 26006
rect 2040 25946 2044 26002
rect 2044 25946 2100 26002
rect 2100 25946 2104 26002
rect 2040 25942 2104 25946
rect 2120 26002 2184 26006
rect 2120 25946 2124 26002
rect 2124 25946 2180 26002
rect 2180 25946 2184 26002
rect 2120 25942 2184 25946
rect 2200 26002 2264 26006
rect 2200 25946 2204 26002
rect 2204 25946 2260 26002
rect 2260 25946 2264 26002
rect 2200 25942 2264 25946
rect 2280 26002 2344 26006
rect 2280 25946 2284 26002
rect 2284 25946 2340 26002
rect 2340 25946 2344 26002
rect 2280 25942 2344 25946
rect 7960 26002 8024 26006
rect 7960 25946 7964 26002
rect 7964 25946 8020 26002
rect 8020 25946 8024 26002
rect 7960 25942 8024 25946
rect 8040 26002 8104 26006
rect 8040 25946 8044 26002
rect 8044 25946 8100 26002
rect 8100 25946 8104 26002
rect 8040 25942 8104 25946
rect 8120 26002 8184 26006
rect 8120 25946 8124 26002
rect 8124 25946 8180 26002
rect 8180 25946 8184 26002
rect 8120 25942 8184 25946
rect 8200 26002 8264 26006
rect 8200 25946 8204 26002
rect 8204 25946 8260 26002
rect 8260 25946 8264 26002
rect 8200 25942 8264 25946
rect 8280 26002 8344 26006
rect 8280 25946 8284 26002
rect 8284 25946 8340 26002
rect 8340 25946 8344 26002
rect 8280 25942 8344 25946
rect 4960 25336 5024 25340
rect 4960 25280 4964 25336
rect 4964 25280 5020 25336
rect 5020 25280 5024 25336
rect 4960 25276 5024 25280
rect 5040 25336 5104 25340
rect 5040 25280 5044 25336
rect 5044 25280 5100 25336
rect 5100 25280 5104 25336
rect 5040 25276 5104 25280
rect 5120 25336 5184 25340
rect 5120 25280 5124 25336
rect 5124 25280 5180 25336
rect 5180 25280 5184 25336
rect 5120 25276 5184 25280
rect 5200 25336 5264 25340
rect 5200 25280 5204 25336
rect 5204 25280 5260 25336
rect 5260 25280 5264 25336
rect 5200 25276 5264 25280
rect 5280 25336 5344 25340
rect 5280 25280 5284 25336
rect 5284 25280 5340 25336
rect 5340 25280 5344 25336
rect 5280 25276 5344 25280
rect 1960 24670 2024 24674
rect 1960 24614 1964 24670
rect 1964 24614 2020 24670
rect 2020 24614 2024 24670
rect 1960 24610 2024 24614
rect 2040 24670 2104 24674
rect 2040 24614 2044 24670
rect 2044 24614 2100 24670
rect 2100 24614 2104 24670
rect 2040 24610 2104 24614
rect 2120 24670 2184 24674
rect 2120 24614 2124 24670
rect 2124 24614 2180 24670
rect 2180 24614 2184 24670
rect 2120 24610 2184 24614
rect 2200 24670 2264 24674
rect 2200 24614 2204 24670
rect 2204 24614 2260 24670
rect 2260 24614 2264 24670
rect 2200 24610 2264 24614
rect 2280 24670 2344 24674
rect 2280 24614 2284 24670
rect 2284 24614 2340 24670
rect 2340 24614 2344 24670
rect 2280 24610 2344 24614
rect 7960 24670 8024 24674
rect 7960 24614 7964 24670
rect 7964 24614 8020 24670
rect 8020 24614 8024 24670
rect 7960 24610 8024 24614
rect 8040 24670 8104 24674
rect 8040 24614 8044 24670
rect 8044 24614 8100 24670
rect 8100 24614 8104 24670
rect 8040 24610 8104 24614
rect 8120 24670 8184 24674
rect 8120 24614 8124 24670
rect 8124 24614 8180 24670
rect 8180 24614 8184 24670
rect 8120 24610 8184 24614
rect 8200 24670 8264 24674
rect 8200 24614 8204 24670
rect 8204 24614 8260 24670
rect 8260 24614 8264 24670
rect 8200 24610 8264 24614
rect 8280 24670 8344 24674
rect 8280 24614 8284 24670
rect 8284 24614 8340 24670
rect 8340 24614 8344 24670
rect 8280 24610 8344 24614
rect 4960 24004 5024 24008
rect 4960 23948 4964 24004
rect 4964 23948 5020 24004
rect 5020 23948 5024 24004
rect 4960 23944 5024 23948
rect 5040 24004 5104 24008
rect 5040 23948 5044 24004
rect 5044 23948 5100 24004
rect 5100 23948 5104 24004
rect 5040 23944 5104 23948
rect 5120 24004 5184 24008
rect 5120 23948 5124 24004
rect 5124 23948 5180 24004
rect 5180 23948 5184 24004
rect 5120 23944 5184 23948
rect 5200 24004 5264 24008
rect 5200 23948 5204 24004
rect 5204 23948 5260 24004
rect 5260 23948 5264 24004
rect 5200 23944 5264 23948
rect 5280 24004 5344 24008
rect 5280 23948 5284 24004
rect 5284 23948 5340 24004
rect 5340 23948 5344 24004
rect 5280 23944 5344 23948
rect 1960 23338 2024 23342
rect 1960 23282 1964 23338
rect 1964 23282 2020 23338
rect 2020 23282 2024 23338
rect 1960 23278 2024 23282
rect 2040 23338 2104 23342
rect 2040 23282 2044 23338
rect 2044 23282 2100 23338
rect 2100 23282 2104 23338
rect 2040 23278 2104 23282
rect 2120 23338 2184 23342
rect 2120 23282 2124 23338
rect 2124 23282 2180 23338
rect 2180 23282 2184 23338
rect 2120 23278 2184 23282
rect 2200 23338 2264 23342
rect 2200 23282 2204 23338
rect 2204 23282 2260 23338
rect 2260 23282 2264 23338
rect 2200 23278 2264 23282
rect 2280 23338 2344 23342
rect 2280 23282 2284 23338
rect 2284 23282 2340 23338
rect 2340 23282 2344 23338
rect 2280 23278 2344 23282
rect 7960 23338 8024 23342
rect 7960 23282 7964 23338
rect 7964 23282 8020 23338
rect 8020 23282 8024 23338
rect 7960 23278 8024 23282
rect 8040 23338 8104 23342
rect 8040 23282 8044 23338
rect 8044 23282 8100 23338
rect 8100 23282 8104 23338
rect 8040 23278 8104 23282
rect 8120 23338 8184 23342
rect 8120 23282 8124 23338
rect 8124 23282 8180 23338
rect 8180 23282 8184 23338
rect 8120 23278 8184 23282
rect 8200 23338 8264 23342
rect 8200 23282 8204 23338
rect 8204 23282 8260 23338
rect 8260 23282 8264 23338
rect 8200 23278 8264 23282
rect 8280 23338 8344 23342
rect 8280 23282 8284 23338
rect 8284 23282 8340 23338
rect 8340 23282 8344 23338
rect 8280 23278 8344 23282
rect 4960 22672 5024 22676
rect 4960 22616 4964 22672
rect 4964 22616 5020 22672
rect 5020 22616 5024 22672
rect 4960 22612 5024 22616
rect 5040 22672 5104 22676
rect 5040 22616 5044 22672
rect 5044 22616 5100 22672
rect 5100 22616 5104 22672
rect 5040 22612 5104 22616
rect 5120 22672 5184 22676
rect 5120 22616 5124 22672
rect 5124 22616 5180 22672
rect 5180 22616 5184 22672
rect 5120 22612 5184 22616
rect 5200 22672 5264 22676
rect 5200 22616 5204 22672
rect 5204 22616 5260 22672
rect 5260 22616 5264 22672
rect 5200 22612 5264 22616
rect 5280 22672 5344 22676
rect 5280 22616 5284 22672
rect 5284 22616 5340 22672
rect 5340 22616 5344 22672
rect 5280 22612 5344 22616
rect 1960 22006 2024 22010
rect 1960 21950 1964 22006
rect 1964 21950 2020 22006
rect 2020 21950 2024 22006
rect 1960 21946 2024 21950
rect 2040 22006 2104 22010
rect 2040 21950 2044 22006
rect 2044 21950 2100 22006
rect 2100 21950 2104 22006
rect 2040 21946 2104 21950
rect 2120 22006 2184 22010
rect 2120 21950 2124 22006
rect 2124 21950 2180 22006
rect 2180 21950 2184 22006
rect 2120 21946 2184 21950
rect 2200 22006 2264 22010
rect 2200 21950 2204 22006
rect 2204 21950 2260 22006
rect 2260 21950 2264 22006
rect 2200 21946 2264 21950
rect 2280 22006 2344 22010
rect 2280 21950 2284 22006
rect 2284 21950 2340 22006
rect 2340 21950 2344 22006
rect 2280 21946 2344 21950
rect 7960 22006 8024 22010
rect 7960 21950 7964 22006
rect 7964 21950 8020 22006
rect 8020 21950 8024 22006
rect 7960 21946 8024 21950
rect 8040 22006 8104 22010
rect 8040 21950 8044 22006
rect 8044 21950 8100 22006
rect 8100 21950 8104 22006
rect 8040 21946 8104 21950
rect 8120 22006 8184 22010
rect 8120 21950 8124 22006
rect 8124 21950 8180 22006
rect 8180 21950 8184 22006
rect 8120 21946 8184 21950
rect 8200 22006 8264 22010
rect 8200 21950 8204 22006
rect 8204 21950 8260 22006
rect 8260 21950 8264 22006
rect 8200 21946 8264 21950
rect 8280 22006 8344 22010
rect 8280 21950 8284 22006
rect 8284 21950 8340 22006
rect 8340 21950 8344 22006
rect 8280 21946 8344 21950
rect 4960 21340 5024 21344
rect 4960 21284 4964 21340
rect 4964 21284 5020 21340
rect 5020 21284 5024 21340
rect 4960 21280 5024 21284
rect 5040 21340 5104 21344
rect 5040 21284 5044 21340
rect 5044 21284 5100 21340
rect 5100 21284 5104 21340
rect 5040 21280 5104 21284
rect 5120 21340 5184 21344
rect 5120 21284 5124 21340
rect 5124 21284 5180 21340
rect 5180 21284 5184 21340
rect 5120 21280 5184 21284
rect 5200 21340 5264 21344
rect 5200 21284 5204 21340
rect 5204 21284 5260 21340
rect 5260 21284 5264 21340
rect 5200 21280 5264 21284
rect 5280 21340 5344 21344
rect 5280 21284 5284 21340
rect 5284 21284 5340 21340
rect 5340 21284 5344 21340
rect 5280 21280 5344 21284
rect 1960 20674 2024 20678
rect 1960 20618 1964 20674
rect 1964 20618 2020 20674
rect 2020 20618 2024 20674
rect 1960 20614 2024 20618
rect 2040 20674 2104 20678
rect 2040 20618 2044 20674
rect 2044 20618 2100 20674
rect 2100 20618 2104 20674
rect 2040 20614 2104 20618
rect 2120 20674 2184 20678
rect 2120 20618 2124 20674
rect 2124 20618 2180 20674
rect 2180 20618 2184 20674
rect 2120 20614 2184 20618
rect 2200 20674 2264 20678
rect 2200 20618 2204 20674
rect 2204 20618 2260 20674
rect 2260 20618 2264 20674
rect 2200 20614 2264 20618
rect 2280 20674 2344 20678
rect 2280 20618 2284 20674
rect 2284 20618 2340 20674
rect 2340 20618 2344 20674
rect 2280 20614 2344 20618
rect 7960 20674 8024 20678
rect 7960 20618 7964 20674
rect 7964 20618 8020 20674
rect 8020 20618 8024 20674
rect 7960 20614 8024 20618
rect 8040 20674 8104 20678
rect 8040 20618 8044 20674
rect 8044 20618 8100 20674
rect 8100 20618 8104 20674
rect 8040 20614 8104 20618
rect 8120 20674 8184 20678
rect 8120 20618 8124 20674
rect 8124 20618 8180 20674
rect 8180 20618 8184 20674
rect 8120 20614 8184 20618
rect 8200 20674 8264 20678
rect 8200 20618 8204 20674
rect 8204 20618 8260 20674
rect 8260 20618 8264 20674
rect 8200 20614 8264 20618
rect 8280 20674 8344 20678
rect 8280 20618 8284 20674
rect 8284 20618 8340 20674
rect 8340 20618 8344 20674
rect 8280 20614 8344 20618
rect 4960 20008 5024 20012
rect 4960 19952 4964 20008
rect 4964 19952 5020 20008
rect 5020 19952 5024 20008
rect 4960 19948 5024 19952
rect 5040 20008 5104 20012
rect 5040 19952 5044 20008
rect 5044 19952 5100 20008
rect 5100 19952 5104 20008
rect 5040 19948 5104 19952
rect 5120 20008 5184 20012
rect 5120 19952 5124 20008
rect 5124 19952 5180 20008
rect 5180 19952 5184 20008
rect 5120 19948 5184 19952
rect 5200 20008 5264 20012
rect 5200 19952 5204 20008
rect 5204 19952 5260 20008
rect 5260 19952 5264 20008
rect 5200 19948 5264 19952
rect 5280 20008 5344 20012
rect 5280 19952 5284 20008
rect 5284 19952 5340 20008
rect 5340 19952 5344 20008
rect 5280 19948 5344 19952
rect 1960 19342 2024 19346
rect 1960 19286 1964 19342
rect 1964 19286 2020 19342
rect 2020 19286 2024 19342
rect 1960 19282 2024 19286
rect 2040 19342 2104 19346
rect 2040 19286 2044 19342
rect 2044 19286 2100 19342
rect 2100 19286 2104 19342
rect 2040 19282 2104 19286
rect 2120 19342 2184 19346
rect 2120 19286 2124 19342
rect 2124 19286 2180 19342
rect 2180 19286 2184 19342
rect 2120 19282 2184 19286
rect 2200 19342 2264 19346
rect 2200 19286 2204 19342
rect 2204 19286 2260 19342
rect 2260 19286 2264 19342
rect 2200 19282 2264 19286
rect 2280 19342 2344 19346
rect 2280 19286 2284 19342
rect 2284 19286 2340 19342
rect 2340 19286 2344 19342
rect 2280 19282 2344 19286
rect 7960 19342 8024 19346
rect 7960 19286 7964 19342
rect 7964 19286 8020 19342
rect 8020 19286 8024 19342
rect 7960 19282 8024 19286
rect 8040 19342 8104 19346
rect 8040 19286 8044 19342
rect 8044 19286 8100 19342
rect 8100 19286 8104 19342
rect 8040 19282 8104 19286
rect 8120 19342 8184 19346
rect 8120 19286 8124 19342
rect 8124 19286 8180 19342
rect 8180 19286 8184 19342
rect 8120 19282 8184 19286
rect 8200 19342 8264 19346
rect 8200 19286 8204 19342
rect 8204 19286 8260 19342
rect 8260 19286 8264 19342
rect 8200 19282 8264 19286
rect 8280 19342 8344 19346
rect 8280 19286 8284 19342
rect 8284 19286 8340 19342
rect 8340 19286 8344 19342
rect 8280 19282 8344 19286
rect 4960 18676 5024 18680
rect 4960 18620 4964 18676
rect 4964 18620 5020 18676
rect 5020 18620 5024 18676
rect 4960 18616 5024 18620
rect 5040 18676 5104 18680
rect 5040 18620 5044 18676
rect 5044 18620 5100 18676
rect 5100 18620 5104 18676
rect 5040 18616 5104 18620
rect 5120 18676 5184 18680
rect 5120 18620 5124 18676
rect 5124 18620 5180 18676
rect 5180 18620 5184 18676
rect 5120 18616 5184 18620
rect 5200 18676 5264 18680
rect 5200 18620 5204 18676
rect 5204 18620 5260 18676
rect 5260 18620 5264 18676
rect 5200 18616 5264 18620
rect 5280 18676 5344 18680
rect 5280 18620 5284 18676
rect 5284 18620 5340 18676
rect 5340 18620 5344 18676
rect 5280 18616 5344 18620
rect 1960 18010 2024 18014
rect 1960 17954 1964 18010
rect 1964 17954 2020 18010
rect 2020 17954 2024 18010
rect 1960 17950 2024 17954
rect 2040 18010 2104 18014
rect 2040 17954 2044 18010
rect 2044 17954 2100 18010
rect 2100 17954 2104 18010
rect 2040 17950 2104 17954
rect 2120 18010 2184 18014
rect 2120 17954 2124 18010
rect 2124 17954 2180 18010
rect 2180 17954 2184 18010
rect 2120 17950 2184 17954
rect 2200 18010 2264 18014
rect 2200 17954 2204 18010
rect 2204 17954 2260 18010
rect 2260 17954 2264 18010
rect 2200 17950 2264 17954
rect 2280 18010 2344 18014
rect 2280 17954 2284 18010
rect 2284 17954 2340 18010
rect 2340 17954 2344 18010
rect 2280 17950 2344 17954
rect 7960 18010 8024 18014
rect 7960 17954 7964 18010
rect 7964 17954 8020 18010
rect 8020 17954 8024 18010
rect 7960 17950 8024 17954
rect 8040 18010 8104 18014
rect 8040 17954 8044 18010
rect 8044 17954 8100 18010
rect 8100 17954 8104 18010
rect 8040 17950 8104 17954
rect 8120 18010 8184 18014
rect 8120 17954 8124 18010
rect 8124 17954 8180 18010
rect 8180 17954 8184 18010
rect 8120 17950 8184 17954
rect 8200 18010 8264 18014
rect 8200 17954 8204 18010
rect 8204 17954 8260 18010
rect 8260 17954 8264 18010
rect 8200 17950 8264 17954
rect 8280 18010 8344 18014
rect 8280 17954 8284 18010
rect 8284 17954 8340 18010
rect 8340 17954 8344 18010
rect 8280 17950 8344 17954
rect 4960 17344 5024 17348
rect 4960 17288 4964 17344
rect 4964 17288 5020 17344
rect 5020 17288 5024 17344
rect 4960 17284 5024 17288
rect 5040 17344 5104 17348
rect 5040 17288 5044 17344
rect 5044 17288 5100 17344
rect 5100 17288 5104 17344
rect 5040 17284 5104 17288
rect 5120 17344 5184 17348
rect 5120 17288 5124 17344
rect 5124 17288 5180 17344
rect 5180 17288 5184 17344
rect 5120 17284 5184 17288
rect 5200 17344 5264 17348
rect 5200 17288 5204 17344
rect 5204 17288 5260 17344
rect 5260 17288 5264 17344
rect 5200 17284 5264 17288
rect 5280 17344 5344 17348
rect 5280 17288 5284 17344
rect 5284 17288 5340 17344
rect 5340 17288 5344 17344
rect 5280 17284 5344 17288
rect 1960 16678 2024 16682
rect 1960 16622 1964 16678
rect 1964 16622 2020 16678
rect 2020 16622 2024 16678
rect 1960 16618 2024 16622
rect 2040 16678 2104 16682
rect 2040 16622 2044 16678
rect 2044 16622 2100 16678
rect 2100 16622 2104 16678
rect 2040 16618 2104 16622
rect 2120 16678 2184 16682
rect 2120 16622 2124 16678
rect 2124 16622 2180 16678
rect 2180 16622 2184 16678
rect 2120 16618 2184 16622
rect 2200 16678 2264 16682
rect 2200 16622 2204 16678
rect 2204 16622 2260 16678
rect 2260 16622 2264 16678
rect 2200 16618 2264 16622
rect 2280 16678 2344 16682
rect 2280 16622 2284 16678
rect 2284 16622 2340 16678
rect 2340 16622 2344 16678
rect 2280 16618 2344 16622
rect 7960 16678 8024 16682
rect 7960 16622 7964 16678
rect 7964 16622 8020 16678
rect 8020 16622 8024 16678
rect 7960 16618 8024 16622
rect 8040 16678 8104 16682
rect 8040 16622 8044 16678
rect 8044 16622 8100 16678
rect 8100 16622 8104 16678
rect 8040 16618 8104 16622
rect 8120 16678 8184 16682
rect 8120 16622 8124 16678
rect 8124 16622 8180 16678
rect 8180 16622 8184 16678
rect 8120 16618 8184 16622
rect 8200 16678 8264 16682
rect 8200 16622 8204 16678
rect 8204 16622 8260 16678
rect 8260 16622 8264 16678
rect 8200 16618 8264 16622
rect 8280 16678 8344 16682
rect 8280 16622 8284 16678
rect 8284 16622 8340 16678
rect 8340 16622 8344 16678
rect 8280 16618 8344 16622
rect 4960 16012 5024 16016
rect 4960 15956 4964 16012
rect 4964 15956 5020 16012
rect 5020 15956 5024 16012
rect 4960 15952 5024 15956
rect 5040 16012 5104 16016
rect 5040 15956 5044 16012
rect 5044 15956 5100 16012
rect 5100 15956 5104 16012
rect 5040 15952 5104 15956
rect 5120 16012 5184 16016
rect 5120 15956 5124 16012
rect 5124 15956 5180 16012
rect 5180 15956 5184 16012
rect 5120 15952 5184 15956
rect 5200 16012 5264 16016
rect 5200 15956 5204 16012
rect 5204 15956 5260 16012
rect 5260 15956 5264 16012
rect 5200 15952 5264 15956
rect 5280 16012 5344 16016
rect 5280 15956 5284 16012
rect 5284 15956 5340 16012
rect 5340 15956 5344 16012
rect 5280 15952 5344 15956
rect 1960 15346 2024 15350
rect 1960 15290 1964 15346
rect 1964 15290 2020 15346
rect 2020 15290 2024 15346
rect 1960 15286 2024 15290
rect 2040 15346 2104 15350
rect 2040 15290 2044 15346
rect 2044 15290 2100 15346
rect 2100 15290 2104 15346
rect 2040 15286 2104 15290
rect 2120 15346 2184 15350
rect 2120 15290 2124 15346
rect 2124 15290 2180 15346
rect 2180 15290 2184 15346
rect 2120 15286 2184 15290
rect 2200 15346 2264 15350
rect 2200 15290 2204 15346
rect 2204 15290 2260 15346
rect 2260 15290 2264 15346
rect 2200 15286 2264 15290
rect 2280 15346 2344 15350
rect 2280 15290 2284 15346
rect 2284 15290 2340 15346
rect 2340 15290 2344 15346
rect 2280 15286 2344 15290
rect 7960 15346 8024 15350
rect 7960 15290 7964 15346
rect 7964 15290 8020 15346
rect 8020 15290 8024 15346
rect 7960 15286 8024 15290
rect 8040 15346 8104 15350
rect 8040 15290 8044 15346
rect 8044 15290 8100 15346
rect 8100 15290 8104 15346
rect 8040 15286 8104 15290
rect 8120 15346 8184 15350
rect 8120 15290 8124 15346
rect 8124 15290 8180 15346
rect 8180 15290 8184 15346
rect 8120 15286 8184 15290
rect 8200 15346 8264 15350
rect 8200 15290 8204 15346
rect 8204 15290 8260 15346
rect 8260 15290 8264 15346
rect 8200 15286 8264 15290
rect 8280 15346 8344 15350
rect 8280 15290 8284 15346
rect 8284 15290 8340 15346
rect 8340 15290 8344 15346
rect 8280 15286 8344 15290
rect 4960 14680 5024 14684
rect 4960 14624 4964 14680
rect 4964 14624 5020 14680
rect 5020 14624 5024 14680
rect 4960 14620 5024 14624
rect 5040 14680 5104 14684
rect 5040 14624 5044 14680
rect 5044 14624 5100 14680
rect 5100 14624 5104 14680
rect 5040 14620 5104 14624
rect 5120 14680 5184 14684
rect 5120 14624 5124 14680
rect 5124 14624 5180 14680
rect 5180 14624 5184 14680
rect 5120 14620 5184 14624
rect 5200 14680 5264 14684
rect 5200 14624 5204 14680
rect 5204 14624 5260 14680
rect 5260 14624 5264 14680
rect 5200 14620 5264 14624
rect 5280 14680 5344 14684
rect 5280 14624 5284 14680
rect 5284 14624 5340 14680
rect 5340 14624 5344 14680
rect 5280 14620 5344 14624
rect 1960 14014 2024 14018
rect 1960 13958 1964 14014
rect 1964 13958 2020 14014
rect 2020 13958 2024 14014
rect 1960 13954 2024 13958
rect 2040 14014 2104 14018
rect 2040 13958 2044 14014
rect 2044 13958 2100 14014
rect 2100 13958 2104 14014
rect 2040 13954 2104 13958
rect 2120 14014 2184 14018
rect 2120 13958 2124 14014
rect 2124 13958 2180 14014
rect 2180 13958 2184 14014
rect 2120 13954 2184 13958
rect 2200 14014 2264 14018
rect 2200 13958 2204 14014
rect 2204 13958 2260 14014
rect 2260 13958 2264 14014
rect 2200 13954 2264 13958
rect 2280 14014 2344 14018
rect 2280 13958 2284 14014
rect 2284 13958 2340 14014
rect 2340 13958 2344 14014
rect 2280 13954 2344 13958
rect 7960 14014 8024 14018
rect 7960 13958 7964 14014
rect 7964 13958 8020 14014
rect 8020 13958 8024 14014
rect 7960 13954 8024 13958
rect 8040 14014 8104 14018
rect 8040 13958 8044 14014
rect 8044 13958 8100 14014
rect 8100 13958 8104 14014
rect 8040 13954 8104 13958
rect 8120 14014 8184 14018
rect 8120 13958 8124 14014
rect 8124 13958 8180 14014
rect 8180 13958 8184 14014
rect 8120 13954 8184 13958
rect 8200 14014 8264 14018
rect 8200 13958 8204 14014
rect 8204 13958 8260 14014
rect 8260 13958 8264 14014
rect 8200 13954 8264 13958
rect 8280 14014 8344 14018
rect 8280 13958 8284 14014
rect 8284 13958 8340 14014
rect 8340 13958 8344 14014
rect 8280 13954 8344 13958
rect 4960 13348 5024 13352
rect 4960 13292 4964 13348
rect 4964 13292 5020 13348
rect 5020 13292 5024 13348
rect 4960 13288 5024 13292
rect 5040 13348 5104 13352
rect 5040 13292 5044 13348
rect 5044 13292 5100 13348
rect 5100 13292 5104 13348
rect 5040 13288 5104 13292
rect 5120 13348 5184 13352
rect 5120 13292 5124 13348
rect 5124 13292 5180 13348
rect 5180 13292 5184 13348
rect 5120 13288 5184 13292
rect 5200 13348 5264 13352
rect 5200 13292 5204 13348
rect 5204 13292 5260 13348
rect 5260 13292 5264 13348
rect 5200 13288 5264 13292
rect 5280 13348 5344 13352
rect 5280 13292 5284 13348
rect 5284 13292 5340 13348
rect 5340 13292 5344 13348
rect 5280 13288 5344 13292
rect 1960 12682 2024 12686
rect 1960 12626 1964 12682
rect 1964 12626 2020 12682
rect 2020 12626 2024 12682
rect 1960 12622 2024 12626
rect 2040 12682 2104 12686
rect 2040 12626 2044 12682
rect 2044 12626 2100 12682
rect 2100 12626 2104 12682
rect 2040 12622 2104 12626
rect 2120 12682 2184 12686
rect 2120 12626 2124 12682
rect 2124 12626 2180 12682
rect 2180 12626 2184 12682
rect 2120 12622 2184 12626
rect 2200 12682 2264 12686
rect 2200 12626 2204 12682
rect 2204 12626 2260 12682
rect 2260 12626 2264 12682
rect 2200 12622 2264 12626
rect 2280 12682 2344 12686
rect 2280 12626 2284 12682
rect 2284 12626 2340 12682
rect 2340 12626 2344 12682
rect 2280 12622 2344 12626
rect 7960 12682 8024 12686
rect 7960 12626 7964 12682
rect 7964 12626 8020 12682
rect 8020 12626 8024 12682
rect 7960 12622 8024 12626
rect 8040 12682 8104 12686
rect 8040 12626 8044 12682
rect 8044 12626 8100 12682
rect 8100 12626 8104 12682
rect 8040 12622 8104 12626
rect 8120 12682 8184 12686
rect 8120 12626 8124 12682
rect 8124 12626 8180 12682
rect 8180 12626 8184 12682
rect 8120 12622 8184 12626
rect 8200 12682 8264 12686
rect 8200 12626 8204 12682
rect 8204 12626 8260 12682
rect 8260 12626 8264 12682
rect 8200 12622 8264 12626
rect 8280 12682 8344 12686
rect 8280 12626 8284 12682
rect 8284 12626 8340 12682
rect 8340 12626 8344 12682
rect 8280 12622 8344 12626
rect 4960 12016 5024 12020
rect 4960 11960 4964 12016
rect 4964 11960 5020 12016
rect 5020 11960 5024 12016
rect 4960 11956 5024 11960
rect 5040 12016 5104 12020
rect 5040 11960 5044 12016
rect 5044 11960 5100 12016
rect 5100 11960 5104 12016
rect 5040 11956 5104 11960
rect 5120 12016 5184 12020
rect 5120 11960 5124 12016
rect 5124 11960 5180 12016
rect 5180 11960 5184 12016
rect 5120 11956 5184 11960
rect 5200 12016 5264 12020
rect 5200 11960 5204 12016
rect 5204 11960 5260 12016
rect 5260 11960 5264 12016
rect 5200 11956 5264 11960
rect 5280 12016 5344 12020
rect 5280 11960 5284 12016
rect 5284 11960 5340 12016
rect 5340 11960 5344 12016
rect 5280 11956 5344 11960
rect 1960 11350 2024 11354
rect 1960 11294 1964 11350
rect 1964 11294 2020 11350
rect 2020 11294 2024 11350
rect 1960 11290 2024 11294
rect 2040 11350 2104 11354
rect 2040 11294 2044 11350
rect 2044 11294 2100 11350
rect 2100 11294 2104 11350
rect 2040 11290 2104 11294
rect 2120 11350 2184 11354
rect 2120 11294 2124 11350
rect 2124 11294 2180 11350
rect 2180 11294 2184 11350
rect 2120 11290 2184 11294
rect 2200 11350 2264 11354
rect 2200 11294 2204 11350
rect 2204 11294 2260 11350
rect 2260 11294 2264 11350
rect 2200 11290 2264 11294
rect 2280 11350 2344 11354
rect 2280 11294 2284 11350
rect 2284 11294 2340 11350
rect 2340 11294 2344 11350
rect 2280 11290 2344 11294
rect 7960 11350 8024 11354
rect 7960 11294 7964 11350
rect 7964 11294 8020 11350
rect 8020 11294 8024 11350
rect 7960 11290 8024 11294
rect 8040 11350 8104 11354
rect 8040 11294 8044 11350
rect 8044 11294 8100 11350
rect 8100 11294 8104 11350
rect 8040 11290 8104 11294
rect 8120 11350 8184 11354
rect 8120 11294 8124 11350
rect 8124 11294 8180 11350
rect 8180 11294 8184 11350
rect 8120 11290 8184 11294
rect 8200 11350 8264 11354
rect 8200 11294 8204 11350
rect 8204 11294 8260 11350
rect 8260 11294 8264 11350
rect 8200 11290 8264 11294
rect 8280 11350 8344 11354
rect 8280 11294 8284 11350
rect 8284 11294 8340 11350
rect 8340 11294 8344 11350
rect 8280 11290 8344 11294
rect 4960 10684 5024 10688
rect 4960 10628 4964 10684
rect 4964 10628 5020 10684
rect 5020 10628 5024 10684
rect 4960 10624 5024 10628
rect 5040 10684 5104 10688
rect 5040 10628 5044 10684
rect 5044 10628 5100 10684
rect 5100 10628 5104 10684
rect 5040 10624 5104 10628
rect 5120 10684 5184 10688
rect 5120 10628 5124 10684
rect 5124 10628 5180 10684
rect 5180 10628 5184 10684
rect 5120 10624 5184 10628
rect 5200 10684 5264 10688
rect 5200 10628 5204 10684
rect 5204 10628 5260 10684
rect 5260 10628 5264 10684
rect 5200 10624 5264 10628
rect 5280 10684 5344 10688
rect 5280 10628 5284 10684
rect 5284 10628 5340 10684
rect 5340 10628 5344 10684
rect 5280 10624 5344 10628
rect 1960 10018 2024 10022
rect 1960 9962 1964 10018
rect 1964 9962 2020 10018
rect 2020 9962 2024 10018
rect 1960 9958 2024 9962
rect 2040 10018 2104 10022
rect 2040 9962 2044 10018
rect 2044 9962 2100 10018
rect 2100 9962 2104 10018
rect 2040 9958 2104 9962
rect 2120 10018 2184 10022
rect 2120 9962 2124 10018
rect 2124 9962 2180 10018
rect 2180 9962 2184 10018
rect 2120 9958 2184 9962
rect 2200 10018 2264 10022
rect 2200 9962 2204 10018
rect 2204 9962 2260 10018
rect 2260 9962 2264 10018
rect 2200 9958 2264 9962
rect 2280 10018 2344 10022
rect 2280 9962 2284 10018
rect 2284 9962 2340 10018
rect 2340 9962 2344 10018
rect 2280 9958 2344 9962
rect 7960 10018 8024 10022
rect 7960 9962 7964 10018
rect 7964 9962 8020 10018
rect 8020 9962 8024 10018
rect 7960 9958 8024 9962
rect 8040 10018 8104 10022
rect 8040 9962 8044 10018
rect 8044 9962 8100 10018
rect 8100 9962 8104 10018
rect 8040 9958 8104 9962
rect 8120 10018 8184 10022
rect 8120 9962 8124 10018
rect 8124 9962 8180 10018
rect 8180 9962 8184 10018
rect 8120 9958 8184 9962
rect 8200 10018 8264 10022
rect 8200 9962 8204 10018
rect 8204 9962 8260 10018
rect 8260 9962 8264 10018
rect 8200 9958 8264 9962
rect 8280 10018 8344 10022
rect 8280 9962 8284 10018
rect 8284 9962 8340 10018
rect 8340 9962 8344 10018
rect 8280 9958 8344 9962
rect 4960 9352 5024 9356
rect 4960 9296 4964 9352
rect 4964 9296 5020 9352
rect 5020 9296 5024 9352
rect 4960 9292 5024 9296
rect 5040 9352 5104 9356
rect 5040 9296 5044 9352
rect 5044 9296 5100 9352
rect 5100 9296 5104 9352
rect 5040 9292 5104 9296
rect 5120 9352 5184 9356
rect 5120 9296 5124 9352
rect 5124 9296 5180 9352
rect 5180 9296 5184 9352
rect 5120 9292 5184 9296
rect 5200 9352 5264 9356
rect 5200 9296 5204 9352
rect 5204 9296 5260 9352
rect 5260 9296 5264 9352
rect 5200 9292 5264 9296
rect 5280 9352 5344 9356
rect 5280 9296 5284 9352
rect 5284 9296 5340 9352
rect 5340 9296 5344 9352
rect 5280 9292 5344 9296
rect 1960 8686 2024 8690
rect 1960 8630 1964 8686
rect 1964 8630 2020 8686
rect 2020 8630 2024 8686
rect 1960 8626 2024 8630
rect 2040 8686 2104 8690
rect 2040 8630 2044 8686
rect 2044 8630 2100 8686
rect 2100 8630 2104 8686
rect 2040 8626 2104 8630
rect 2120 8686 2184 8690
rect 2120 8630 2124 8686
rect 2124 8630 2180 8686
rect 2180 8630 2184 8686
rect 2120 8626 2184 8630
rect 2200 8686 2264 8690
rect 2200 8630 2204 8686
rect 2204 8630 2260 8686
rect 2260 8630 2264 8686
rect 2200 8626 2264 8630
rect 2280 8686 2344 8690
rect 2280 8630 2284 8686
rect 2284 8630 2340 8686
rect 2340 8630 2344 8686
rect 2280 8626 2344 8630
rect 7960 8686 8024 8690
rect 7960 8630 7964 8686
rect 7964 8630 8020 8686
rect 8020 8630 8024 8686
rect 7960 8626 8024 8630
rect 8040 8686 8104 8690
rect 8040 8630 8044 8686
rect 8044 8630 8100 8686
rect 8100 8630 8104 8686
rect 8040 8626 8104 8630
rect 8120 8686 8184 8690
rect 8120 8630 8124 8686
rect 8124 8630 8180 8686
rect 8180 8630 8184 8686
rect 8120 8626 8184 8630
rect 8200 8686 8264 8690
rect 8200 8630 8204 8686
rect 8204 8630 8260 8686
rect 8260 8630 8264 8686
rect 8200 8626 8264 8630
rect 8280 8686 8344 8690
rect 8280 8630 8284 8686
rect 8284 8630 8340 8686
rect 8340 8630 8344 8686
rect 8280 8626 8344 8630
rect 4960 8020 5024 8024
rect 4960 7964 4964 8020
rect 4964 7964 5020 8020
rect 5020 7964 5024 8020
rect 4960 7960 5024 7964
rect 5040 8020 5104 8024
rect 5040 7964 5044 8020
rect 5044 7964 5100 8020
rect 5100 7964 5104 8020
rect 5040 7960 5104 7964
rect 5120 8020 5184 8024
rect 5120 7964 5124 8020
rect 5124 7964 5180 8020
rect 5180 7964 5184 8020
rect 5120 7960 5184 7964
rect 5200 8020 5264 8024
rect 5200 7964 5204 8020
rect 5204 7964 5260 8020
rect 5260 7964 5264 8020
rect 5200 7960 5264 7964
rect 5280 8020 5344 8024
rect 5280 7964 5284 8020
rect 5284 7964 5340 8020
rect 5340 7964 5344 8020
rect 5280 7960 5344 7964
rect 1960 7354 2024 7358
rect 1960 7298 1964 7354
rect 1964 7298 2020 7354
rect 2020 7298 2024 7354
rect 1960 7294 2024 7298
rect 2040 7354 2104 7358
rect 2040 7298 2044 7354
rect 2044 7298 2100 7354
rect 2100 7298 2104 7354
rect 2040 7294 2104 7298
rect 2120 7354 2184 7358
rect 2120 7298 2124 7354
rect 2124 7298 2180 7354
rect 2180 7298 2184 7354
rect 2120 7294 2184 7298
rect 2200 7354 2264 7358
rect 2200 7298 2204 7354
rect 2204 7298 2260 7354
rect 2260 7298 2264 7354
rect 2200 7294 2264 7298
rect 2280 7354 2344 7358
rect 2280 7298 2284 7354
rect 2284 7298 2340 7354
rect 2340 7298 2344 7354
rect 2280 7294 2344 7298
rect 7960 7354 8024 7358
rect 7960 7298 7964 7354
rect 7964 7298 8020 7354
rect 8020 7298 8024 7354
rect 7960 7294 8024 7298
rect 8040 7354 8104 7358
rect 8040 7298 8044 7354
rect 8044 7298 8100 7354
rect 8100 7298 8104 7354
rect 8040 7294 8104 7298
rect 8120 7354 8184 7358
rect 8120 7298 8124 7354
rect 8124 7298 8180 7354
rect 8180 7298 8184 7354
rect 8120 7294 8184 7298
rect 8200 7354 8264 7358
rect 8200 7298 8204 7354
rect 8204 7298 8260 7354
rect 8260 7298 8264 7354
rect 8200 7294 8264 7298
rect 8280 7354 8344 7358
rect 8280 7298 8284 7354
rect 8284 7298 8340 7354
rect 8340 7298 8344 7354
rect 8280 7294 8344 7298
rect 4960 6688 5024 6692
rect 4960 6632 4964 6688
rect 4964 6632 5020 6688
rect 5020 6632 5024 6688
rect 4960 6628 5024 6632
rect 5040 6688 5104 6692
rect 5040 6632 5044 6688
rect 5044 6632 5100 6688
rect 5100 6632 5104 6688
rect 5040 6628 5104 6632
rect 5120 6688 5184 6692
rect 5120 6632 5124 6688
rect 5124 6632 5180 6688
rect 5180 6632 5184 6688
rect 5120 6628 5184 6632
rect 5200 6688 5264 6692
rect 5200 6632 5204 6688
rect 5204 6632 5260 6688
rect 5260 6632 5264 6688
rect 5200 6628 5264 6632
rect 5280 6688 5344 6692
rect 5280 6632 5284 6688
rect 5284 6632 5340 6688
rect 5340 6632 5344 6688
rect 5280 6628 5344 6632
rect 1960 6022 2024 6026
rect 1960 5966 1964 6022
rect 1964 5966 2020 6022
rect 2020 5966 2024 6022
rect 1960 5962 2024 5966
rect 2040 6022 2104 6026
rect 2040 5966 2044 6022
rect 2044 5966 2100 6022
rect 2100 5966 2104 6022
rect 2040 5962 2104 5966
rect 2120 6022 2184 6026
rect 2120 5966 2124 6022
rect 2124 5966 2180 6022
rect 2180 5966 2184 6022
rect 2120 5962 2184 5966
rect 2200 6022 2264 6026
rect 2200 5966 2204 6022
rect 2204 5966 2260 6022
rect 2260 5966 2264 6022
rect 2200 5962 2264 5966
rect 2280 6022 2344 6026
rect 2280 5966 2284 6022
rect 2284 5966 2340 6022
rect 2340 5966 2344 6022
rect 2280 5962 2344 5966
rect 7960 6022 8024 6026
rect 7960 5966 7964 6022
rect 7964 5966 8020 6022
rect 8020 5966 8024 6022
rect 7960 5962 8024 5966
rect 8040 6022 8104 6026
rect 8040 5966 8044 6022
rect 8044 5966 8100 6022
rect 8100 5966 8104 6022
rect 8040 5962 8104 5966
rect 8120 6022 8184 6026
rect 8120 5966 8124 6022
rect 8124 5966 8180 6022
rect 8180 5966 8184 6022
rect 8120 5962 8184 5966
rect 8200 6022 8264 6026
rect 8200 5966 8204 6022
rect 8204 5966 8260 6022
rect 8260 5966 8264 6022
rect 8200 5962 8264 5966
rect 8280 6022 8344 6026
rect 8280 5966 8284 6022
rect 8284 5966 8340 6022
rect 8340 5966 8344 6022
rect 8280 5962 8344 5966
rect 4960 5356 5024 5360
rect 4960 5300 4964 5356
rect 4964 5300 5020 5356
rect 5020 5300 5024 5356
rect 4960 5296 5024 5300
rect 5040 5356 5104 5360
rect 5040 5300 5044 5356
rect 5044 5300 5100 5356
rect 5100 5300 5104 5356
rect 5040 5296 5104 5300
rect 5120 5356 5184 5360
rect 5120 5300 5124 5356
rect 5124 5300 5180 5356
rect 5180 5300 5184 5356
rect 5120 5296 5184 5300
rect 5200 5356 5264 5360
rect 5200 5300 5204 5356
rect 5204 5300 5260 5356
rect 5260 5300 5264 5356
rect 5200 5296 5264 5300
rect 5280 5356 5344 5360
rect 5280 5300 5284 5356
rect 5284 5300 5340 5356
rect 5340 5300 5344 5356
rect 5280 5296 5344 5300
rect 1960 4690 2024 4694
rect 1960 4634 1964 4690
rect 1964 4634 2020 4690
rect 2020 4634 2024 4690
rect 1960 4630 2024 4634
rect 2040 4690 2104 4694
rect 2040 4634 2044 4690
rect 2044 4634 2100 4690
rect 2100 4634 2104 4690
rect 2040 4630 2104 4634
rect 2120 4690 2184 4694
rect 2120 4634 2124 4690
rect 2124 4634 2180 4690
rect 2180 4634 2184 4690
rect 2120 4630 2184 4634
rect 2200 4690 2264 4694
rect 2200 4634 2204 4690
rect 2204 4634 2260 4690
rect 2260 4634 2264 4690
rect 2200 4630 2264 4634
rect 2280 4690 2344 4694
rect 2280 4634 2284 4690
rect 2284 4634 2340 4690
rect 2340 4634 2344 4690
rect 2280 4630 2344 4634
rect 7960 4690 8024 4694
rect 7960 4634 7964 4690
rect 7964 4634 8020 4690
rect 8020 4634 8024 4690
rect 7960 4630 8024 4634
rect 8040 4690 8104 4694
rect 8040 4634 8044 4690
rect 8044 4634 8100 4690
rect 8100 4634 8104 4690
rect 8040 4630 8104 4634
rect 8120 4690 8184 4694
rect 8120 4634 8124 4690
rect 8124 4634 8180 4690
rect 8180 4634 8184 4690
rect 8120 4630 8184 4634
rect 8200 4690 8264 4694
rect 8200 4634 8204 4690
rect 8204 4634 8260 4690
rect 8260 4634 8264 4690
rect 8200 4630 8264 4634
rect 8280 4690 8344 4694
rect 8280 4634 8284 4690
rect 8284 4634 8340 4690
rect 8340 4634 8344 4690
rect 8280 4630 8344 4634
rect 4960 4024 5024 4028
rect 4960 3968 4964 4024
rect 4964 3968 5020 4024
rect 5020 3968 5024 4024
rect 4960 3964 5024 3968
rect 5040 4024 5104 4028
rect 5040 3968 5044 4024
rect 5044 3968 5100 4024
rect 5100 3968 5104 4024
rect 5040 3964 5104 3968
rect 5120 4024 5184 4028
rect 5120 3968 5124 4024
rect 5124 3968 5180 4024
rect 5180 3968 5184 4024
rect 5120 3964 5184 3968
rect 5200 4024 5264 4028
rect 5200 3968 5204 4024
rect 5204 3968 5260 4024
rect 5260 3968 5264 4024
rect 5200 3964 5264 3968
rect 5280 4024 5344 4028
rect 5280 3968 5284 4024
rect 5284 3968 5340 4024
rect 5340 3968 5344 4024
rect 5280 3964 5344 3968
rect 1960 3358 2024 3362
rect 1960 3302 1964 3358
rect 1964 3302 2020 3358
rect 2020 3302 2024 3358
rect 1960 3298 2024 3302
rect 2040 3358 2104 3362
rect 2040 3302 2044 3358
rect 2044 3302 2100 3358
rect 2100 3302 2104 3358
rect 2040 3298 2104 3302
rect 2120 3358 2184 3362
rect 2120 3302 2124 3358
rect 2124 3302 2180 3358
rect 2180 3302 2184 3358
rect 2120 3298 2184 3302
rect 2200 3358 2264 3362
rect 2200 3302 2204 3358
rect 2204 3302 2260 3358
rect 2260 3302 2264 3358
rect 2200 3298 2264 3302
rect 2280 3358 2344 3362
rect 2280 3302 2284 3358
rect 2284 3302 2340 3358
rect 2340 3302 2344 3358
rect 2280 3298 2344 3302
rect 7960 3358 8024 3362
rect 7960 3302 7964 3358
rect 7964 3302 8020 3358
rect 8020 3302 8024 3358
rect 7960 3298 8024 3302
rect 8040 3358 8104 3362
rect 8040 3302 8044 3358
rect 8044 3302 8100 3358
rect 8100 3302 8104 3358
rect 8040 3298 8104 3302
rect 8120 3358 8184 3362
rect 8120 3302 8124 3358
rect 8124 3302 8180 3358
rect 8180 3302 8184 3358
rect 8120 3298 8184 3302
rect 8200 3358 8264 3362
rect 8200 3302 8204 3358
rect 8204 3302 8260 3358
rect 8260 3302 8264 3358
rect 8200 3298 8264 3302
rect 8280 3358 8344 3362
rect 8280 3302 8284 3358
rect 8284 3302 8340 3358
rect 8340 3302 8344 3358
rect 8280 3298 8344 3302
rect 4960 2692 5024 2696
rect 4960 2636 4964 2692
rect 4964 2636 5020 2692
rect 5020 2636 5024 2692
rect 4960 2632 5024 2636
rect 5040 2692 5104 2696
rect 5040 2636 5044 2692
rect 5044 2636 5100 2692
rect 5100 2636 5104 2692
rect 5040 2632 5104 2636
rect 5120 2692 5184 2696
rect 5120 2636 5124 2692
rect 5124 2636 5180 2692
rect 5180 2636 5184 2692
rect 5120 2632 5184 2636
rect 5200 2692 5264 2696
rect 5200 2636 5204 2692
rect 5204 2636 5260 2692
rect 5260 2636 5264 2692
rect 5200 2632 5264 2636
rect 5280 2692 5344 2696
rect 5280 2636 5284 2692
rect 5284 2636 5340 2692
rect 5340 2636 5344 2692
rect 5280 2632 5344 2636
<< metal4 >>
rect 1952 26006 2352 26022
rect 1952 25942 1960 26006
rect 2024 25942 2040 26006
rect 2104 25942 2120 26006
rect 2184 25942 2200 26006
rect 2264 25942 2280 26006
rect 2344 25942 2352 26006
rect 1952 24674 2352 25942
rect 1952 24610 1960 24674
rect 2024 24610 2040 24674
rect 2104 24610 2120 24674
rect 2184 24610 2200 24674
rect 2264 24610 2280 24674
rect 2344 24610 2352 24674
rect 1952 23342 2352 24610
rect 1952 23278 1960 23342
rect 2024 23278 2040 23342
rect 2104 23278 2120 23342
rect 2184 23278 2200 23342
rect 2264 23278 2280 23342
rect 2344 23278 2352 23342
rect 1952 22010 2352 23278
rect 1952 21946 1960 22010
rect 2024 21946 2040 22010
rect 2104 21946 2120 22010
rect 2184 21946 2200 22010
rect 2264 21946 2280 22010
rect 2344 21946 2352 22010
rect 1952 20678 2352 21946
rect 1952 20614 1960 20678
rect 2024 20614 2040 20678
rect 2104 20614 2120 20678
rect 2184 20614 2200 20678
rect 2264 20614 2280 20678
rect 2344 20614 2352 20678
rect 1952 19346 2352 20614
rect 1952 19282 1960 19346
rect 2024 19282 2040 19346
rect 2104 19282 2120 19346
rect 2184 19282 2200 19346
rect 2264 19282 2280 19346
rect 2344 19282 2352 19346
rect 1952 18014 2352 19282
rect 1952 17950 1960 18014
rect 2024 17950 2040 18014
rect 2104 17950 2120 18014
rect 2184 17950 2200 18014
rect 2264 17950 2280 18014
rect 2344 17950 2352 18014
rect 1952 16682 2352 17950
rect 1952 16618 1960 16682
rect 2024 16618 2040 16682
rect 2104 16618 2120 16682
rect 2184 16618 2200 16682
rect 2264 16618 2280 16682
rect 2344 16618 2352 16682
rect 1952 15350 2352 16618
rect 1952 15286 1960 15350
rect 2024 15286 2040 15350
rect 2104 15286 2120 15350
rect 2184 15286 2200 15350
rect 2264 15286 2280 15350
rect 2344 15286 2352 15350
rect 1952 14018 2352 15286
rect 1952 13954 1960 14018
rect 2024 13954 2040 14018
rect 2104 13954 2120 14018
rect 2184 13954 2200 14018
rect 2264 13954 2280 14018
rect 2344 13954 2352 14018
rect 1952 12686 2352 13954
rect 1952 12622 1960 12686
rect 2024 12622 2040 12686
rect 2104 12622 2120 12686
rect 2184 12622 2200 12686
rect 2264 12622 2280 12686
rect 2344 12622 2352 12686
rect 1952 11354 2352 12622
rect 1952 11290 1960 11354
rect 2024 11290 2040 11354
rect 2104 11290 2120 11354
rect 2184 11290 2200 11354
rect 2264 11290 2280 11354
rect 2344 11290 2352 11354
rect 1952 10022 2352 11290
rect 1952 9958 1960 10022
rect 2024 9958 2040 10022
rect 2104 9958 2120 10022
rect 2184 9958 2200 10022
rect 2264 9958 2280 10022
rect 2344 9958 2352 10022
rect 1952 8690 2352 9958
rect 1952 8626 1960 8690
rect 2024 8626 2040 8690
rect 2104 8626 2120 8690
rect 2184 8626 2200 8690
rect 2264 8626 2280 8690
rect 2344 8626 2352 8690
rect 1952 7358 2352 8626
rect 1952 7294 1960 7358
rect 2024 7294 2040 7358
rect 2104 7294 2120 7358
rect 2184 7294 2200 7358
rect 2264 7294 2280 7358
rect 2344 7294 2352 7358
rect 1952 6026 2352 7294
rect 1952 5962 1960 6026
rect 2024 5962 2040 6026
rect 2104 5962 2120 6026
rect 2184 5962 2200 6026
rect 2264 5962 2280 6026
rect 2344 5962 2352 6026
rect 1952 4694 2352 5962
rect 1952 4630 1960 4694
rect 2024 4630 2040 4694
rect 2104 4630 2120 4694
rect 2184 4630 2200 4694
rect 2264 4630 2280 4694
rect 2344 4630 2352 4694
rect 1952 3362 2352 4630
rect 1952 3298 1960 3362
rect 2024 3298 2040 3362
rect 2104 3298 2120 3362
rect 2184 3298 2200 3362
rect 2264 3298 2280 3362
rect 2344 3298 2352 3362
rect 1952 2616 2352 3298
rect 4952 25340 5352 26022
rect 4952 25276 4960 25340
rect 5024 25276 5040 25340
rect 5104 25276 5120 25340
rect 5184 25276 5200 25340
rect 5264 25276 5280 25340
rect 5344 25276 5352 25340
rect 4952 24008 5352 25276
rect 4952 23944 4960 24008
rect 5024 23944 5040 24008
rect 5104 23944 5120 24008
rect 5184 23944 5200 24008
rect 5264 23944 5280 24008
rect 5344 23944 5352 24008
rect 4952 22676 5352 23944
rect 4952 22612 4960 22676
rect 5024 22612 5040 22676
rect 5104 22612 5120 22676
rect 5184 22612 5200 22676
rect 5264 22612 5280 22676
rect 5344 22612 5352 22676
rect 4952 21344 5352 22612
rect 4952 21280 4960 21344
rect 5024 21280 5040 21344
rect 5104 21280 5120 21344
rect 5184 21280 5200 21344
rect 5264 21280 5280 21344
rect 5344 21280 5352 21344
rect 4952 20012 5352 21280
rect 4952 19948 4960 20012
rect 5024 19948 5040 20012
rect 5104 19948 5120 20012
rect 5184 19948 5200 20012
rect 5264 19948 5280 20012
rect 5344 19948 5352 20012
rect 4952 18680 5352 19948
rect 4952 18616 4960 18680
rect 5024 18616 5040 18680
rect 5104 18616 5120 18680
rect 5184 18616 5200 18680
rect 5264 18616 5280 18680
rect 5344 18616 5352 18680
rect 4952 17348 5352 18616
rect 4952 17284 4960 17348
rect 5024 17284 5040 17348
rect 5104 17284 5120 17348
rect 5184 17284 5200 17348
rect 5264 17284 5280 17348
rect 5344 17284 5352 17348
rect 4952 16016 5352 17284
rect 4952 15952 4960 16016
rect 5024 15952 5040 16016
rect 5104 15952 5120 16016
rect 5184 15952 5200 16016
rect 5264 15952 5280 16016
rect 5344 15952 5352 16016
rect 4952 14684 5352 15952
rect 4952 14620 4960 14684
rect 5024 14620 5040 14684
rect 5104 14620 5120 14684
rect 5184 14620 5200 14684
rect 5264 14620 5280 14684
rect 5344 14620 5352 14684
rect 4952 13352 5352 14620
rect 4952 13288 4960 13352
rect 5024 13288 5040 13352
rect 5104 13288 5120 13352
rect 5184 13288 5200 13352
rect 5264 13288 5280 13352
rect 5344 13288 5352 13352
rect 4952 12020 5352 13288
rect 4952 11956 4960 12020
rect 5024 11956 5040 12020
rect 5104 11956 5120 12020
rect 5184 11956 5200 12020
rect 5264 11956 5280 12020
rect 5344 11956 5352 12020
rect 4952 10688 5352 11956
rect 4952 10624 4960 10688
rect 5024 10624 5040 10688
rect 5104 10624 5120 10688
rect 5184 10624 5200 10688
rect 5264 10624 5280 10688
rect 5344 10624 5352 10688
rect 4952 9356 5352 10624
rect 4952 9292 4960 9356
rect 5024 9292 5040 9356
rect 5104 9292 5120 9356
rect 5184 9292 5200 9356
rect 5264 9292 5280 9356
rect 5344 9292 5352 9356
rect 4952 8024 5352 9292
rect 4952 7960 4960 8024
rect 5024 7960 5040 8024
rect 5104 7960 5120 8024
rect 5184 7960 5200 8024
rect 5264 7960 5280 8024
rect 5344 7960 5352 8024
rect 4952 6692 5352 7960
rect 4952 6628 4960 6692
rect 5024 6628 5040 6692
rect 5104 6628 5120 6692
rect 5184 6628 5200 6692
rect 5264 6628 5280 6692
rect 5344 6628 5352 6692
rect 4952 5360 5352 6628
rect 4952 5296 4960 5360
rect 5024 5296 5040 5360
rect 5104 5296 5120 5360
rect 5184 5296 5200 5360
rect 5264 5296 5280 5360
rect 5344 5296 5352 5360
rect 4952 4028 5352 5296
rect 4952 3964 4960 4028
rect 5024 3964 5040 4028
rect 5104 3964 5120 4028
rect 5184 3964 5200 4028
rect 5264 3964 5280 4028
rect 5344 3964 5352 4028
rect 4952 2696 5352 3964
rect 4952 2632 4960 2696
rect 5024 2632 5040 2696
rect 5104 2632 5120 2696
rect 5184 2632 5200 2696
rect 5264 2632 5280 2696
rect 5344 2632 5352 2696
rect 4952 2616 5352 2632
rect 7952 26006 8352 26022
rect 7952 25942 7960 26006
rect 8024 25942 8040 26006
rect 8104 25942 8120 26006
rect 8184 25942 8200 26006
rect 8264 25942 8280 26006
rect 8344 25942 8352 26006
rect 7952 24674 8352 25942
rect 7952 24610 7960 24674
rect 8024 24610 8040 24674
rect 8104 24610 8120 24674
rect 8184 24610 8200 24674
rect 8264 24610 8280 24674
rect 8344 24610 8352 24674
rect 7952 23342 8352 24610
rect 7952 23278 7960 23342
rect 8024 23278 8040 23342
rect 8104 23278 8120 23342
rect 8184 23278 8200 23342
rect 8264 23278 8280 23342
rect 8344 23278 8352 23342
rect 7952 22010 8352 23278
rect 7952 21946 7960 22010
rect 8024 21946 8040 22010
rect 8104 21946 8120 22010
rect 8184 21946 8200 22010
rect 8264 21946 8280 22010
rect 8344 21946 8352 22010
rect 7952 20678 8352 21946
rect 7952 20614 7960 20678
rect 8024 20614 8040 20678
rect 8104 20614 8120 20678
rect 8184 20614 8200 20678
rect 8264 20614 8280 20678
rect 8344 20614 8352 20678
rect 7952 19346 8352 20614
rect 7952 19282 7960 19346
rect 8024 19282 8040 19346
rect 8104 19282 8120 19346
rect 8184 19282 8200 19346
rect 8264 19282 8280 19346
rect 8344 19282 8352 19346
rect 7952 18014 8352 19282
rect 7952 17950 7960 18014
rect 8024 17950 8040 18014
rect 8104 17950 8120 18014
rect 8184 17950 8200 18014
rect 8264 17950 8280 18014
rect 8344 17950 8352 18014
rect 7952 16682 8352 17950
rect 7952 16618 7960 16682
rect 8024 16618 8040 16682
rect 8104 16618 8120 16682
rect 8184 16618 8200 16682
rect 8264 16618 8280 16682
rect 8344 16618 8352 16682
rect 7952 15350 8352 16618
rect 7952 15286 7960 15350
rect 8024 15286 8040 15350
rect 8104 15286 8120 15350
rect 8184 15286 8200 15350
rect 8264 15286 8280 15350
rect 8344 15286 8352 15350
rect 7952 14018 8352 15286
rect 7952 13954 7960 14018
rect 8024 13954 8040 14018
rect 8104 13954 8120 14018
rect 8184 13954 8200 14018
rect 8264 13954 8280 14018
rect 8344 13954 8352 14018
rect 7952 12686 8352 13954
rect 7952 12622 7960 12686
rect 8024 12622 8040 12686
rect 8104 12622 8120 12686
rect 8184 12622 8200 12686
rect 8264 12622 8280 12686
rect 8344 12622 8352 12686
rect 7952 11354 8352 12622
rect 7952 11290 7960 11354
rect 8024 11290 8040 11354
rect 8104 11290 8120 11354
rect 8184 11290 8200 11354
rect 8264 11290 8280 11354
rect 8344 11290 8352 11354
rect 7952 10022 8352 11290
rect 7952 9958 7960 10022
rect 8024 9958 8040 10022
rect 8104 9958 8120 10022
rect 8184 9958 8200 10022
rect 8264 9958 8280 10022
rect 8344 9958 8352 10022
rect 7952 8690 8352 9958
rect 7952 8626 7960 8690
rect 8024 8626 8040 8690
rect 8104 8626 8120 8690
rect 8184 8626 8200 8690
rect 8264 8626 8280 8690
rect 8344 8626 8352 8690
rect 7952 7358 8352 8626
rect 7952 7294 7960 7358
rect 8024 7294 8040 7358
rect 8104 7294 8120 7358
rect 8184 7294 8200 7358
rect 8264 7294 8280 7358
rect 8344 7294 8352 7358
rect 7952 6026 8352 7294
rect 7952 5962 7960 6026
rect 8024 5962 8040 6026
rect 8104 5962 8120 6026
rect 8184 5962 8200 6026
rect 8264 5962 8280 6026
rect 8344 5962 8352 6026
rect 7952 4694 8352 5962
rect 7952 4630 7960 4694
rect 8024 4630 8040 4694
rect 8104 4630 8120 4694
rect 8184 4630 8200 4694
rect 8264 4630 8280 4694
rect 8344 4630 8352 4694
rect 7952 3362 8352 4630
rect 7952 3298 7960 3362
rect 8024 3298 8040 3362
rect 8104 3298 8120 3362
rect 8184 3298 8200 3362
rect 8264 3298 8280 3362
rect 8344 3298 8352 3362
rect 7952 2616 8352 3298
use sky130_fd_sc_hs__and2_1  _18_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749223325
transform 1 0 8064 0 1 22644
box -38 -49 518 715
use sky130_fd_sc_hs__clkbuf_1  _19_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 9024 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__or4bb_1  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 4800 0 1 6660
box -38 -49 998 715
use sky130_fd_sc_hs__nand2_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749010377
transform 1 0 5568 0 -1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__or3b_1  _22_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 4512 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__o21a_1  _23_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 2400 0 -1 7992
box -38 -49 614 715
use sky130_fd_sc_hs__and2_1  _24_
timestamp 1749223325
transform 1 0 1920 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__a21bo_1  _25_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 3744 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__clkbuf_1  _26_
timestamp 1704896540
transform 1 0 1536 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__nor2_1  _27_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 5472 0 1 6660
box -38 -49 326 715
use sky130_fd_sc_hs__xor2_1  _28_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 5472 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__and2_1  _29_
timestamp 1749223325
transform -1 0 6912 0 -1 5328
box -38 -49 518 715
use sky130_fd_sc_hs__clkbuf_1  _30_
timestamp 1704896540
transform 1 0 1728 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__and3_1  _31_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 6336 0 1 5328
box -38 -49 614 715
use sky130_fd_sc_hs__a21oi_1  _32_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 6720 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__nor3_1  _33_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 1536 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__xor2_1  _34_
timestamp 1704896540
transform 1 0 4800 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__and2_1  _35_
timestamp 1749223325
transform 1 0 2400 0 -1 6660
box -38 -49 518 715
use sky130_fd_sc_hs__clkbuf_1  _36_
timestamp 1704896540
transform -1 0 5184 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__dfxtp_1  _37_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 1920 0 1 6660
box -38 -49 1670 715
use sky130_fd_sc_hs__dfxtp_4  _38_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 2880 0 -1 6660
box -38 -49 1958 715
use sky130_fd_sc_hs__dfrtp_1  _39_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 1536 0 1 17316
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _40_
timestamp 1704896540
transform 1 0 3840 0 1 17316
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _41_
timestamp 1704896540
transform -1 0 4896 0 -1 18648
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _42_
timestamp 1704896540
transform -1 0 4704 0 -1 11988
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _43_
timestamp 1704896540
transform 1 0 2688 0 -1 13320
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _44_
timestamp 1704896540
transform 1 0 5088 0 1 11988
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _45_
timestamp 1704896540
transform 1 0 6432 0 -1 11988
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _46_
timestamp 1704896540
transform 1 0 6528 0 1 9324
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _47_
timestamp 1704896540
transform 1 0 6624 0 -1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _48_
timestamp 1704896540
transform 1 0 6720 0 1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_2  _49_ $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 6048 0 1 15984
box -38 -49 2342 715
use sky130_fd_sc_hs__dfxtp_1  _50_
timestamp 1704896540
transform -1 0 3840 0 -1 5328
box -38 -49 1670 715
use sky130_fd_sc_hs__dfxtp_1  _51_
timestamp 1704896540
transform 1 0 3840 0 -1 3996
box -38 -49 1670 715
use sky130_fd_sc_hs__dfxtp_1  _52_
timestamp 1704896540
transform 1 0 3840 0 -1 5328
box -38 -49 1670 715
use sky130_fd_sc_hs__dfxtp_1  _53_
timestamp 1704896540
transform 1 0 2112 0 1 5328
box -38 -49 1670 715
use sky130_fd_sc_hs__dfrtp_1  _54_
timestamp 1704896540
transform 1 0 4128 0 -1 23976
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _55_
timestamp 1704896540
transform 1 0 5088 0 1 22644
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _56_
timestamp 1704896540
transform 1 0 4896 0 1 21312
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _57_
timestamp 1704896540
transform 1 0 4800 0 1 23976
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _58_
timestamp 1704896540
transform 1 0 3840 0 1 15984
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _59_
timestamp 1704896540
transform 1 0 3744 0 -1 17316
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _60_
timestamp 1704896540
transform 1 0 2208 0 -1 21312
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _61_
timestamp 1704896540
transform -1 0 3744 0 1 22644
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _62_
timestamp 1704896540
transform -1 0 3744 0 1 21312
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _63_
timestamp 1704896540
transform 1 0 2208 0 -1 22644
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _64_
timestamp 1704896540
transform 1 0 7776 0 -1 9324
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _65_
timestamp 1704896540
transform 1 0 7392 0 -1 7992
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _66_
timestamp 1704896540
transform 1 0 6720 0 1 7992
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _67_
timestamp 1704896540
transform 1 0 5952 0 1 6660
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _68_
timestamp 1704896540
transform 1 0 4512 0 1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _69_
timestamp 1704896540
transform 1 0 3360 0 -1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _70_
timestamp 1704896540
transform 1 0 1536 0 1 10656
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _71_
timestamp 1704896540
transform 1 0 1536 0 1 11988
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _72_
timestamp 1704896540
transform -1 0 3744 0 1 15984
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _73_
timestamp 1704896540
transform -1 0 3840 0 -1 15984
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _74_
timestamp 1704896540
transform 1 0 7680 0 -1 23976
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _75_
timestamp 1704896540
transform 1 0 7680 0 -1 22644
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _76_
timestamp 1704896540
transform 1 0 7488 0 -1 18648
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _77_
timestamp 1704896540
transform 1 0 7488 0 -1 15984
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _78_
timestamp 1704896540
transform 1 0 6720 0 1 14652
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _79_
timestamp 1704896540
transform 1 0 7392 0 -1 17316
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _80_
timestamp 1704896540
transform 1 0 7392 0 -1 14652
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _81_
timestamp 1704896540
transform 1 0 6912 0 -1 21312
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _82_
timestamp 1704896540
transform 1 0 6912 0 -1 19980
box -38 -49 2246 715
use sky130_fd_sc_hs__dfrtp_1  _83_
timestamp 1704896540
transform 1 0 6720 0 1 19980
box -38 -49 2246 715
use sky130_fd_sc_hs__clkbuf_16  clkbuf_0_CLK $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 3840 0 1 5328
box -38 -49 1958 715
use sky130_fd_sc_hs__clkbuf_16  clkbuf_1_0__f_CLK
timestamp 1704896540
transform 1 0 4512 0 1 3996
box -38 -49 1958 715
use sky130_fd_sc_hs__clkbuf_16  clkbuf_1_1__f_CLK
timestamp 1704896540
transform -1 0 3744 0 1 7992
box -38 -49 1958 715
use sky130_fd_sc_hs__fill_2  FILLER_0_0_16 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 2688 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_0_18 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 2880 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_0_23 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 3360 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_0_28
timestamp 1704896540
transform 1 0 3840 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_0_30
timestamp 1704896540
transform 1 0 4032 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_0_35 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 4512 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_0_47
timestamp 1704896540
transform 1 0 5664 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_0_51
timestamp 1704896540
transform 1 0 6048 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_0_53
timestamp 1704896540
transform 1 0 6240 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_0_59
timestamp 1704896540
transform 1 0 6816 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_0_71
timestamp 1704896540
transform 1 0 7968 0 1 2664
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_0_79
timestamp 1704896540
transform 1 0 8736 0 1 2664
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_1_4
timestamp 1704896540
transform 1 0 1536 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_1_6
timestamp 1704896540
transform 1 0 1728 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_1_11
timestamp 1704896540
transform 1 0 2208 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_1_19
timestamp 1704896540
transform 1 0 2976 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3744 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_1_45
timestamp 1704896540
transform 1 0 5472 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_1_53
timestamp 1704896540
transform 1 0 6240 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_1_55
timestamp 1704896540
transform 1 0 6432 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_1_63
timestamp 1704896540
transform 1 0 7200 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_1_71
timestamp 1704896540
transform 1 0 7968 0 -1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_1_79
timestamp 1704896540
transform 1 0 8736 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_1_83
timestamp 1704896540
transform 1 0 9120 0 -1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_1_85
timestamp 1704896540
transform 1 0 9312 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_2_8
timestamp 1704896540
transform 1 0 1920 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_2_16
timestamp 1704896540
transform 1 0 2688 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_2_24
timestamp 1704896540
transform 1 0 3456 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_2_26
timestamp 1704896540
transform 1 0 3648 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_2_28
timestamp 1704896540
transform 1 0 3840 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_2_32
timestamp 1704896540
transform 1 0 4224 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_2_34
timestamp 1704896540
transform 1 0 4416 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_2_55
timestamp 1704896540
transform 1 0 6432 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_2_63
timestamp 1704896540
transform 1 0 7200 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_2_71
timestamp 1704896540
transform 1 0 7968 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_2_79
timestamp 1704896540
transform 1 0 8736 0 1 3996
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_2_82
timestamp 1704896540
transform 1 0 9024 0 1 3996
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_2_90
timestamp 1704896540
transform 1 0 9792 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  FILLER_0_3_4
timestamp 1704896540
transform 1 0 1536 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_3_8
timestamp 1704896540
transform 1 0 1920 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_3_10
timestamp 1704896540
transform 1 0 2112 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_3_53
timestamp 1704896540
transform 1 0 6240 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_3_60
timestamp 1704896540
transform 1 0 6912 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_3_68
timestamp 1704896540
transform 1 0 7680 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_3_76
timestamp 1704896540
transform 1 0 8448 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_3_84
timestamp 1704896540
transform 1 0 9216 0 -1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_3_92
timestamp 1704896540
transform 1 0 9984 0 -1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_4_4
timestamp 1704896540
transform 1 0 1536 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_4_58
timestamp 1704896540
transform 1 0 6720 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_4_66
timestamp 1704896540
transform 1 0 7488 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_4_74
timestamp 1704896540
transform 1 0 8256 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_4_78
timestamp 1704896540
transform 1 0 8640 0 1 5328
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_4_80
timestamp 1704896540
transform 1 0 8832 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_4_82
timestamp 1704896540
transform 1 0 9024 0 1 5328
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_4_90
timestamp 1704896540
transform 1 0 9792 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  FILLER_0_5_49
timestamp 1704896540
transform 1 0 5856 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_5_53
timestamp 1704896540
transform 1 0 6240 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_5_55
timestamp 1704896540
transform 1 0 6432 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_5_63
timestamp 1704896540
transform 1 0 7200 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_5_71
timestamp 1704896540
transform 1 0 7968 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_5_79
timestamp 1704896540
transform 1 0 8736 0 -1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_5_87
timestamp 1704896540
transform 1 0 9504 0 -1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_5_89
timestamp 1704896540
transform 1 0 9696 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_6_25
timestamp 1704896540
transform 1 0 3552 0 1 6660
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_6_45
timestamp 1704896540
transform 1 0 5472 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_6_49
timestamp 1704896540
transform 1 0 5856 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_6_73
timestamp 1704896540
transform 1 0 8160 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_6_82
timestamp 1704896540
transform 1 0 9024 0 1 6660
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_6_90
timestamp 1704896540
transform 1 0 9792 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_7_4
timestamp 1704896540
transform 1 0 1536 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_7_12
timestamp 1704896540
transform 1 0 2304 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_7_35
timestamp 1704896540
transform 1 0 4512 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_7_43
timestamp 1704896540
transform 1 0 5280 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_7_51
timestamp 1704896540
transform 1 0 6048 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_7_53
timestamp 1704896540
transform 1 0 6240 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6432 0 -1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_7_63
timestamp 1704896540
transform 1 0 7200 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_7_88
timestamp 1704896540
transform 1 0 9600 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_7_92
timestamp 1704896540
transform 1 0 9984 0 -1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_8_4
timestamp 1704896540
transform 1 0 1536 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_8_6
timestamp 1704896540
transform 1 0 1728 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_8_28
timestamp 1704896540
transform 1 0 3840 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_8_36
timestamp 1704896540
transform 1 0 4608 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_8_44
timestamp 1704896540
transform 1 0 5376 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_8_52
timestamp 1704896540
transform 1 0 6144 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_8_56
timestamp 1704896540
transform 1 0 6528 0 1 7992
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_8_82
timestamp 1704896540
transform 1 0 9024 0 1 7992
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_9_4
timestamp 1704896540
transform 1 0 1536 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_9_12
timestamp 1704896540
transform 1 0 2304 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_9_20
timestamp 1704896540
transform 1 0 3072 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_9_28
timestamp 1704896540
transform 1 0 3840 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_9_36
timestamp 1704896540
transform 1 0 4608 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_9_44
timestamp 1704896540
transform 1 0 5376 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_9_52
timestamp 1704896540
transform 1 0 6144 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_9_55
timestamp 1704896540
transform 1 0 6432 0 -1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_9_63
timestamp 1704896540
transform 1 0 7200 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_9_67
timestamp 1704896540
transform 1 0 7584 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_9_92
timestamp 1704896540
transform 1 0 9984 0 -1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_4
timestamp 1704896540
transform 1 0 1536 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_12
timestamp 1704896540
transform 1 0 2304 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_10_20
timestamp 1704896540
transform 1 0 3072 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_10_24
timestamp 1704896540
transform 1 0 3456 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_10_26
timestamp 1704896540
transform 1 0 3648 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_28
timestamp 1704896540
transform 1 0 3840 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_36
timestamp 1704896540
transform 1 0 4608 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_44
timestamp 1704896540
transform 1 0 5376 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_10_52
timestamp 1704896540
transform 1 0 6144 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_10_79
timestamp 1704896540
transform 1 0 8736 0 1 9324
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_10_82
timestamp 1704896540
transform 1 0 9024 0 1 9324
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_10_90
timestamp 1704896540
transform 1 0 9792 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_11_10
timestamp 1704896540
transform 1 0 2112 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_11_18
timestamp 1704896540
transform 1 0 2880 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_11_22
timestamp 1704896540
transform 1 0 3264 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_11_46
timestamp 1704896540
transform 1 0 5568 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_11_55
timestamp 1704896540
transform 1 0 6432 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_11_80
timestamp 1704896540
transform 1 0 8832 0 -1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_11_88
timestamp 1704896540
transform 1 0 9600 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_11_92
timestamp 1704896540
transform 1 0 9984 0 -1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_12_28
timestamp 1704896540
transform 1 0 3840 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_12_32
timestamp 1704896540
transform 1 0 4224 0 1 10656
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_12_34
timestamp 1704896540
transform 1 0 4416 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_12_82
timestamp 1704896540
transform 1 0 9024 0 1 10656
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_4
timestamp 1704896540
transform 1 0 1536 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_13_12
timestamp 1704896540
transform 1 0 2304 0 -1 11988
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_37
timestamp 1704896540
transform 1 0 4704 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_45
timestamp 1704896540
transform 1 0 5472 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_13_53
timestamp 1704896540
transform 1 0 6240 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_78
timestamp 1704896540
transform 1 0 8640 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_13_86
timestamp 1704896540
transform 1 0 9408 0 -1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_14_28
timestamp 1704896540
transform 1 0 3840 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_14_36
timestamp 1704896540
transform 1 0 4608 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_14_40
timestamp 1704896540
transform 1 0 4992 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_14_64
timestamp 1704896540
transform 1 0 7296 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_14_72
timestamp 1704896540
transform 1 0 8064 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__fill_1  FILLER_0_14_80
timestamp 1704896540
transform 1 0 8832 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_14_82
timestamp 1704896540
transform 1 0 9024 0 1 11988
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_14_90
timestamp 1704896540
transform 1 0 9792 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_15_4
timestamp 1704896540
transform 1 0 1536 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_15_12
timestamp 1704896540
transform 1 0 2304 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_15_39
timestamp 1704896540
transform 1 0 4896 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_15_47
timestamp 1704896540
transform 1 0 5664 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_15_51
timestamp 1704896540
transform 1 0 6048 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_15_53
timestamp 1704896540
transform 1 0 6240 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_15_55
timestamp 1704896540
transform 1 0 6432 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_15_63
timestamp 1704896540
transform 1 0 7200 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_15_71
timestamp 1704896540
transform 1 0 7968 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_15_79
timestamp 1704896540
transform 1 0 8736 0 -1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_15_87
timestamp 1704896540
transform 1 0 9504 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_15_91
timestamp 1704896540
transform 1 0 9888 0 -1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_15_93
timestamp 1704896540
transform 1 0 10080 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_4
timestamp 1704896540
transform 1 0 1536 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_12
timestamp 1704896540
transform 1 0 2304 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_16_20
timestamp 1704896540
transform 1 0 3072 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_16_24
timestamp 1704896540
transform 1 0 3456 0 1 13320
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_16_26
timestamp 1704896540
transform 1 0 3648 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_28
timestamp 1704896540
transform 1 0 3840 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_36
timestamp 1704896540
transform 1 0 4608 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_44
timestamp 1704896540
transform 1 0 5376 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_52
timestamp 1704896540
transform 1 0 6144 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_60
timestamp 1704896540
transform 1 0 6912 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_68
timestamp 1704896540
transform 1 0 7680 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_16_76
timestamp 1704896540
transform 1 0 8448 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_16_80
timestamp 1704896540
transform 1 0 8832 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_16_82
timestamp 1704896540
transform 1 0 9024 0 1 13320
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_17_8
timestamp 1704896540
transform 1 0 1920 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_17_16
timestamp 1704896540
transform 1 0 2688 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_17_24
timestamp 1704896540
transform 1 0 3456 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_17_32
timestamp 1704896540
transform 1 0 4224 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_17_40
timestamp 1704896540
transform 1 0 4992 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_17_48
timestamp 1704896540
transform 1 0 5760 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_17_52
timestamp 1704896540
transform 1 0 6144 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_17_55
timestamp 1704896540
transform 1 0 6432 0 -1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_17_63
timestamp 1704896540
transform 1 0 7200 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_17_88
timestamp 1704896540
transform 1 0 9600 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_17_92
timestamp 1704896540
transform 1 0 9984 0 -1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_18_4
timestamp 1704896540
transform 1 0 1536 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_18_12
timestamp 1704896540
transform 1 0 2304 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_18_20
timestamp 1704896540
transform 1 0 3072 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_18_24
timestamp 1704896540
transform 1 0 3456 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_18_26
timestamp 1704896540
transform 1 0 3648 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_18_28
timestamp 1704896540
transform 1 0 3840 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_18_36
timestamp 1704896540
transform 1 0 4608 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_18_44
timestamp 1704896540
transform 1 0 5376 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_18_52
timestamp 1704896540
transform 1 0 6144 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_18_56
timestamp 1704896540
transform 1 0 6528 0 1 14652
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_18_82
timestamp 1704896540
transform 1 0 9024 0 1 14652
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_18_90
timestamp 1704896540
transform 1 0 9792 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_19_4
timestamp 1704896540
transform 1 0 1536 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_19_28
timestamp 1704896540
transform 1 0 3840 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_19_36
timestamp 1704896540
transform 1 0 4608 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_19_44
timestamp 1704896540
transform 1 0 5376 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_19_52
timestamp 1704896540
transform 1 0 6144 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_19_55
timestamp 1704896540
transform 1 0 6432 0 -1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_19_63
timestamp 1704896540
transform 1 0 7200 0 -1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_19_65
timestamp 1704896540
transform 1 0 7392 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_19_89
timestamp 1704896540
transform 1 0 9696 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_20_75
timestamp 1704896540
transform 1 0 8352 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_20_79
timestamp 1704896540
transform 1 0 8736 0 1 15984
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_20_82
timestamp 1704896540
transform 1 0 9024 0 1 15984
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_20_90
timestamp 1704896540
transform 1 0 9792 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_21_4
timestamp 1704896540
transform 1 0 1536 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_21_12
timestamp 1704896540
transform 1 0 2304 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_21_20
timestamp 1704896540
transform 1 0 3072 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_21_24
timestamp 1704896540
transform 1 0 3456 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_21_26
timestamp 1704896540
transform 1 0 3648 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__decap_4  FILLER_0_21_50
timestamp 1704896540
transform 1 0 5952 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_21_55
timestamp 1704896540
transform 1 0 6432 0 -1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_21_63
timestamp 1704896540
transform 1 0 7200 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_21_88
timestamp 1704896540
transform 1 0 9600 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_21_92
timestamp 1704896540
transform 1 0 9984 0 -1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_22_51
timestamp 1704896540
transform 1 0 6048 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_22_59
timestamp 1704896540
transform 1 0 6816 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_22_67
timestamp 1704896540
transform 1 0 7584 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_22_75
timestamp 1704896540
transform 1 0 8352 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_22_79
timestamp 1704896540
transform 1 0 8736 0 1 17316
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_22_82
timestamp 1704896540
transform 1 0 9024 0 1 17316
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_22_90
timestamp 1704896540
transform 1 0 9792 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_23_4
timestamp 1704896540
transform 1 0 1536 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_23_12
timestamp 1704896540
transform 1 0 2304 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_23_39
timestamp 1704896540
transform 1 0 4896 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_23_47
timestamp 1704896540
transform 1 0 5664 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_23_51
timestamp 1704896540
transform 1 0 6048 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_23_53
timestamp 1704896540
transform 1 0 6240 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_23_55
timestamp 1704896540
transform 1 0 6432 0 -1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_23_63
timestamp 1704896540
transform 1 0 7200 0 -1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_23_65
timestamp 1704896540
transform 1 0 7392 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_1  FILLER_0_23_89
timestamp 1704896540
transform 1 0 9696 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_24_8
timestamp 1704896540
transform 1 0 1920 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_24_16
timestamp 1704896540
transform 1 0 2688 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_24_24
timestamp 1704896540
transform 1 0 3456 0 1 18648
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_24_26
timestamp 1704896540
transform 1 0 3648 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_24_28
timestamp 1704896540
transform 1 0 3840 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_24_36
timestamp 1704896540
transform 1 0 4608 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_24_44
timestamp 1704896540
transform 1 0 5376 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_24_52
timestamp 1704896540
transform 1 0 6144 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_24_60
timestamp 1704896540
transform 1 0 6912 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_24_68
timestamp 1704896540
transform 1 0 7680 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_24_76
timestamp 1704896540
transform 1 0 8448 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_24_80
timestamp 1704896540
transform 1 0 8832 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_24_82
timestamp 1704896540
transform 1 0 9024 0 1 18648
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_24_90
timestamp 1704896540
transform 1 0 9792 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_25_4
timestamp 1704896540
transform 1 0 1536 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_25_12
timestamp 1704896540
transform 1 0 2304 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_25_20
timestamp 1704896540
transform 1 0 3072 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_25_28
timestamp 1704896540
transform 1 0 3840 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_25_36
timestamp 1704896540
transform 1 0 4608 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_25_44
timestamp 1704896540
transform 1 0 5376 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_25_52
timestamp 1704896540
transform 1 0 6144 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__decap_4  FILLER_0_25_55
timestamp 1704896540
transform 1 0 6432 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_25_59
timestamp 1704896540
transform 1 0 6816 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_25_83
timestamp 1704896540
transform 1 0 9120 0 -1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_25_91
timestamp 1704896540
transform 1 0 9888 0 -1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_25_93
timestamp 1704896540
transform 1 0 10080 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_26_4
timestamp 1704896540
transform 1 0 1536 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_26_12
timestamp 1704896540
transform 1 0 2304 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_26_20
timestamp 1704896540
transform 1 0 3072 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_26_24
timestamp 1704896540
transform 1 0 3456 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_26_26
timestamp 1704896540
transform 1 0 3648 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_26_28
timestamp 1704896540
transform 1 0 3840 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_26_36
timestamp 1704896540
transform 1 0 4608 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_26_44
timestamp 1704896540
transform 1 0 5376 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_26_52
timestamp 1704896540
transform 1 0 6144 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_26_56
timestamp 1704896540
transform 1 0 6528 0 1 19980
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_26_82
timestamp 1704896540
transform 1 0 9024 0 1 19980
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_27_4
timestamp 1704896540
transform 1 0 1536 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_27_8
timestamp 1704896540
transform 1 0 1920 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_27_10
timestamp 1704896540
transform 1 0 2112 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_27_34
timestamp 1704896540
transform 1 0 4416 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_27_42
timestamp 1704896540
transform 1 0 5184 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_27_50
timestamp 1704896540
transform 1 0 5952 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  FILLER_0_27_55
timestamp 1704896540
transform 1 0 6432 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_27_59
timestamp 1704896540
transform 1 0 6816 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_27_83
timestamp 1704896540
transform 1 0 9120 0 -1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_27_91
timestamp 1704896540
transform 1 0 9888 0 -1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_27_93
timestamp 1704896540
transform 1 0 10080 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_28_28
timestamp 1704896540
transform 1 0 3840 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_28_36
timestamp 1704896540
transform 1 0 4608 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_28_38
timestamp 1704896540
transform 1 0 4800 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_28_62
timestamp 1704896540
transform 1 0 7104 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_28_70
timestamp 1704896540
transform 1 0 7872 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_28_78
timestamp 1704896540
transform 1 0 8640 0 1 21312
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_28_80
timestamp 1704896540
transform 1 0 8832 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_28_82
timestamp 1704896540
transform 1 0 9024 0 1 21312
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_28_90
timestamp 1704896540
transform 1 0 9792 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__fill_2  FILLER_0_29_8
timestamp 1704896540
transform 1 0 1920 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_29_10
timestamp 1704896540
transform 1 0 2112 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_29_34
timestamp 1704896540
transform 1 0 4416 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_29_42
timestamp 1704896540
transform 1 0 5184 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_29_50
timestamp 1704896540
transform 1 0 5952 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_29_55
timestamp 1704896540
transform 1 0 6432 0 -1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_29_63
timestamp 1704896540
transform 1 0 7200 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_29_67
timestamp 1704896540
transform 1 0 7584 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_29_91
timestamp 1704896540
transform 1 0 9888 0 -1 22644
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_29_93
timestamp 1704896540
transform 1 0 10080 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_30_28
timestamp 1704896540
transform 1 0 3840 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_30_36
timestamp 1704896540
transform 1 0 4608 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_30_40
timestamp 1704896540
transform 1 0 4992 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_30_64
timestamp 1704896540
transform 1 0 7296 0 1 22644
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_30_77
timestamp 1704896540
transform 1 0 8544 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  FILLER_0_30_86
timestamp 1704896540
transform 1 0 9408 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_31_4
timestamp 1704896540
transform 1 0 1536 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_31_12
timestamp 1704896540
transform 1 0 2304 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_31_20
timestamp 1704896540
transform 1 0 3072 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_31_28
timestamp 1704896540
transform 1 0 3840 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_31_30
timestamp 1704896540
transform 1 0 4032 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_31_55
timestamp 1704896540
transform 1 0 6432 0 -1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_31_63
timestamp 1704896540
transform 1 0 7200 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__fill_1  FILLER_0_31_67
timestamp 1704896540
transform 1 0 7584 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_31_91
timestamp 1704896540
transform 1 0 9888 0 -1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_31_93
timestamp 1704896540
transform 1 0 10080 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_8
timestamp 1704896540
transform 1 0 1920 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_16
timestamp 1704896540
transform 1 0 2688 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_32_24
timestamp 1704896540
transform 1 0 3456 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_32_26
timestamp 1704896540
transform 1 0 3648 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_28
timestamp 1704896540
transform 1 0 3840 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_32_36
timestamp 1704896540
transform 1 0 4608 0 1 23976
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_61
timestamp 1704896540
transform 1 0 7008 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_69
timestamp 1704896540
transform 1 0 7776 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__decap_4  FILLER_0_32_77
timestamp 1704896540
transform 1 0 8544 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__fill_8  FILLER_0_32_82
timestamp 1704896540
transform 1 0 9024 0 1 23976
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_12
timestamp 1704896540
transform 1 0 2304 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_20
timestamp 1704896540
transform 1 0 3072 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_28
timestamp 1704896540
transform 1 0 3840 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_36
timestamp 1704896540
transform 1 0 4608 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_44
timestamp 1704896540
transform 1 0 5376 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_33_52
timestamp 1704896540
transform 1 0 6144 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_55
timestamp 1704896540
transform 1 0 6432 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_63
timestamp 1704896540
transform 1 0 7200 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_8  FILLER_0_33_71
timestamp 1704896540
transform 1 0 7968 0 -1 25308
box -38 -49 806 715
use sky130_fd_sc_hs__fill_2  FILLER_0_33_79
timestamp 1704896540
transform 1 0 8736 0 -1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_33_81
timestamp 1704896540
transform 1 0 8928 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_8
timestamp 1704896540
transform 1 0 1920 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_14
timestamp 1704896540
transform 1 0 2496 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_20
timestamp 1704896540
transform 1 0 3072 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_34_26
timestamp 1704896540
transform 1 0 3648 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_32
timestamp 1704896540
transform 1 0 4224 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_38
timestamp 1704896540
transform 1 0 4800 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_44
timestamp 1704896540
transform 1 0 5376 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_55
timestamp 1704896540
transform 1 0 6432 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_34_57
timestamp 1704896540
transform 1 0 6624 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_62
timestamp 1704896540
transform 1 0 7104 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_68
timestamp 1704896540
transform 1 0 7680 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_74
timestamp 1704896540
transform 1 0 8256 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_1  FILLER_0_34_80
timestamp 1704896540
transform 1 0 8832 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_86
timestamp 1704896540
transform 1 0 9408 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__fill_2  FILLER_0_34_92
timestamp 1704896540
transform 1 0 9984 0 1 25308
box -38 -49 230 715
use sky130_fd_sc_hs__clkbuf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 1920 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_2  input2
timestamp 1704896540
transform -1 0 1920 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__buf_8  input3 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform 1 0 1536 0 1 2664
box -38 -49 1190 715
use sky130_fd_sc_hs__clkbuf_4  input4 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 2112 0 -1 10656
box -38 -49 614 715
use sky130_fd_sc_hs__clkbuf_1  output5
timestamp 1704896540
transform 1 0 5952 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output6
timestamp 1704896540
transform -1 0 7104 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output7
timestamp 1704896540
transform -1 0 7680 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output8
timestamp 1704896540
transform -1 0 8256 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output9
timestamp 1704896540
transform -1 0 8832 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output10
timestamp 1704896540
transform -1 0 9408 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output11
timestamp 1704896540
transform -1 0 9984 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output12
timestamp 1704896540
transform 1 0 9792 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output13
timestamp 1704896540
transform 1 0 9408 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output14
timestamp 1704896540
transform 1 0 9792 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output15
timestamp 1704896540
transform 1 0 9024 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output16
timestamp 1704896540
transform -1 0 1920 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output17
timestamp 1704896540
transform -1 0 1920 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output18
timestamp 1704896540
transform 1 0 9408 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output19
timestamp 1704896540
transform 1 0 9792 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output20
timestamp 1704896540
transform 1 0 9792 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output21
timestamp 1704896540
transform 1 0 9792 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output22
timestamp 1704896540
transform 1 0 9792 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output23
timestamp 1704896540
transform 1 0 9792 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output24
timestamp 1704896540
transform 1 0 9792 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output25
timestamp 1704896540
transform 1 0 9792 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output26
timestamp 1704896540
transform 1 0 9792 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output27
timestamp 1704896540
transform 1 0 9792 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output28
timestamp 1704896540
transform -1 0 1920 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output29
timestamp 1704896540
transform -1 0 2208 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output30
timestamp 1704896540
transform -1 0 3360 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output31
timestamp 1704896540
transform -1 0 4512 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output32
timestamp 1704896540
transform -1 0 5664 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output33
timestamp 1704896540
transform -1 0 6816 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output34
timestamp 1704896540
transform -1 0 7968 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output35
timestamp 1704896540
transform -1 0 9408 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output36
timestamp 1704896540
transform -1 0 10176 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output37
timestamp 1704896540
transform 1 0 9408 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output38
timestamp 1704896540
transform -1 0 2304 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output39
timestamp 1704896540
transform -1 0 1920 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output40
timestamp 1704896540
transform -1 0 1920 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output41
timestamp 1704896540
transform -1 0 2496 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output42
timestamp 1704896540
transform -1 0 3072 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output43
timestamp 1704896540
transform -1 0 3648 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output44
timestamp 1704896540
transform -1 0 4224 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output45
timestamp 1704896540
transform -1 0 4800 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output46
timestamp 1704896540
transform -1 0 5376 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__clkbuf_1  output47
timestamp 1704896540
transform -1 0 5952 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_0_Left_35
timestamp 1704896540
transform 1 0 1152 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 10560 0 1 2664
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_1_Left_36
timestamp 1704896540
transform 1 0 1152 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 10560 0 -1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_2_Left_37
timestamp 1704896540
transform 1 0 1152 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 10560 0 1 3996
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_3_Left_38
timestamp 1704896540
transform 1 0 1152 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 10560 0 -1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_4_Left_39
timestamp 1704896540
transform 1 0 1152 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 10560 0 1 5328
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_5_Left_40
timestamp 1704896540
transform 1 0 1152 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 10560 0 -1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_6_Left_41
timestamp 1704896540
transform 1 0 1152 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 10560 0 1 6660
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_7_Left_42
timestamp 1704896540
transform 1 0 1152 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 10560 0 -1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_8_Left_43
timestamp 1704896540
transform 1 0 1152 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 10560 0 1 7992
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_9_Left_44
timestamp 1704896540
transform 1 0 1152 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 10560 0 -1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_10_Left_45
timestamp 1704896540
transform 1 0 1152 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 10560 0 1 9324
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_11_Left_46
timestamp 1704896540
transform 1 0 1152 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 10560 0 -1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_12_Left_47
timestamp 1704896540
transform 1 0 1152 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 10560 0 1 10656
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_13_Left_48
timestamp 1704896540
transform 1 0 1152 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 10560 0 -1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_14_Left_49
timestamp 1704896540
transform 1 0 1152 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 10560 0 1 11988
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_15_Left_50
timestamp 1704896540
transform 1 0 1152 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 10560 0 -1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_16_Left_51
timestamp 1704896540
transform 1 0 1152 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 10560 0 1 13320
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_17_Left_52
timestamp 1704896540
transform 1 0 1152 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 10560 0 -1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_18_Left_53
timestamp 1704896540
transform 1 0 1152 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 10560 0 1 14652
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_19_Left_54
timestamp 1704896540
transform 1 0 1152 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 10560 0 -1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_20_Left_55
timestamp 1704896540
transform 1 0 1152 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 10560 0 1 15984
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_21_Left_56
timestamp 1704896540
transform 1 0 1152 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 10560 0 -1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_22_Left_57
timestamp 1704896540
transform 1 0 1152 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 10560 0 1 17316
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_23_Left_58
timestamp 1704896540
transform 1 0 1152 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 10560 0 -1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_24_Left_59
timestamp 1704896540
transform 1 0 1152 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 10560 0 1 18648
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_25_Left_60
timestamp 1704896540
transform 1 0 1152 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 10560 0 -1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_26_Left_61
timestamp 1704896540
transform 1 0 1152 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 10560 0 1 19980
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_27_Left_62
timestamp 1704896540
transform 1 0 1152 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 10560 0 -1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_28_Left_63
timestamp 1704896540
transform 1 0 1152 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 10560 0 1 21312
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_29_Left_64
timestamp 1704896540
transform 1 0 1152 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_29_Right_29
timestamp 1704896540
transform -1 0 10560 0 -1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_30_Left_65
timestamp 1704896540
transform 1 0 1152 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_30_Right_30
timestamp 1704896540
transform -1 0 10560 0 1 22644
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_31_Left_66
timestamp 1704896540
transform 1 0 1152 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_31_Right_31
timestamp 1704896540
transform -1 0 10560 0 -1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_32_Left_67
timestamp 1704896540
transform 1 0 1152 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_32_Right_32
timestamp 1704896540
transform -1 0 10560 0 1 23976
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_33_Left_68
timestamp 1704896540
transform 1 0 1152 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_33_Right_33
timestamp 1704896540
transform -1 0 10560 0 -1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_34_Left_69
timestamp 1704896540
transform 1 0 1152 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__decap_4  PHY_EDGE_ROW_34_Right_34
timestamp 1704896540
transform -1 0 10560 0 1 25308
box -38 -49 422 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749010377
transform 1 0 3744 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1749010377
transform 1 0 6336 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1749010377
transform 1 0 8928 0 1 2664
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_73
timestamp 1749010377
transform 1 0 6336 0 -1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_74
timestamp 1749010377
transform 1 0 3744 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_75
timestamp 1749010377
transform 1 0 8928 0 1 3996
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_76
timestamp 1749010377
transform 1 0 6336 0 -1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_77
timestamp 1749010377
transform 1 0 3744 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_78
timestamp 1749010377
transform 1 0 8928 0 1 5328
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_79
timestamp 1749010377
transform 1 0 6336 0 -1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_80
timestamp 1749010377
transform 1 0 3744 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_81
timestamp 1749010377
transform 1 0 8928 0 1 6660
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp 1749010377
transform 1 0 6336 0 -1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp 1749010377
transform 1 0 3744 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_84
timestamp 1749010377
transform 1 0 8928 0 1 7992
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_85
timestamp 1749010377
transform 1 0 6336 0 -1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_86
timestamp 1749010377
transform 1 0 3744 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_87
timestamp 1749010377
transform 1 0 8928 0 1 9324
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_88
timestamp 1749010377
transform 1 0 6336 0 -1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_89
timestamp 1749010377
transform 1 0 3744 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_90
timestamp 1749010377
transform 1 0 8928 0 1 10656
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_91
timestamp 1749010377
transform 1 0 6336 0 -1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_92
timestamp 1749010377
transform 1 0 3744 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_93
timestamp 1749010377
transform 1 0 8928 0 1 11988
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_94
timestamp 1749010377
transform 1 0 6336 0 -1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_95
timestamp 1749010377
transform 1 0 3744 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_96
timestamp 1749010377
transform 1 0 8928 0 1 13320
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_97
timestamp 1749010377
transform 1 0 6336 0 -1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_98
timestamp 1749010377
transform 1 0 3744 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_99
timestamp 1749010377
transform 1 0 8928 0 1 14652
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_100
timestamp 1749010377
transform 1 0 6336 0 -1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_101
timestamp 1749010377
transform 1 0 3744 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_102
timestamp 1749010377
transform 1 0 8928 0 1 15984
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_103
timestamp 1749010377
transform 1 0 6336 0 -1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_104
timestamp 1749010377
transform 1 0 3744 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_105
timestamp 1749010377
transform 1 0 8928 0 1 17316
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_106
timestamp 1749010377
transform 1 0 6336 0 -1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_107
timestamp 1749010377
transform 1 0 3744 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_108
timestamp 1749010377
transform 1 0 8928 0 1 18648
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_109
timestamp 1749010377
transform 1 0 6336 0 -1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_110
timestamp 1749010377
transform 1 0 3744 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_111
timestamp 1749010377
transform 1 0 8928 0 1 19980
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_112
timestamp 1749010377
transform 1 0 6336 0 -1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_113
timestamp 1749010377
transform 1 0 3744 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_114
timestamp 1749010377
transform 1 0 8928 0 1 21312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_115
timestamp 1749010377
transform 1 0 6336 0 -1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_116
timestamp 1749010377
transform 1 0 3744 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_117
timestamp 1749010377
transform 1 0 8928 0 1 22644
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_118
timestamp 1749010377
transform 1 0 6336 0 -1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_119
timestamp 1749010377
transform 1 0 3744 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_120
timestamp 1749010377
transform 1 0 8928 0 1 23976
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_121
timestamp 1749010377
transform 1 0 6336 0 -1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_122
timestamp 1749010377
transform 1 0 3744 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_123
timestamp 1749010377
transform 1 0 6336 0 1 25308
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_124
timestamp 1749010377
transform 1 0 8928 0 1 25308
box -38 -49 134 715
<< labels >>
flabel metal2 s 6068 28074 6124 28874 0 FreeSans 224 90 0 0 CF[0]
port 0 nsew signal output
flabel metal2 s 6644 28074 6700 28874 0 FreeSans 224 90 0 0 CF[1]
port 1 nsew signal output
flabel metal2 s 7220 28074 7276 28874 0 FreeSans 224 90 0 0 CF[2]
port 2 nsew signal output
flabel metal2 s 7796 28074 7852 28874 0 FreeSans 224 90 0 0 CF[3]
port 3 nsew signal output
flabel metal2 s 8372 28074 8428 28874 0 FreeSans 224 90 0 0 CF[4]
port 4 nsew signal output
flabel metal2 s 8948 28074 9004 28874 0 FreeSans 224 90 0 0 CF[5]
port 5 nsew signal output
flabel metal2 s 9524 28074 9580 28874 0 FreeSans 224 90 0 0 CF[6]
port 6 nsew signal output
flabel metal2 s 10100 28074 10156 28874 0 FreeSans 224 90 0 0 CF[7]
port 7 nsew signal output
flabel metal2 s 10676 28074 10732 28874 0 FreeSans 224 90 0 0 CF[8]
port 8 nsew signal output
flabel metal2 s 11252 28074 11308 28874 0 FreeSans 224 90 0 0 CF[9]
port 9 nsew signal output
flabel metal3 s 10922 27246 11722 27366 0 FreeSans 480 0 0 0 CKO
port 10 nsew signal output
flabel metal3 s 0 22510 800 22630 0 FreeSans 480 0 0 0 CKS
port 11 nsew signal output
flabel metal3 s 0 26654 800 26774 0 FreeSans 480 0 0 0 CKSB
port 12 nsew signal output
flabel metal3 s 0 5934 800 6054 0 FreeSans 480 0 0 0 CLK
port 13 nsew signal input
flabel metal3 s 0 18366 800 18486 0 FreeSans 480 0 0 0 CMP_N
port 14 nsew signal input
flabel metal3 s 0 14222 800 14342 0 FreeSans 480 0 0 0 CMP_P
port 15 nsew signal input
flabel metal3 s 10922 1198 11722 1318 0 FreeSans 480 0 0 0 DATA[0]
port 16 nsew signal output
flabel metal3 s 10922 3566 11722 3686 0 FreeSans 480 0 0 0 DATA[1]
port 17 nsew signal output
flabel metal3 s 10922 5934 11722 6054 0 FreeSans 480 0 0 0 DATA[2]
port 18 nsew signal output
flabel metal3 s 10922 8302 11722 8422 0 FreeSans 480 0 0 0 DATA[3]
port 19 nsew signal output
flabel metal3 s 10922 10670 11722 10790 0 FreeSans 480 0 0 0 DATA[4]
port 20 nsew signal output
flabel metal3 s 10922 13038 11722 13158 0 FreeSans 480 0 0 0 DATA[5]
port 21 nsew signal output
flabel metal3 s 10922 15406 11722 15526 0 FreeSans 480 0 0 0 DATA[6]
port 22 nsew signal output
flabel metal3 s 10922 17774 11722 17894 0 FreeSans 480 0 0 0 DATA[7]
port 23 nsew signal output
flabel metal3 s 10922 20142 11722 20262 0 FreeSans 480 0 0 0 DATA[8]
port 24 nsew signal output
flabel metal3 s 10922 22510 11722 22630 0 FreeSans 480 0 0 0 DATA[9]
port 25 nsew signal output
flabel metal3 s 0 1790 800 1910 0 FreeSans 480 0 0 0 EN
port 26 nsew signal input
flabel metal3 s 0 10078 800 10198 0 FreeSans 480 0 0 0 RDY
port 27 nsew signal input
flabel metal2 s 596 0 652 800 0 FreeSans 224 90 0 0 SWN[0]
port 28 nsew signal output
flabel metal2 s 1748 0 1804 800 0 FreeSans 224 90 0 0 SWN[1]
port 29 nsew signal output
flabel metal2 s 2900 0 2956 800 0 FreeSans 224 90 0 0 SWN[2]
port 30 nsew signal output
flabel metal2 s 4052 0 4108 800 0 FreeSans 224 90 0 0 SWN[3]
port 31 nsew signal output
flabel metal2 s 5204 0 5260 800 0 FreeSans 224 90 0 0 SWN[4]
port 32 nsew signal output
flabel metal2 s 6356 0 6412 800 0 FreeSans 224 90 0 0 SWN[5]
port 33 nsew signal output
flabel metal2 s 7508 0 7564 800 0 FreeSans 224 90 0 0 SWN[6]
port 34 nsew signal output
flabel metal2 s 8660 0 8716 800 0 FreeSans 224 90 0 0 SWN[7]
port 35 nsew signal output
flabel metal2 s 9812 0 9868 800 0 FreeSans 224 90 0 0 SWN[8]
port 36 nsew signal output
flabel metal2 s 10964 0 11020 800 0 FreeSans 224 90 0 0 SWN[9]
port 37 nsew signal output
flabel metal2 s 308 28074 364 28874 0 FreeSans 224 90 0 0 SWP[0]
port 38 nsew signal output
flabel metal2 s 884 28074 940 28874 0 FreeSans 224 90 0 0 SWP[1]
port 39 nsew signal output
flabel metal2 s 1460 28074 1516 28874 0 FreeSans 224 90 0 0 SWP[2]
port 40 nsew signal output
flabel metal2 s 2036 28074 2092 28874 0 FreeSans 224 90 0 0 SWP[3]
port 41 nsew signal output
flabel metal2 s 2612 28074 2668 28874 0 FreeSans 224 90 0 0 SWP[4]
port 42 nsew signal output
flabel metal2 s 3188 28074 3244 28874 0 FreeSans 224 90 0 0 SWP[5]
port 43 nsew signal output
flabel metal2 s 3764 28074 3820 28874 0 FreeSans 224 90 0 0 SWP[6]
port 44 nsew signal output
flabel metal2 s 4340 28074 4396 28874 0 FreeSans 224 90 0 0 SWP[7]
port 45 nsew signal output
flabel metal2 s 4916 28074 4972 28874 0 FreeSans 224 90 0 0 SWP[8]
port 46 nsew signal output
flabel metal2 s 5492 28074 5548 28874 0 FreeSans 224 90 0 0 SWP[9]
port 47 nsew signal output
flabel metal4 s 4952 2616 5352 26022 0 FreeSans 1920 90 0 0 VGND
port 48 nsew ground bidirectional
flabel metal4 s 1952 2616 2352 26022 0 FreeSans 1920 90 0 0 VPWR
port 49 nsew power bidirectional
flabel metal4 s 7952 2616 8352 26022 0 FreeSans 1920 90 0 0 VPWR
port 49 nsew power bidirectional
rlabel metal1 5856 25308 5856 25308 0 VGND
rlabel metal1 5856 25974 5856 25974 0 VPWR
rlabel metal2 6199 28194 6199 28194 0 CF[0]
rlabel metal2 6727 28194 6727 28194 0 CF[1]
rlabel metal2 7303 28194 7303 28194 0 CF[2]
rlabel metal2 7879 28194 7879 28194 0 CF[3]
rlabel metal2 8455 28194 8455 28194 0 CF[4]
rlabel metal2 9031 28194 9031 28194 0 CF[5]
rlabel metal2 9607 28194 9607 28194 0 CF[6]
rlabel metal2 10128 26688 10128 26688 0 CF[7]
rlabel metal1 10224 25123 10224 25123 0 CF[8]
rlabel metal1 10704 24457 10704 24457 0 CF[9]
rlabel metal2 9360 26251 9360 26251 0 CKO
rlabel metal1 1440 22533 1440 22533 0 CKS
rlabel metal1 1536 25197 1536 25197 0 CKSB
rlabel metal2 3888 5753 3888 5753 0 CLK
rlabel metal3 1191 18426 1191 18426 0 CMP_N
rlabel metal3 807 14282 807 14282 0 CMP_P
rlabel metal2 9744 2090 9744 2090 0 DATA[0]
rlabel via2 10128 3607 10128 3607 0 DATA[1]
rlabel metal2 10128 6049 10128 6049 0 DATA[2]
rlabel via2 10128 8343 10128 8343 0 DATA[3]
rlabel via2 10128 10748 10128 10748 0 DATA[4]
rlabel metal2 10128 13264 10128 13264 0 DATA[5]
rlabel via2 10128 15447 10128 15447 0 DATA[6]
rlabel metal2 10128 17963 10128 17963 0 DATA[7]
rlabel via2 10128 20183 10128 20183 0 DATA[8]
rlabel metal2 10128 22662 10128 22662 0 DATA[9]
rlabel metal3 1143 1850 1143 1850 0 EN
rlabel metal3 807 10138 807 10138 0 RDY
rlabel metal1 1104 4107 1104 4107 0 SWN[0]
rlabel metal2 1831 666 1831 666 0 SWN[1]
rlabel metal2 2928 1801 2928 1801 0 SWN[2]
rlabel metal2 4080 1801 4080 1801 0 SWN[3]
rlabel metal2 5232 1043 5232 1043 0 SWN[4]
rlabel metal2 6384 1801 6384 1801 0 SWN[5]
rlabel metal2 7591 666 7591 666 0 SWN[6]
rlabel metal2 8688 1801 8688 1801 0 SWN[7]
rlabel metal2 9840 1801 9840 1801 0 SWN[8]
rlabel metal2 10992 2060 10992 2060 0 SWN[9]
rlabel metal1 1152 25123 1152 25123 0 SWP[0]
rlabel metal1 1248 24457 1248 24457 0 SWP[1]
rlabel metal2 1543 28194 1543 28194 0 SWP[2]
rlabel metal1 2016 25863 2016 25863 0 SWP[3]
rlabel metal1 2688 25863 2688 25863 0 SWP[4]
rlabel metal2 3271 28194 3271 28194 0 SWP[5]
rlabel metal2 3847 28194 3847 28194 0 SWP[6]
rlabel metal2 4423 28194 4423 28194 0 SWP[7]
rlabel metal2 4999 28194 4999 28194 0 SWP[8]
rlabel metal1 5568 25863 5568 25863 0 SWP[9]
rlabel metal1 2400 7067 2400 7067 0 _00_
rlabel metal2 3312 6586 3312 6586 0 _01_
rlabel metal1 4416 4921 4416 4921 0 _02_
rlabel metal1 3936 3737 3936 3737 0 _03_
rlabel metal2 4272 5587 4272 5587 0 _04_
rlabel metal2 3984 6290 3984 6290 0 _05_
rlabel metal1 8784 22977 8784 22977 0 _06_
rlabel metal2 3888 6475 3888 6475 0 _07_
rlabel metal1 5232 7030 5232 7030 0 _08_
rlabel metal1 3504 7733 3504 7733 0 _09_
rlabel metal1 3312 7881 3312 7881 0 _10_
rlabel metal2 3024 7289 3024 7289 0 _11_
rlabel metal1 6672 5106 6672 5106 0 _12_
rlabel metal2 1776 5254 1776 5254 0 _13_
rlabel via2 5136 6308 5136 6308 0 _14_
rlabel metal2 2448 5994 2448 5994 0 _15_
rlabel metal1 4272 6475 4272 6475 0 _16_
rlabel metal1 5040 6919 5040 6919 0 _17_
rlabel metal1 5808 5069 5808 5069 0 clk_div_0.COUNT\[0\]
rlabel metal2 5520 5587 5520 5587 0 clk_div_0.COUNT\[1\]
rlabel metal1 5088 5217 5088 5217 0 clk_div_0.COUNT\[2\]
rlabel metal2 4848 5920 4848 5920 0 clk_div_0.COUNT\[3\]
rlabel metal2 4560 5032 4560 5032 0 clknet_0_CLK
rlabel metal2 3888 4699 3888 4699 0 clknet_1_0__leaf_CLK
rlabel metal1 1920 6993 1920 6993 0 clknet_1_1__leaf_CLK
rlabel metal1 7152 20276 7152 20276 0 cyclic_flag_0.FINAL
rlabel metal1 6384 6919 6384 6919 0 net1
rlabel metal1 4368 16317 4368 16317 0 net10
rlabel metal1 6480 9583 6480 9583 0 net11
rlabel metal1 6048 21645 6048 21645 0 net12
rlabel metal1 5520 22940 5520 22940 0 net13
rlabel metal1 5880 23643 5880 23643 0 net14
rlabel metal2 9360 23976 9360 23976 0 net15
rlabel metal1 5911 23569 5911 23569 0 net16
rlabel metal1 2928 7622 2928 7622 0 net17
rlabel metal1 9408 2997 9408 2997 0 net18
rlabel metal1 9456 19425 9456 19425 0 net19
rlabel metal1 3744 21645 3744 21645 0 net2
rlabel metal1 9792 6327 9792 6327 0 net20
rlabel metal1 9648 8325 9648 8325 0 net21
rlabel metal1 9744 10989 9744 10989 0 net22
rlabel metal2 9840 14208 9840 14208 0 net23
rlabel metal1 9696 15651 9696 15651 0 net24
rlabel metal1 9696 18315 9696 18315 0 net25
rlabel metal2 9840 21201 9840 21201 0 net26
rlabel metal2 9840 23199 9840 23199 0 net27
rlabel metal1 1728 15429 1728 15429 0 net28
rlabel metal1 2112 16095 2112 16095 0 net29
rlabel metal2 5808 5809 5808 5809 0 net3
rlabel metal1 3408 12099 3408 12099 0 net30
rlabel metal1 4560 2997 4560 2997 0 net31
rlabel metal1 5520 10101 5520 10101 0 net32
rlabel metal1 6624 2997 6624 2997 0 net33
rlabel metal2 7920 4884 7920 4884 0 net34
rlabel metal1 9024 8103 9024 8103 0 net35
rlabel metal1 9840 2997 9840 2997 0 net36
rlabel metal1 9648 8769 9648 8769 0 net37
rlabel metal2 4272 23754 4272 23754 0 net38
rlabel metal2 1776 20720 1776 20720 0 net39
rlabel metal1 3120 17649 3120 17649 0 net4
rlabel metal1 2208 22755 2208 22755 0 net40
rlabel metal1 3600 21201 3600 21201 0 net41
rlabel metal1 4416 17205 4416 17205 0 net42
rlabel metal1 4800 25789 4800 25789 0 net43
rlabel metal2 6768 24975 6768 24975 0 net44
rlabel metal1 4752 25604 4752 25604 0 net45
rlabel metal1 6480 22977 6480 22977 0 net46
rlabel metal1 6048 23865 6048 23865 0 net47
rlabel metal1 3168 22311 3168 22311 0 net5
rlabel metal2 3312 23421 3312 23421 0 net6
rlabel metal1 3360 22977 3360 22977 0 net7
rlabel metal2 2640 23014 2640 23014 0 net8
rlabel metal1 4800 16983 4800 16983 0 net9
<< properties >>
string FIXED_BBOX 0 0 11722 28874
<< end >>
