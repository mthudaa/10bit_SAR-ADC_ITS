magic
tech sky130A
magscale 1 2
timestamp 1749010377
<< locali >>
rect 151 -3707 379 -3667
rect 536 -3717 657 -3677
rect 1009 -3716 1326 -3676
rect 1976 -3717 2190 -3677
rect -435 -4469 -301 -4429
rect 126 -4453 379 -4413
rect 532 -4443 628 -4403
rect 1009 -4443 1326 -4403
rect 1972 -4443 2190 -4403
<< viali >>
rect -351 -3701 -291 -3641
rect -171 -3700 -111 -3640
rect 23 -3707 63 -3667
rect 882 -3728 942 -3668
rect 2415 -3724 2475 -3664
rect 2824 -3718 2864 -3678
rect -251 -3894 -211 -3854
rect -251 -4266 -211 -4226
rect -631 -4462 -571 -4402
rect -171 -4478 -111 -4418
rect 13 -4463 73 -4403
rect 678 -4453 738 -4393
rect 2415 -4456 2475 -4396
rect 2824 -4442 2864 -4402
<< metal1 >>
rect 1060 -3423 1070 -3363
rect 1130 -3423 1140 -3363
rect -181 -3567 -171 -3507
rect -111 -3567 678 -3507
rect 738 -3567 748 -3507
rect 2578 -3577 2588 -3497
rect 2668 -3517 2678 -3497
rect 2668 -3577 2927 -3517
rect -363 -3641 -279 -3635
rect -641 -3701 -631 -3641
rect -571 -3701 -351 -3641
rect -291 -3701 -279 -3641
rect -363 -3707 -279 -3701
rect -183 -3640 -99 -3634
rect -183 -3700 -171 -3640
rect -111 -3700 -99 -3640
rect -183 -3706 -99 -3700
rect 3 -3717 13 -3657
rect 73 -3717 83 -3657
rect 870 -3668 954 -3662
rect 870 -3728 882 -3668
rect 942 -3728 954 -3668
rect 870 -3734 954 -3728
rect 2403 -3664 2487 -3658
rect 2403 -3724 2415 -3664
rect 2475 -3724 2487 -3664
rect 2403 -3730 2487 -3724
rect 2812 -3678 2927 -3668
rect 2812 -3718 2824 -3678
rect 2864 -3718 2927 -3678
rect 2812 -3728 2927 -3718
rect -263 -3854 13 -3844
rect -263 -3894 -251 -3854
rect -211 -3894 13 -3854
rect -263 -3904 13 -3894
rect 73 -3904 83 -3844
rect 2405 -3904 2415 -3844
rect 2475 -3904 2927 -3844
rect 2791 -4100 2873 -4026
rect -263 -4226 13 -4216
rect -263 -4266 -251 -4226
rect -211 -4266 13 -4226
rect -263 -4276 13 -4266
rect 73 -4276 83 -4216
rect 666 -4393 750 -4387
rect -643 -4402 -559 -4396
rect -643 -4462 -631 -4402
rect -571 -4462 -559 -4402
rect 1 -4403 85 -4397
rect -643 -4468 -559 -4462
rect -183 -4418 -99 -4412
rect -183 -4478 -171 -4418
rect -111 -4478 -99 -4418
rect 1 -4463 13 -4403
rect 73 -4463 85 -4403
rect 666 -4453 678 -4393
rect 738 -4453 750 -4393
rect 666 -4459 750 -4453
rect 2403 -4396 2487 -4390
rect 2403 -4456 2415 -4396
rect 2475 -4456 2487 -4396
rect 2812 -4402 2927 -4392
rect 2812 -4442 2824 -4402
rect 2864 -4442 2927 -4402
rect 2812 -4452 2927 -4442
rect 2403 -4462 2487 -4456
rect 1 -4469 85 -4463
rect -183 -4484 -99 -4478
rect 2405 -4607 2415 -4547
rect 2475 -4607 2927 -4547
rect 1060 -4756 1070 -4696
rect 1130 -4756 1140 -4696
rect 2783 -4764 2865 -4690
<< via1 >>
rect 1070 -3423 1130 -3363
rect -171 -3567 -111 -3507
rect 678 -3567 738 -3507
rect 2588 -3577 2668 -3497
rect -631 -3701 -571 -3641
rect -171 -3700 -111 -3640
rect 13 -3667 73 -3657
rect 13 -3707 23 -3667
rect 23 -3707 63 -3667
rect 63 -3707 73 -3667
rect 13 -3717 73 -3707
rect 882 -3728 942 -3668
rect 2415 -3724 2475 -3664
rect 13 -3904 73 -3844
rect 2415 -3904 2475 -3844
rect 13 -4276 73 -4216
rect -631 -4462 -571 -4402
rect -171 -4478 -111 -4418
rect 13 -4463 73 -4403
rect 678 -4453 738 -4393
rect 2415 -4456 2475 -4396
rect 2415 -4607 2475 -4547
rect 1070 -4756 1130 -4696
<< metal2 >>
rect 1070 -3363 1130 -3353
rect -631 -3507 -571 -3497
rect -631 -3641 -571 -3567
rect -631 -4402 -571 -3701
rect -171 -3507 -111 -3497
rect -171 -3640 -111 -3567
rect 678 -3507 738 -3497
rect -171 -3710 -111 -3700
rect 13 -3657 73 -3647
rect 13 -3844 73 -3717
rect 13 -3914 73 -3904
rect 13 -4216 73 -4206
rect 13 -4403 73 -4276
rect -631 -4472 -571 -4462
rect -171 -4418 -111 -4408
rect 678 -4393 738 -3567
rect 678 -4463 738 -4453
rect 882 -3668 942 -3658
rect 13 -4473 73 -4463
rect -171 -4551 -111 -4478
rect 882 -4551 942 -3728
rect -171 -4611 942 -4551
rect 1070 -4696 1130 -3423
rect 2588 -3497 2668 -3487
rect 2588 -3587 2668 -3577
rect 2415 -3664 2475 -3654
rect 2415 -3844 2475 -3724
rect 2415 -3914 2475 -3904
rect 2415 -4396 2475 -4386
rect 2415 -4547 2475 -4456
rect 2415 -4617 2475 -4607
rect 1070 -4766 1130 -4756
<< via2 >>
rect -631 -3567 -571 -3507
rect 2588 -3577 2668 -3497
<< metal3 >>
rect 2578 -3497 2678 -3492
rect -641 -3507 2588 -3497
rect -641 -3567 -631 -3507
rect -571 -3567 2588 -3507
rect -641 -3577 2588 -3567
rect 2668 -3577 2678 -3497
rect 2578 -3582 2678 -3577
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749010377
transform 1 0 -87 0 -1 -3394
box -38 -49 326 715
use sky130_fd_sc_hs__inv_1  sky130_fd_sc_hs__inv_1_1
timestamp 1749010377
transform 1 0 297 0 -1 -3394
box -38 -49 326 715
use sky130_fd_sc_hs__inv_4  sky130_fd_sc_hs__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749010377
transform 1 0 585 0 -1 -3394
box -38 -49 518 715
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749010377
transform 1 0 1161 0 -1 -3394
box -38 -49 902 715
use sky130_fd_sc_hs__inv_8  sky130_fd_sc_hs__inv_8_1
timestamp 1749010377
transform 1 0 2025 0 -1 -3394
box -38 -49 902 715
use sky130_fd_sc_hs__nand2_1  sky130_fd_sc_hs__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749010377
transform -1 0 -87 0 -1 -3394
box -38 -49 326 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749010377
transform 1 0 201 0 1 -4726
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_1
timestamp 1749010377
transform 1 0 1065 0 1 -4726
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_2
timestamp 1749010377
transform 1 0 201 0 -1 -3394
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_3
timestamp 1749010377
transform 1 0 1065 0 -1 -3394
box -38 -49 134 715
use sky130_fd_sc_hs__nand2_1  x1
timestamp 1749010377
transform 1 0 -375 0 1 -4726
box -38 -49 326 715
use sky130_fd_sc_hs__inv_1  x3
timestamp 1749010377
transform 1 0 -663 0 1 -4726
box -38 -49 326 715
use sky130_fd_sc_hs__inv_1  x4
timestamp 1749010377
transform 1 0 -87 0 1 -4726
box -38 -49 326 715
use sky130_fd_sc_hs__inv_1  x6
timestamp 1749010377
transform 1 0 297 0 1 -4726
box -38 -49 326 715
use sky130_fd_sc_hs__inv_4  x8
timestamp 1749010377
transform 1 0 585 0 1 -4726
box -38 -49 518 715
use sky130_fd_sc_hs__inv_8  x10
timestamp 1749010377
transform 1 0 1161 0 1 -4726
box -38 -49 902 715
use sky130_fd_sc_hs__inv_8  x12
timestamp 1749010377
transform 1 0 2025 0 1 -4726
box -38 -49 902 715
<< labels >>
flabel metal1 2878 -3567 2918 -3527 0 FreeSans 400 0 0 0 IN
port 0 nsew
flabel metal1 2878 -3717 2918 -3677 0 FreeSans 400 0 0 0 CLK0
port 1 nsew
flabel metal1 2876 -3894 2916 -3854 0 FreeSans 400 0 0 0 CLKB0
port 2 nsew
flabel metal1 2876 -4443 2916 -4403 0 FreeSans 400 0 0 0 CLK1
port 3 nsew
flabel metal1 2877 -4597 2917 -4557 0 FreeSans 400 0 0 0 CLKB1
port 4 nsew
flabel metal1 2820 -4082 2860 -4042 0 FreeSans 400 0 0 0 VDD
port 5 nsew
flabel metal1 2807 -4748 2847 -4708 0 FreeSans 400 0 0 0 VSS
port 6 nsew
flabel space 2503 -3833 2543 -3793 0 FreeSans 400 0 0 0 VSS
port 7 nsew
<< end >>
