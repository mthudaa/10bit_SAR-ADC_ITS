magic
tech sky130A
magscale 1 2
timestamp 1749411235
<< viali >>
rect 8835 -8 8869 26
rect 10702 21 10736 55
rect 20924 2 20958 36
rect 22791 -8 22825 26
<< metal1 >>
rect 11222 6278 11232 6374
rect 11328 6278 11338 6374
rect 12158 6119 14974 6375
rect 16686 6119 19502 6375
rect 20322 6278 20332 6374
rect 20428 6278 20438 6374
rect 11318 264 11328 360
rect 11424 264 11434 360
rect 12158 264 14974 520
rect 16686 264 19502 520
rect 20226 264 20236 360
rect 20332 264 20342 360
rect 20754 116 20764 168
rect 20816 116 20826 168
rect 10685 55 11048 64
rect 8823 26 8881 32
rect -1 -8 8835 26
rect 8869 -8 8881 26
rect 10685 21 10702 55
rect 10736 21 11048 55
rect 10685 12 11048 21
rect 11100 12 11110 64
rect 20754 -7 20764 45
rect 20816 36 20975 45
rect 20816 2 20924 36
rect 20958 2 20975 36
rect 20816 -7 20975 2
rect 22779 26 22837 32
rect 8823 -14 8881 -8
rect 22779 -8 22791 26
rect 22825 -8 31660 26
rect 22779 -14 22837 -8
rect 10838 -403 10848 -305
rect 10946 -403 10956 -305
rect 20704 -403 20714 -305
rect 20812 -403 20822 -305
<< via1 >>
rect 11232 6278 11328 6374
rect 20332 6278 20428 6374
rect 11328 264 11424 360
rect 20236 264 20332 360
rect 20764 116 20816 168
rect 11048 12 11100 64
rect 20764 -7 20816 45
rect 10848 -403 10946 -305
rect 20714 -403 20812 -305
<< metal2 >>
rect 11232 6374 11328 6384
rect 11232 6268 11328 6278
rect 20332 6374 20428 6384
rect 20332 6268 20428 6278
rect 11328 360 11424 370
rect 11328 254 11424 264
rect 20236 360 20332 370
rect 20236 254 20332 264
rect 20764 168 20816 178
rect 20340 116 20764 168
rect 11048 64 11100 74
rect 11100 12 11353 64
rect 20764 45 20816 116
rect 11048 2 11100 12
rect 20764 -17 20816 -7
rect 10848 -305 10946 -295
rect 10848 -413 10946 -403
rect 20714 -305 20812 -295
rect 20714 -413 20812 -403
<< via2 >>
rect 11232 6278 11328 6374
rect 20332 6278 20428 6374
rect 11328 264 11424 360
rect 20236 264 20332 360
rect 10848 -403 10946 -305
rect 20714 -403 20812 -305
<< metal3 >>
rect 11222 6374 11338 6379
rect 20322 6374 20438 6379
rect 11222 6278 11232 6374
rect 11328 6278 20332 6374
rect 20428 6278 20438 6374
rect 11222 6273 11338 6278
rect 15782 744 15878 6278
rect 20322 6273 20438 6278
rect 15772 648 15782 744
rect 15878 648 15888 744
rect 11318 360 11434 365
rect 20226 360 20342 365
rect 11318 264 11328 360
rect 11424 264 20236 360
rect 20332 264 20342 360
rect 11318 259 11434 264
rect 20226 259 20342 264
rect 10838 -305 10956 -300
rect 20704 -305 20822 -300
rect 10838 -403 10848 -305
rect 10946 -307 20714 -305
rect 10946 -403 15782 -307
rect 15878 -403 20714 -307
rect 20812 -403 20822 -305
rect 10838 -408 10956 -403
rect 20704 -408 20822 -403
<< via3 >>
rect 15782 648 15878 744
rect 15782 -403 15878 -307
<< metal4 >>
rect 15781 744 15879 745
rect 15781 648 15782 744
rect 15878 648 15879 744
rect 15781 647 15879 648
rect 15782 -306 15878 647
rect 15781 -307 15879 -306
rect 15781 -403 15782 -307
rect 15878 -403 15879 -307
rect 15781 -404 15879 -403
use sky130_fd_sc_hs__buf_16  sky130_fd_sc_hs__buf_16_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1704896540
transform -1 0 10848 0 -1 312
box -38 -49 2150 715
use sky130_fd_sc_hs__buf_16  sky130_fd_sc_hs__buf_16_1
timestamp 1704896540
transform 1 0 20812 0 -1 312
box -38 -49 2150 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hs/mag
timestamp 1749010377
transform -1 0 8736 0 -1 312
box -38 -49 134 715
use sky130_fd_sc_hs__tapvpwrvgnd_1  sky130_fd_sc_hs__tapvpwrvgnd_1_1
timestamp 1749010377
transform -1 0 23020 0 -1 312
box -38 -49 134 715
use th_sw  th_sw_0
timestamp 1749388026
transform 1 0 369 0 1 132
box -369 -132 15509 6243
use th_sw  th_sw_1
timestamp 1749388026
transform -1 0 31291 0 1 132
box -369 -132 15509 6243
<< labels >>
flabel metal1 -1 -8 33 26 0 FreeSans 400 0 0 0 CKB
port 0 nsew
flabel metal1 31626 -8 31660 26 0 FreeSans 400 0 0 0 CK
port 1 nsew
flabel metal3 15832 6306 15866 6340 0 FreeSans 400 0 0 0 VDD
port 2 nsew
flabel metal3 15706 294 15740 328 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal1 13525 6222 13559 6256 0 FreeSans 400 0 0 0 VIN
port 4 nsew
flabel metal1 18101 6222 18135 6256 0 FreeSans 400 0 0 0 VIP
port 5 nsew
flabel metal1 13533 411 13567 445 0 FreeSans 400 0 0 0 VCN
port 6 nsew
flabel metal1 18092 413 18126 447 0 FreeSans 400 0 0 0 VCP
port 7 nsew
<< end >>
