magic
tech sky130A
magscale 1 2
timestamp 1749046477
<< metal1 >>
rect -608 1136 -400 1234
rect -348 1136 282 1234
rect 334 1136 542 1234
rect -514 872 -504 924
rect -452 872 -317 924
rect 283 828 490 880
rect 542 828 552 880
rect -618 723 -608 775
rect -556 723 -317 775
rect 283 723 386 775
rect 438 723 448 775
rect -608 -34 542 64
rect -514 -759 -504 -707
rect -452 -759 -317 -707
rect 283 -759 490 -707
rect 542 -759 552 -707
rect -618 -908 -608 -856
rect -556 -908 -318 -856
rect 283 -864 386 -812
rect 438 -864 448 -812
rect -608 -1204 -400 -1106
rect -348 -1204 282 -1106
rect 334 -1204 542 -1106
<< via1 >>
rect -400 1136 -348 1234
rect 282 1136 334 1234
rect -504 872 -452 924
rect 490 828 542 880
rect -608 723 -556 775
rect 386 723 438 775
rect -504 -759 -452 -707
rect 490 -759 542 -707
rect -608 -908 -556 -856
rect 386 -864 438 -812
rect -400 -1204 -348 -1106
rect 282 -1204 334 -1106
<< metal2 >>
rect -400 1234 -348 1244
rect -504 924 -452 934
rect -608 775 -556 785
rect -608 -856 -556 723
rect -504 -707 -452 872
rect -504 -769 -452 -759
rect -608 -918 -556 -908
rect -400 -1106 -348 1136
rect -400 -1214 -348 -1204
rect 282 1234 334 1244
rect 282 -1106 334 1136
rect 490 880 542 890
rect 386 775 438 785
rect 386 -812 438 723
rect 490 -707 542 828
rect 490 -769 542 -759
rect 386 -874 438 -864
rect 282 -1214 334 -1204
use pd_in_half  pd_in_half_0
timestamp 1749043030
transform 1 0 -496 0 -1 793
box 96 -441 830 827
use pd_in_half  pd_in_half_1
timestamp 1749043030
transform 1 0 -496 0 1 -763
box 96 -441 830 827
<< labels >>
flabel metal2 -596 -434 -566 -404 0 FreeSans 400 0 0 0 INP
port 0 nsew
flabel metal2 -492 -509 -462 -479 0 FreeSans 400 0 0 0 INN
port 1 nsew
flabel metal1 -2 0 28 30 0 FreeSans 400 0 0 0 VDD
port 2 nsew
flabel metal1 -30 -1169 0 -1139 0 FreeSans 400 0 0 0 VSS
port 3 nsew
flabel metal2 395 409 425 439 0 FreeSans 400 0 0 0 A
port 4 nsew
flabel metal2 498 410 528 440 0 FreeSans 400 0 0 0 B
port 5 nsew
<< end >>
